

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
DKaw2YF5X/sI0l9aLdTgbK/M5GUdtEMTnIFmxvSMohXCNpaRunL9ipaA59Dc71YrenIGtec5QT4M
zCoGKmFbyA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
QRHRuF+/6jbJdc98CuDuU1RSPkw4Mrd2rWInSv90clZq9I1OTAA5/xdv3Hk99Vg2prXDV3YjNqoB
pcpnTJxql+YZ6VAzN0qCk+oUeO1cCu3qiinofcBjVXCdgYxomUKUeE7FJeYz3Js2G/kJGoeHFW9U
+zAl6jadwyF9Jbvv+i4=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Lb7wQIOJLuT7MorOQ8eHbXO7nLYJ4w6DRb/CRc0KXgD29tV/pKu8nH2e+iVICJbGwJJtQ3k8P1j/
LscOU8Hk23tTbvsi/KP4jYIAhUNpSlUfm6H0KJ2yht05tm7/nGOSq+YwUD5ni46LH6TZmw9wRjLo
RAHSpBohLboc3y/hVTXta9kQmKPnqAmdZWZqkVyyS5o93+63/fdqbFaxxtwx1mXeZDQ2+2zbTCKf
tbrO065IQsNhLqpQ6GmWS0y4Yk762FiY/PW8xLoCZ1V1Fh8ocFk7LKyATUlQjo3T4vsNks0JLfh6
k4wW0gpjLf86zBHim396ye0D0jCoECOhPpGtaQ==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ZXacKhqAwgw8zLrWO0Oej9oQ1uNqsfSW24Ju9AdSqiO9hJgeX3QSs/Auka01BXmxZF02hREfAK/G
6uXtwOuytUDW3C0vu69znjuzfKa65iqAvitXfuV2wV2SBDUohxstI576S9cHfGPfoJ7tVzjIg2t8
+fXxMYGWVW/hL5Dt3LeBc+ul5BEG9/vwugVmMP2uMG9nGEtDEQeLb7bWAsdsP6jyz5L4K49swiWc
6TrDCW/53r7o1y18s7qcumMrH+8e09lZWlV7gV/qSGCmNFjNoXkvbq7X5+RT29nF6kaEY/1Y1wcM
sqDv/0rI3Yh5PZatD+o2YnHnz7Es16C87EBZrw==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pkb010SLYsAhKXcWm+QlAA9Be33Kx3pWG3KQ8c4OXZxiNI+ziOzdNGDZkUALVJhYeeODAczIsICK
xPobg5BZJdmnFjXMkYzJiVNc7H8OtQ+xwCOlZfGQy0nG30bs3aCt+0ciZZz0ed8EJ3QfOUNUrA8S
ACDctQvzk535zqal7JGqVOcbax0rksASegZXl9TYHMAWSFXsQNDtHG7HCq8QaEGySiiJnEz1Zygi
CXmAaOXrSZ/75eRU/jV0Zmfl2uX9M3RD4WyT2L0mtTPVI1Jo5riNKDciMqi09G5yCgGBizlVK0Le
ynsKW0Fvo5j+TrmGuES2+DcsvwzxQUmrQ9n9YA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
saU9xQVocYCNVhmm+/jaIKt7f7lGDiBCwD7GUeN8jk+fV3dDx7VH8BXnwqh3bO2UtgQTq4TYazR5
PsEJU9lk5Y+2uIztywixaUOcY0t6PGvi6DZ5S1UapcNaqz1GzVDJNMdFrGWeodfXgyVpIeng6Jtk
EKceFNW0p1SgbLjlCjU=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pbTosJ4LwLIDFDsIbDQWyryoCwFpua23V6z9HaJa95eQ/VgCaYwQRc0pJmp/UgRFI8GxRIcCfLjR
nDQiDTQUzYsgXuFi39wSqyum1ybk+zJc/c0tfa3zo7fAh7WEKBR6EfegxJoOfQ6umn8yMUOq35ku
5cQGVgAH0mV2j7kgcszzSTcMNu1shLKlPJejpCdXAsAct77F4/JiYgr35R62Nw5TiOPHxLGWKlD0
S4rOzGqDzYI4jb5eYbnrBMtpHWXse9ybFZPj47SvpsioKcFIHeUE7GrNOvNDQPdNPahScNll6gSb
fa6tuXH+3Q3DQNGg7RW23POGEp2w+WE6Kef4qQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 74224)
`protect data_block
0pR4qYYHrD92Vr2lltbDGBYi94yA5NimRwES1b2SJNOcuW0dbY2DWegKuGXMbI+wlmb0QzXCX3m4
uxs0DjvI9veZcNFHdAlsLjcQIJlYHEzKBEMvZ/nVYjtEq0+r3G2HDX2cOn/axZ1tHlSH3+vW2jIu
fEdc3J1yxR8Qqlqs/yNzfe3UeyultfOgRRgzhqu3pban25qNyVOW9qU4vlETy+hLjjegdRCc8P8b
h14jKQkC4/ynl/fVzCiT4etTlYzArNsNG3m1KdGnzHpyrIv7f6Kmg/t2p+rrNeJampUBIPiNXA8Q
xLFSwRyHhQ+dP/2AVQnc3HAPs9se2rt1dTDJFPFlmoLjjGtG4bXP+hSx2Fula0rlf9FhoWc1/ezP
Kmvmhf10h6ueREoY2m2nb+Nj9eIlkm68d1rmAcWHx+sGPJat/un1yUOE4WPrf4dG5gAQrqMHfXSH
jOrtoA5X2ukdz09cHSUx0Gxh1coPZBGEiDMn1hudbm8eq7Cp66pFMPfgJyubVbvBeBa7cB2xSsWq
yqIBdEax1GMpnwRp47q2Ft6417vQ64kzKiyK326S4OCQdzDjGV65O5mRfvmH8b3qlLFHiA5iPcuI
d2H4EZu/STykKCz7KKKKukqwb0uehkLB2efy2qzJGsCOBhx/uqSTSI3aLhDDtP2EOnJ/tEFkZV6P
mUahSaMHujmjPiWNLzPV3zjPGr/+gcPEhM0SDrUscBU4eRK49NaAfj0Fz5DPcstYMRgoHqOvUj8u
eOpJL7I/y4K7i3a/HPWNIeOwXzTpo8jQYENwg1rulbOkY3O/EDvL5DEat+J2noqVa1/NfA00FdDK
dz+hOv33C7YOA/mOT9wQ2rHHkbr0PZ+aXsEurZ8zS0HAvEBmthjvJ4kXEkXNY5h3/J4/xzTfmiJ0
QQjMs5qI7EVuxk9L2F72ZLVNV3WB6KVfMix31V33fahyuFrjAyp8c4LN/iAljwW0xxH1CGw++ibX
T1QOtLVHT+2Rk10Xp5xNM3FbJSz8kcc0m6Ffxn8s+1Y2yS3vtx1utzXBJId2yNtBCIWJ60QqXsxl
P99T1NUO5Nq7QQnCJCvC/fhSBzjgZRsIUAW8PvS5/0ovWZxf7XgvTtAXAdhrHNkJNRZl5UuL5S7A
uGs36vZbDGV2/bEkT6bapmfFJZvgDamTHO8sTZ9baiXWIPG+tnmQts6m6QLkZMiTLGEzFIPyZU5d
2DYd3xxxh8fDux4Elsz3ESz10GZyiCDJ/iHAHxj9iVHUsCzeGXqwWnnbZF5Nh+GaWqFcQLq9opB/
ea7TFFyPUEyH1pdRhiIA255oAoqD0ZYPHFJkHnA460erCz9DjlRpO8saqOi6EF5xFMWV4UkeyBqk
W6lfnkZEBEHQEUTLCOQaX6MCm5aOg6TLM9VuJ6vQQ6WHCoern7vKoUgh1OMoR2LtBKFug4tF56Af
avvWReyIezuBpLa4IEEx2i1C1yCiaDIcK4kPrZ8qqgNPDSEteODgzZtqxiWP1BCqlWyXSa8XVUIy
JlrNMlG1Nlrfh5ZadCM7yoyd6Fn7Qn/+3KjqVZkS/DG9kAVKNMCO//2Wz0oEYH55QHd24JKJAloH
mh4Vh97IignRgU4jYPSbpXEFQ7TyTRjBDnaeLXVw1H+lPOrYylWGTQqyRWD4Mg7vbSFRlGe54G9e
ofP62dS3PXrk9hrc9iAtVOUs1mgX6b77p9GQBqmF1OeYPO491hNV8MqWr+KgiGgydbDLrbv7hgl1
Ub+0z0al7rfyodDrk3+X3Pyp9brVY/IBLvfLF4kerZpIBt1LX2labdiSQ0YEFc5B1WPnBOiFH2Od
u0pvAEax3jC3Zyhk4XqM/ioLCHjayaErd5nk5eBySsySQnair2ObxZP0zra+wpVqVPSjVxoQFMtM
X23ggNoEuABBagETw9+pfd08ybayBRY8x3bSC1iUqZtZR5IyCsMVKUjvKXDx/wcPsmWyGz89n6rm
MANItc56suSM3SBX3mgyroxkC6hNMQzQOfR7KbP1ddf6IlfP/UCrOkdzCXc4yIc8pxh6AfEjMk7g
pedXRAZIHH8QTn2Fd6zTsY4v1hlmQnuGwEq5qhWs9MT/EzWIgw3zYDWBgMtv5HwxdJ18IBkl+pjC
nCAcqZ42EuK/BFLl25bHiTnzZLwcdU78iMWkK2VaFs0HdddyTKokFFsG2si/vwYdyoVOZWvmC3YA
y7+v+8rWZqbNo9mq7L1D8rIDnpGgkOKh/eudjDh+SEcwQjuOlbDYas0mVPHLa03Vi+PkK1AHRbJo
MqyVu9pK3D6lkacal1m78ycO3xCF9fgdahw+BAO6b5mbUg2PwfCG2y3HP3kja6g9tpMfqwuVqpXU
AaE6GYOOojmFZgYnmA5wD09UoDbbuxCyKQF3gCeFRniv4WtxiWsSw40cImXsQfesCpCSbHRNr5jg
C//DHxemPkW394uDja8HrTY5qNXPZpgMUVI0hqCaZFe8j8Z81URdKEGTkxqw/O9VHhI21nt4SUew
O5lUwuvdG2F8ptIHYBDe0bTHCjFwkdhERqFtvfurtwMR+ewMevP9eyBIquS+1fBmb5ZXgUUydCE7
nHHV0nmA1K0BoiSKPtooPG+i3z5h0uheIQi8kzZtSJva4zJiKnOW/3ZfFNbBe2nKTKV1FjmOx0es
+gDetMquR8utC+nVDMNWYxSK6cifME0Elx5WcPFUFi5WsgJVsMa1jnVaJvr/p8piSjXLlbDh5WN/
h++/FX50+WIkb6PP3oW6N9W0l+bIi5XYHJBZojAt2ysK82r26En6pccWIiIN8u4SyBDXOFEpGAfV
RXeR4N99mWDSLe5r9qR9CPw7E/Atz1fR5S81t0/SJSesvCDPJWqIWR5lxueSM0EIvjxkXgpbU6CR
QkmQBdc3iypEUSS7BUBrNAqHOetlMB/raEwsQApTt2S6OrE+pNE8+u1J5P7zlZVamZq4dtboOKoR
erEo+bSXx81HMZufaaQ2qNmPJz3mcmolshNMFpINKjb+rPvm01h33LV8ryBmItwMZOj5XYe6ChjT
WP3TRGUnSHkxSs6LPu47AbVJdFRVuDZJW9HvwSWlMnfQVmMomrXAdtATKShupZ8+EHcaERQUIJPo
mvHIO9tYoGMcztTa2qQegUhB/r7LtHSVJxILDLKQbsAsljspWAycwTHuT+s5YI/lagiuUkfZeZ31
UKBlrYpFh9CLWKy3EuLs6D40rPuAUgN5YHZUmFqT+hcRY+DQjrpngx3PSGl4DWCdIuX4WIRpnKk1
7whcfd6nvTCclyMWBOYtylET2qNd0yXnurvGW/9q0sB0rCyrCviKEQs+LJwI0IIQk9TW6GFW71S3
6rk8xGFL7bRJ0ghkmMaJURrF4d0DQWGOGNwKy7sX7rs+nwZYn1YDsHmYOW92wXFR9LrjtsufEuw6
eNwWjQx4abIh3VjP6PZ25tI+d7zhbggmbVjgZO6ID1PyWqvp7xL9vBF7aHykoOjpI3pe6geaeLs8
JHRP82xIzHdtvB7dNV1hpDps5sk3phXukfhWomDPzsBmO+PHyvkKzQInmmn3eR7SzDPaVAdZAnh9
pY0TerPPr/IkxZMbLdab7F4fQp+fSMAG7r6Q4kTjhlR2j18kw+A0tHed+PZd8moX0zdQ1Ay6Rw9R
O69C+ttmrOy9eAOpALVzNzeXdaKgnTNjHbzQWhY7si5ok0uQdPEcqJZFxp6il19KV0lrogIfafUI
YNtrOWf/v03lt5M9CWWkjzUVKUHNKoep7trl1f7XX6+xdG06QeZpCgeWKzAzVr2JSjeMegEYBZ0e
0t3iZ1TZQiG7NTlg3Fg4w0egCKfrFfTl0msXDs7iKahWDShn9ZkS6wUDmM8WDTpI4tLI4CJY9OHq
OwGG0e3G0V8p9z2lm8f77d+AQ256p3H3w8D54CbA6GGFK71wae0676vLsMNoB8ZY5ctn3fMkV1ej
qR5SQWYjJofdXsZvcgwTxGSjo+gRh/GBFFLtqyWrY1lQUiWxlO5v/Nx8uCFqRezfHHYxwH5875aZ
B+yCKXOSQPwoFc2AlFTPksGEK+rjrWvIcK4voDcfhe8M9ZNimo8FCj5DsIacJDE7EDeX8RsGu+dJ
/WooCJEPUC0QJ+u9PCkd+Cb4DeKInC9y64CBHYF4QfRBTICGIDojv48yScpcHkALgK8mZkJNtX8G
jTlw2dA1bl0Dh0hXhZblQ06lQ36UCS3WqZ+oHg/K7W/umY3e1WjjGnpG16Jc8/PftleegwK3xPl2
UQk+UZU9jqbaTQj+LStFQy+IKMJ6hPz4moFq12OT4OKXgBdGoUfh4odDjr8X9oZilHvEcAi8LW/s
ALlsucn4/8ZkzaAqf8hOsKE330s30HDuYfMfUaS1VRz2kHBMc/tBoV8upr599vhfwH15621n6wtB
Ds8j1L1UKs4wg97chaXY7u4abInNTCnOZkwhHGff2sL0O40q/owfttEm0ooVutCS+TeQl3ZMeZig
PUdiMHAEHOgttwPrYHJM4ylrSxsVS8WfN6p5pJFa8dQ6lI5pRaizY06sDsLVmfq865YQ17RXfF5u
5Td5ely+zU1btOts768SUd5rct+mYSHXj0y7/vL40cW7QMaKjSYZIMrcnMPynDphqSOeGVXCR3Vu
CJVDkGeahVnCar2sBHQPceOYtfH2B0nuOi8UKrGv8m0o9BHX26tjY3WrlrcoybNcrSy8AIYjnc86
UKjKrFnoDfTvH+prYiAiSWMwYGYpEBOy/5Ysw8SpCRK7x16reT1eow3KXtGnrP54EgnKod7s8dLJ
hCO+btX5uS2iNZyiOFMngj6ih4QRAWuAp9s54GzsbkLeXIqkSk92x/tKJLqYy+4bLm6tAMqCa1PD
cHEhuOkGBgxKw66qS27n1ujLCzrnr/zzGxOybYLhdUz9MZtW0HHo3jBULECKEoLgi8ZAIU7i9lNY
WYHChnu4VbeNa78qylQLOewjjEMYZJwPt5jJ0XhDCyye9HCk+zXdYrymLG6ujlwr4DohnnKMFT0O
pXbBTxHj3qqwF+zpn0uOpYAn8ODbCOYF+DhKDn+HrgYpNQQmAtckYkigQSytbD6NnBEhcDrIdjCg
5dv78qUcrbcTFVi1xOr8GlZ//nOPJww7SiCuHFPf1EnEG449EF5l9w/psSM1F3tp1oRteP92pqRX
eezybcrH43C94NLaHSYA2bUUu8uOJTzbFBIzQw+k2JLXYat6T8FwD/WECa7eosQ1t3MBaItmpFxm
+QfF6vWyCcNHjDIaB92SGOjQzwzeT0FUtDaJxV/p6ZmWecftIUzCmTohmfJfzt4bA4iBgwcHJQSp
1ZIYiBV44v9i5at01c9SsmrpeMtu52Ax8rpyckX00Gl6n6E+wVFpeHx5ztersDbGujimgGmyt9Ih
zcoOY+e33kAzXhxjZGT/CSj8fkTtT6zDVY7nUHZTkU1jfUKTqAwvjAwa42uHqomsJcT9JT8yTvAZ
fm/q9kZx6Q+bCwUQgyjgTdyi93GbRfYXJK6FZHRqQ9LU8ChmV4IDDAfLty5E8pCJWHETHidhMwmL
V3edc321XMl6pe8clN3SGpxFJBHyWttbKaqCFgJCtRUBJ6oUaiKdyP2A4O94TxwTg5mX8tjK1cSh
zSzbzn4frioB8gtu7n3ZoViT90EXy97u0B6LJZH7rfo9XcsREAvVSgDQEEfcgztQryZBkWaHg8f4
eL5TA9JzMTpF3I1G4HRh9t2HRd5ZJJIALlfMpBnwyvQ6eDHDfoEB0qh26f/vXSDlAQWW1CSOwQKS
gS5RKKqT4inOd1I6uhw5gV1jq/EgrlIYe4tSHMlXSjNgprvNhNa6DGA1RsD23RPrpkDPDUmRiR0H
F6KoyICecmUrikzHchfnHVhfU5ChJ7k168yEycGNpdk/p8pcJzOF7IYA4OdrjozLKHRpGnsnUkYE
OBkbFdoWgfuZKw8WArQCsLevkiAqR1SFVsOh1UuDQj03Xy2e6tG0RbycI+RzDboqPNpVkv9oNFBx
lVx1EtfaFgRwXwUMDHOxB8Pq/Nt/VSScpHiRe4W3Qt+ArSr7Xvsvp2r2Rt3MxHH4rSvewv/BdbCC
sujqdgN/HXJiY5hB1fbqmpeLAOFzpddgW7qnF7sfuez3RAaxK3jZrclkEa3mAKqs8CWBoilZ0r4g
pbNpgMss09Jo8E2mS3503+5S9P6MTVaGJK5nqhk4FGtlIQ/caUsK20zTwNmQ85TDM2WtEGbuQ50O
/e9gmJxcJ03AdkKFQ2idiU9i9mvWHm0Unvhi74DefedslWF54w+dTY/gFQaOWMEJ0zRRf7OZw2MO
FNmgmMQElofKVPcb49iYEnEblpZC299dacN3cqZoki7KTQ8lImJFAp3mrU6hgreX7ncGZYGF83on
d92U3kBNaWuZokXkTlGmkTzbQPcVcfMPAM3l3eleHGdZPbXUuJdX56a5DAb34KsxfSA60njeW6wS
rb1KEJf0jZZEw0LRcCPZ84O6neXlOTxyd/O8ISg4+IFdsAYpDfSoKbqA3d8at3PsM6yj3K6GjPi3
m8ziYH/xSTeP4hlnSj49O1K8qtSnDaOO2IAJ5JwfJ2VjGTvenpIsPnud9llSKxQbRk6Ne+rW4AOe
HvUd+VG2EbaDlpcbhn5wdL5/mZG30mOacNXdaR74wRGQ+LBVYBK5B6rWAM3fqHIV9sXNQne/s0AU
9PiTGCM9tKAzOUETGNistukzkfyHkibfCSpLnWDKXG/LMAs863gaw+Uf2sy0zLpT0b0xJNFEZh/6
f5dqbcY7tzXbmvUP18uvgM/3TnhoGtGwEuXAT225ANjbGQ3l6O9TCSwFk/cyX0ZDkcI3HY60Jua6
08kIQsUmvBoMuUCJwoK+8csUQdXoJ8Nu3jemXBO94ekj3c4q6EPVLf2+5JwqtKDPgQSZyXeuCuY0
8okcstVRbOZtspL60WhfrDruUO8sZGp+yFivrftArkxVkQ1SwqXAVkOD3j5bhm1bkK6Zw0tlO5Ba
xRIVQ437EDViy0+Gv2rhetI0ouLJH3rV88W0P8Q2sXQZ5sfTMJ9CWDShG2A0JTY7MsPO6WrcoObm
wFHPPRJptttP7AwyWe5Th1L6LI57S9VV7dp31rx9JqnHNoAspBS1v14eH4zC7rS27pyK0N/7AmXH
zEeQ+B3xnyu6y3U+gab6kvM4KzH8+qA2ZfsNc5QBtIHsy5PEALf4rVWDN+bjoEVGE5s3YEZt9p+Q
296/VoBJ7Rg6XGacbmQMT7MmKDTkbRmgVOh6mAXSTkOvRcKIf+Qs+ayM8OBWcK0yt5DDewJGDEdM
3DSzpiieLAdqACpmsTZev8AGarSKrWMMcCNVv8GRxCCLtp66uMJQjgxEhstv8c4JPRg3+1uTeGWQ
YFFJTqTgv9K48qaTaoF4O03+RUa4cmkutcSd4aanC9q1S3dnM0OfNz7sBqKsx9Ho8tfxBPQV0qfu
9fbvztS2VYbhMDXCLhxurWe/DEkfoDx0O4amXpS/rDZiL0kTqKirXZ3s4Hce9jm/kfIE4Oa3Z9np
w8MWl+jg58DaKsRrv6Tgqnd0I4gi6sK9wpB79rK4J+Gh2/oyUIZCZEGtKNQ9fzBvi/yen1gEoH0D
qFVdPVvZIUhxVEIijRGYjkxCWUH2P4SlhPyiAaHE1NNKc6G5/me5Qz7d6lpzvQF8W4WGMFR9HCHu
4YasDSm4UtTOEfWfpw+K2Nop2LDjjG727ut2KYMbTJrv/CazCRdwAuKEc3MCPiKB8kFrCItLibBl
B24D++1mHpLN/U96qL/SJIxjyRlC6jFkz+VisKhSUNo7lvel35XQcvKztwVA1zgCo2aF83bPh3to
PZSTwCbYljyIvkM0fQhcOvFRUToIS556rzSW1DncC55AXmKgVWtHSdU919WtjV9y0qacpEw6riIi
KCGhmu36oTKhVsC6WMJ7L54E5dyWAnmtIjZmIv7gVm9SxQ+TlhXIcpXMb2h3bNAZCO6SZCsxTjVA
WGgoPz4HZrVR0aS+0UwJSLP9fmXtLiIBS6RAwOyAObbtEclxcLkuPMwY2dUG4jDgd7NfAfXAXQXs
scL1gCIobW5iaLXCR/q5T7BVCLLkVt9vDf2qt7+Mr9zCYtUj1p2+B3ifeSZu60HAvVk4iS+gSxx+
Tg8kzyk5qNGYyOrk14fBLK1J/9rqSEa0ozd/sr32odY3lYuuLB10HbuGlKAf+bV3/nMXN34u2NoV
t7MPREtKw1THt/LfNuh+ikoCvdnL6MIIOQBmf6DraWKjEFp3EA1TF4gPCg3iNhVSmezcAj2kuCO9
o1ubhxyY2Y2CCODdicci7eSF2C4OMmX6uDA0yf2X+il9Yhd63Z+xShY8UYWUM8GzU2JsMF1W5nnz
778cdSKIwBN3UzD5OK4/xegLj5qE+utScB7wQ4yqIrtQswBC7N+tYzA1yaPBpH5MUXL0j2TPP2Z5
ZlDs4DFKhI0ZX5C+eRjncIGhfdstYLWX157DN1siIFnA0+uJxfCENAiZv3zXNftNKAUICUix1dw8
TseL4WDPeylKzTyNyak1OegVSHU7uFtSN7GdgYAMx46RxtMw6yRXKgs8je+7mvZFXwTPdicqTZwq
v24mKHtYytDr+yv1TOaAtFUJaBuQnWN3t+Ptquh6LbbdpNC2Ica5Lp9kwQlbSMflavaoBAoYZ8zn
tnynRa7jVhoVViyelfYqqEEhppEL0ivQtA9emmyNnZekZXe2yeIUHAHPmWnwny1UoNaWxfcOtFAU
fp5bR4JBgOXthmTOAbYUbC7tiR9q6yMwepKOzP7XCPZCRLVIS9gkOmbR5LKt3MQ2YZc/NBOsLKB5
pvxzMUSBQkvfCUOWE+EYvlyF92podDwuKBkF8G6PrrE5kqNYOklwwUUx4VeV+6T2KoWNzWvVxbqT
KrK455DTs6XSGxV+zkpzhscgsbxxGOTL+1Vs83Z5loRy/BqieL0p0JgX0W8FbulWr2OXeiapKLwZ
kIBzVL6w2XaNXCjE6s0LMSfEBgYGwVjLghy9OwrPysWZHNZFZczSZ8AsUC3Idbbhp9fC4+Av8T3K
DSfY6iB44hMQemHl9n/Gj2I7kW0fWfPBWMJIMRaULv2THYvQBbhO3eeQ0IYiYM0AAYCNTYKYpEq8
sITHU16fPBWS1dpy3XLpQ5L3z0WAdB99TxfsdipjDG4mT8FlcJYaIz1SQXyCcBrH96qRk9l1hOxe
nMitieXUoF4yLMAnOuz/oUGS07I4a6DJgNMi2U/1ztzNwFpBJqNHcWLAUbPsCUor10MuocM9Hr3j
HSaLn+shZXQXH97Hs0dDCDDiN9HGuPaqF4x1tSemGefE6l+aHaFXErHpple8cVZRURb4PQ/+VkJ1
Q52Ff0GX33uaiFuakD1Ql2FAfDOyfLfts24KQUgcGVwSZTUOK1Hk09+FqoIczTzjgSe6YEo3p8gQ
WdmpC0kIEkLJahpKVxd0hMnF3zxSH+Yl5qeuBgGaQsMCZpC+EABdZ/Si02ePmfP9uT1H/QKykAHl
3M6EBccHchubOawcqP0Txe3vLNJs+ABMaa5lhNnqN0x96HHs8FdaL30BW1IW+iqnlw5Q4u5FtzKz
plJ8V4/r8Xo2fAQMi0+g0fUzPwJgN9ZDIx2QTzRyrAixCVk+a+6fu+ViJChoV7xQ7o9gFJttmuVw
GTNtE7HmmOEBY/waFDUdg9LXX3F8uxdDtjMZVbcdg6qNsqZ0+eH6W4Zmeq9UDjJilFoUkc4IYMph
52ke+S5eLLabWPOiIF8EoXXCrfTBmYcszwlFIjOyB1o7YzXhi0LSPLqd7CfiQq8chXWVaznAM5zm
R91fkcTmaa/lsdJ7OR2efJnCQPUYRBRLoejXhpoKs23vAUp10raXrBO5zHaP7Q7OLmC0OLFji4t1
JP9yvfPDF+h4LRhkUvxvuKcjMPz6ZN/nlFkacHJeXAlSn5RQByAWkoBWbKcyIQPbVZQtqbDkWktI
Tu0q7kYLxA3JK9PqyPHWfGX4YP5bJWzSCTtV1baYCBVS+sLKiDdq8kj3OrCb5dJuoqY6Y8/wa2ZP
iWfsZhg+7cFLdG1UFsjATrt65OAxfouCocLo3NDtfBl3NnS8XBUNTLnprxUN+8O1qTirbaKG8nre
p6qkuXEJdArOxA3Yl+D+z9MTbnESXBh7zWJCtqCQjEt24PO02B2s6W23Bi6KfTMRtw36GpWuWEj3
pzQn74eZfIFBTSQb4+GbYbM1Oo4VbsuNd8G4wO3qHkWczoGhoIteGdZnWpqKShFEXwXuJjWm/OaN
JbEo0pml+cqjwsPjaHt1hz8h5IJIiPB6hOOFoLcyUXZfKMs/w88yYvhTrHzvAVU7FKR3pGTQJO2v
zm/flWiYfAkNQRajvQEIAFkPC2bSccyRv1bFZDlVRD1oGF+LLVkSDI9DugLVB30QKjIC4dDWF3Oi
rK5P4AWMR6ytBC5LOeKX6ZeS38ncpWq2NAH3J/3PtaUmN5YXudx3HtLwqhCwLS0gEBkSogoWGYj2
zMk4457ZXITti2IgRuV/vul7NFMFeTLo7aAvFepFXi6RVq8rbJJE8pCCz78cevOU1t1SRF+yb5hH
/JCW94NmagSAsWPSw5xZZbXrvKDaH4ra/WmfM/B0u1kmYxBTkrkpjVM+ncx5EBxcu0EaDjamiMro
ut7Z5wh/z5GYMA42ub8vX5vE+mEKGbsHTCjf2Ygk/J+OkTVz4ASJeX9fqpZjTfBdb8tPvtut7m2j
Sw808D+kB5zNwz2X1BjlopfBoHDRYPp4a6ccS4Q7OWum3vwStYztyu42my93BTE8/6e4jlJWSsog
vuhUIUlP2rW6NNqkV844e/4F4ODHQvqQChrIiv1puqb0pKrs1AQFYAeLrvbVJ+NtDFeLaarMrAfJ
aRyaerSrSN/gTggBkyyvbZEWgVZ4wqx8L8Rx0WCc3RKCks5b4AOUm6Bpb+b8pEWTxhftC8/JsYZr
/AVo2fOSUuQ7+DPwh0v/O69UfJ7eL/DOrF87zD3Gi8L/pCNTS5xskoSZeq5YSNCg69QtKIqAV/f5
K4vYKXZHg4d/Fm4/ukxFghLlpCt3hNM+Ec6Yt7ptmUR4v1kh2CmPwHx3Ngil9qSG6Jf5PGahIneN
g6N7ET6ItKw9X8HY4UFEKFR6Anr+OsWGRT6pXxW43ODC7YGLsVwFALngzpvMBTJheO0btZfyJnkm
G2RBpE8P+FUYxxKKslECGlbbfsWIOMpQvK/MzE5kgx5WOwru5STQxNEfjZRJKZ3U5PfcFGZa2P0f
oRPd2eTM/zJXLlVW1fVotH1QmPa8yLC7kNp8q5pkVY31bwyn4RoDPgbuS+03qOv77EppaPwxKSRc
UgkAqdVnx1K5wkTZ7PvfEp8w7TZOpYWJG0GkVOI9L6SQgoKkOuPQAWEGHV/wAEQT08FsTtA6HLPn
vW4a+Ss/OSdxsfzWp7sNK1Vnro778ti5zHP9wIfxU4s6/FQpx0DPl3kOD/egiKRRa63HHPEmcEG3
3fTiMA/8U3euMSv3yTeb4Xn2U/DBFEdl6MFfFcGBCwQgens1afVpC/Wr+i1+3o35zHG4ZbPqHWeL
L96jwU459hQ1ngpbPI0uoORgU2HoQFBo/KNvJ1o/dboGZWU3ERh7vdVptrIMh6Xa6POjWz3mlbuo
HgCX6Q/D7JSQZ/Gd4vKu7AmmMHzCQZJQ9rdU/LLQLi6ccOVRFLXJi2pkK2nZVbCRiO2YLrhKUijL
Cqcpy1yBQomFDX1I7I65Sl7bulzeRqHxHDNiRn4xC/TASmit6zvL05AbS4TiQMWBjOixF9GpGmRj
X8tBECZRhgKF5O8DMq97ZdqrV7/pIkzssdaUwN8Kq8D4PuJ2Xr4e54PS+sMToezVU2GuXUgGO/gu
mhpAowjSKi4Ltr8yewORcGBCJi3EBb3cOgfTgGvKTg+qJ1LWt1EW1nPPCf+m6Ro/0mkN19g0SABT
O3anD6QlWZYZNmtp+2KJ/IBlATFzzANqvPNQCnxmzun8va4HCVMu1E7Cf2NY7tnZ0aJNlWTWv7z9
latLY1MOBHwB08WZ3bXn0Qo4Ao5S1voJDAU2gus8VoQCQqDRaithCNZOFl7TxW865e4PK9IxN7eZ
C1v8CrNu/WwlKalnglDwPHQ4gMyvTOrVuBcijOPtByCrO65dWYettd6KsZ8gxfEjuJcsEKMTyOyn
+410hlNP6LgE8Oolu9UMO4tQQon7e3PrzHPm4790AA7lVstBvM8+gSFUgqTV/buwP70hcSWaS8sG
LHkWfSGKqPOajjAV3bD2dY8tvyvIcJgORqC1G45+cYLVpaFPkEx9PEOTmHIpVdVlGo1RDHBcPVXi
th+POZFLL4JJnbY0x8qEL9bkk7S3hehMleFGvrfvWKG8DO8ZeDf2L0UBnr/Q3nFKFwrLhgLo5Tuh
AbvgRS6AQNH9938n6Vdn+53KOdwj6MeKb4uU5lAeLg7YnNRC/GbX1zs6eWvESGOyL+dVDBnnVayl
wWqr0VpaQwwEtPP2UZAvg8O0rEosv+RRoV5Quv2E/mQRjnsLrJN5VgXi9+oSIe3IMU8FTJ94TrPm
N6B3ujFoGariFdA75q1K4KZuziYffKLdKyNTPUQ3ol205q1weuGYLr+DPeHrlWbrSuH6AyrUDPm3
Rsy5BpNHeQHvh79Ssnm5G/TvZYUubnba2MCbWPJhShsyqctIhb3ntcDjkfEP0idYq/bfig9Bq8hV
Kep/a1dy6P4wZWW1lxsXPj4UbXDU7J81yvmqZJJfs01eN+Wzo3InxbUj605w0K4iG6jqiCsH1Shz
82luhwrZ5/3Wy1RALvflxT5YLkjoYJ+agxBMz5eZTeS9WUM5Al/n5CA58H9rr1N6nJGaQS9DLMub
h5TxyxKRowKPvfRydhGM0DaN/ZqJfm8T1zREa8nxQ0gtz3QJyIRYFfqbHy0CLRe8CbOgeBGNEsuP
hCC57SKCkns+e/r953SCwgcc0u50SBgQ8KGoTITYDiJTzMXbXbcp6DvTAyWGXMh1OYZ9iLH6lR7j
73ag2gSjcaJ1bh0UAnlcks7oIOCXizCdPL1eKuegNazM4T7xWHjS2YC5PIqRaKv/jSYGoYa1HHzY
iWIxhRZ4xsCv/JbYrG+bBiJcNJ7YTEfXZEk+8nB8RDMrvXaCHZqx63seU6ejazOYSaGTY+enXK+T
0yP/DqsuXmYXXPJVJR1PbVinavHGic/zSLSWFte1C9B6YECducjKMtJmd4a8PqcvCE1gCJCUgn5d
pQSZBgJ0LJO9W/XxyNacO7n07K/SqgJtVHQXmWJgfRxUe5luSz3DNMFTm276izURFke299ntH4Ld
aVTnYWxy6i/lP/vq3qemqA4LIUOrYq9tZq0LhYDGF1pi2+GPTHot7Zgb/W4ZbjcZa+v0Flt1eFgJ
kzgcHQY1f8iUgf9gAuIIC2ZdbGDZzG+7TNqjDsAvEKBrcvvulT9V2s0XAqguNs/UlqcIG5DuEaOk
jHBfC2tTfvKgE1eq+f5YXGcXyfbtsJZxAORXBft9MoufPBB0QAU105BPZh2fBqBywaGykazEFzd9
bZLzHx0NNBSUDGoY3fE7oKuscF1Cn2qX4isEJezJo8NX1b5oiCDvDTCHb/H56q21q+H7xMjqIFV0
PZcGz/tIvCtMewYZ0UgcvARXKjNTD1UN09BoDhFCbqcaKfbLLQ9yyeYPN9TS6BiZVMyaNSZ7Qvph
M5zTwxk3dHWdEl9RPNIXjoGmQmWEKx0HMSY+9GVVOThVih0PUWr18fC0bj1N/flIq0cA+FycmMtW
9n0ArgEw/Y5Y2j8gjTN03ulfPXJP13/Zdti7/sE/70oodbUeAtKgC7DAi5+OwUt2YyYBqJEb4w/B
4qXfrkLSS93OCB+FAaL4/YhBoGSIve09m7/KfJoFeaMKxSQeo6INZLb5VB2ps3HSxj+FYD+KLe/Y
TmmrU/IlRmWXrB4kc03xivm3k7XQs+OiLjiRhHe9uTXU7A1LTONmXUPPp8hOCx5Ld/MJugeCSvl0
5JI11PjE1pKI/n0AoXtgG7LXuUOhoivVbxaAmVFIhlcy4L7yzVai2SfYNcXjtvMCv2TIi0Tdfti9
CEPIOpvV40KCJqMCkrMU7MyC61KsaCSAyfnNnq7g/aaQxe7sEK8MawH1DSCs6vksMRBnKA7zCgsX
LFcOjsQldPBVr7o9HSnG4Il8ZkrDjbL1e4tHGrruqF+18JN/IxTMCAn1Z5vT4J9WMuxj0WT+Occv
BoDhb1FyjxabCGER6eEc7b81jdCpAKC2XVVsttlKSFyEbpjikPQi78/L8/YiUa8+pEJPdr5x0zrG
hMb1iveCsHVkxw9A4V171z+ST8AgS74+FSHeallSr8WAMASwhmK0tGRiKOlq8tXGDE7RNCOZJQ87
zLH3Dmjs860KZ+WHozVK9QMB8u705+SzzKs7gFGtb4C+BePZXhXjY6oFeDYvOwx3o3SGBml1tLal
y+X0l8uDFm+OYWo8mlPZFLREu8MsdSW4B13Tl1k8HfM8iBwF2BgaAV/sEbN3+3e30296+bm5vpQr
mdeLyHBsYxydYFS+kPJD/jV6c67UGEpsD2DN4c9+Yg5dstrXlS8gU9EV/ERMk2AvNKu9TylmURe3
vKu8pMF59/m1ElbUEYqLABBt/fdEuKEDXF1knYz24UQZ5w+7PR7NiBR1lNldEir5aRmbKGKrs/eR
Poof5u7tveHsFMTOr2RxyPCFFYqvNIVngh/8Jml5sMZF8524QII/3tVspNCs2c/MYnxtwREgi8bJ
IWf4C6+jhSlJ7h4ZB+3kbvBdCN5KxfPnt5PCdfQsqJLLFL9indtPRxPEbGXABkPNW3j9GnBLUouQ
uQ0yzFD0/kK9gGChKQ5aeKRVHPXrfHLd1PtgYT0cxpd5TRx2KFgIIM+CA95KSw6tfNNVqf58/N6w
kYo0OSuhqv58DJ6InLwvY6gSHe2YXD2nwbhFUDzrgdw7/THC+7vZ3eyn8GUZnb80vN0ffRQqYR3q
HBcn/kkva95aGp+3k1LWdjPRRc0hCnEtWKKteKVBmpuwzND/1j1fxNzUHkEytbceKLftg7zYaD0w
nvn7dgved3xVBzmPHCP5KsSkGy22JqVA4NU3gG9R47iVltQvj42HOE0AV5Z3tIeyUXHwvt98jiM2
OXMJ+0TGXhUM6/w9PrN5Utz0x2pzRKJg9x+ARQf7jyvY/2Dhb59ww09XJIF1wSqUv0CA9ZZJYS4L
/JHbsvp9blwREnQAdcgtBXXWFhZuJZPkwEQzUcXYWmCD38J3YNqlZGMIl1N9cFCKS1JpBF+RUNB/
EO6eEEusediUOyKL1xc/wbEsX6WPM0A1Vsm5JUpkeIVwNFAZkIfMQRzB9COWia0SLNmWuY5yy4SV
DL64G5j/271fr/ud3nrxLzr2OMyErg7NyDlL3YImO+DRn1CQJpeVe42l/8ESQIH8A+i8tVgUJ1AE
xPTofmE19nuCrbgrQp9ezUjjNBL9Th4YtUuaDJVDGXlQAke69CoYN1YQzU1C3671X47tHCaVEATs
b66480HLneKccBN2UxlWFci5wsOvLimq/g6W/L2b33+QJaa1j3IFLvJpbmAPa4YsxZnen5KJeCDZ
630WhvncIsFTXo2YzL9gc3dH8eU2v5JL92WxN4ILwymDgB0xk2SoVypHzZdWx9f78aahdwfJEJgP
1OQHZaDZeWcTLv0znyelwItRyhTYECyIBBlz52bMjZo/EeTWkAk1iiQ/qOByEPsF0Bg3RU12QAzd
u4cZzf0w5KO71FIaN8aTh8iFw76UI6VGNVnyO4P4ZcpCAz4Yd+1mjEBuCXWReWqRdkLsDr2au6tT
BEXEWpLlWXGheJVC67Kr4fU4LO9YhXhH6fgOtCbjtJHNS8ETnbbXB4djp20dQoZVO8ONVkqzxOb5
FfUA2RM5nflTR52mtmdv0V3PtRqRuRuEqUMJm4M7elRmxg/2AlforMNUFvEeCma40LnKctmWjW0F
mm2PD/RMgXpaGmLu/LLrTj88IiJqoe/KRNyRO8iFG6Rmrtk81+EMOC4+KJoLe1zJ5zy78kAwsHhq
EOt2rgYMzotGO3cWFWo1f0PLdvhHF7DP46W5oxmviPl9Q9wxMTEMDj//IwdLH8hBCBtTih0MBC3X
eS3FjUoYrVhFRPkOP/gcGNhN1IeO4J4zpvwwNRYhB3TMS2EBpdAlEr9ZmmTv2UHuXtE4QByS5vXf
7C8W+SKEiSfhmeVWcJKBe30JczKUyQ0ZAdkJv32exRMk0HNMO1KqYVK7TYQBhES+W9LTX6O8D5Bt
jVb+mXagDy5RrKlSUWjSbsCYcVaPUJlxjrw0lcY0dCCMiSWkBU8Z1ZYo+LSWHLrD6HQTgT8f9lyN
uuuQtw7Vekk9N0cNa0Tyz/fNWEjIUXYCsOoFrZBjQLX+teVH/xQUoZzk+G0S5ubgxvMzUQbg0FIA
XIPauiUNZ1/fQvudZp0k+KohjG34cpYtFJOeGrKkPeFbQ5XcB3HJzRxtyGFey2tY23Yu/Vbluutx
XybIWkaKo+zh87IVgB0K5wsFfemDlVt5u/uEz9o5i1UBHXt1WmxeBLra6cMMr4QoNk5Nmc1MmeoA
aRBi9/eW5ouZYOM0O1aelCzzCS1w2JVjQmV+xXE1IyG1zggRmaAgGSCJ+nyTXOdfJ9Xyh8B8Hkyx
R5vOvJSUPwhL/V6zS1aKqB3WoFO9zLIwl/U8b75T96VHHM/vXNPk+ncpXfx7KKzCwo2CcU42VPNV
L740M1gUMyszsQCPJF/w4MU8S9mKxKrr5G7rJ28P1UIUDPaAJsN2jeSpidvlzSWhibAWRiyGTwMD
A3c0ASoGH+771FLbzli4z/fHFl2r0Wi+0aTiQHleK+1NXMnRZx+t92HVyCRsTTNmajtAP8aQ6MsO
8oY1e1G/T9J0yRv7e4uZo8d7pB6fniKa54c2kweYM/EDfyK/0iRt622wrncmtTZfThfJf5uh5eAV
5j6PZTsBag9ZGmPh4U//RMtPHFbo4ubkhp2oiguFX8DFhqLXXCm46cPyU/fQ8Vt3WqYmoKuYaPt7
PhoR33nW9cnB4jAoBQwDl7lnH9G7MW1SEYbWKfONVKpXGSCrSojAzwHfLX98TFPmtRkLBoBCh+Am
peYhyobaVGhV4fcXauPORO/lcnmFcTklsaLDL6rE3lLpwMWUXmUBbqjlyocm7QFJRfd0rAUo7S6G
WBPBE5vP9hrWC76LKervN8yFNo2DDKBkbJaRHcSR8OopI1AaPGPnoynFRU2LvPm5Q45j/SMurZfc
cR0vefEt/Lgk4XAFIC0F+Iz+1baj8Teu+yyLE9BzXnbM/tnquVKTYKdCo3Ig0ONpqrcjUUNruSvT
M76EmcdWgdy4BpiQyTe8n813EFdQZbbg4TxZ/cdKRvl3ETxHC883UfzRSFZUojgFICXeDZO/O4Yq
Q96sey1VfTu+4l7wiF5LF6HG39MoorZbv1hIiDMSEhQBB4N9OY71lCuImOkO8bxdGdZYotkSTXvG
qeZfwxlX2nAfBypdMEdzI3bGhxHxQdcE35lEwOKoyzvG+SJz/2HCQuXJFs0rQG0dAHN1e3UNJES3
fdRrXPaDVv4Dt1B3F/Gm/4i0rDu7lHBkvaQaVkfoxH5F4VtOWjNJc4zkl8AAiDtJP7JRB0+Dmi6Y
qs9xfnYq7Z5r1f00YoTlcBygmx/c147fHNRR1fx4fpuWTSEIjskefb5AjAJxwwGifysGrylG/kfh
pYQQcWGN1gK6tmyxiObvWAwi22EmKWScv1sFzkYwaD5JHYvPRAvcIS96vZVyyFpDbtI15TVI/ohk
ev2xjXn/qg/uAUu24OevfP4qcFARURJcw7jiyhJLu0jxYt7z6Zq3CtoR9u8ti6eD+9H1SBkOoVQZ
rwviCG+n26duByspQE0p19n5fRsvkS9pltHpCGVVciUwSvh8rgtwRaEKTsGqNr8BA69yK/E1xH5Y
P2bYE2QhV0kEVy8RATRCJwroa66Qk53CmgqBkgdi3klUnIIgCJtC9AlJwaSKSfUJaZYHkTCzIyZ8
9wMm+AwTwZKjs6XHg+Td32v/Xui+a4ads0szBnblLvQ+kkycQPuUa4qIApQ2uiRNq6Nj1xcTwGbB
kFzykIEvc2yNUMeBKl4aKztgYd3mufhGOM/XnQIx27JEOy5CfPc6+otLi5YSQdkeRptKiKuzXa2S
RbmjzswU/rwCFIAc1pvJvVtS+obU+viChtMcsCXK4i23UfL6M47t1K6+3O7dkZiqTAsl/E9QAoWu
B5KpzeO+dpSw99GxavQEVkbjNr3Co8AN6zSMnrDrS4nCTLqE5mJp89KKhVcMfE1XsgiFglFgdJcp
N/JwgXuPALJlCaskuHHDWLtqn3uxybzAC4GG3CfiosPvhZl7iUaFahOrpyUsyD+XrB6ueiLPl818
J6NkCAM+vW/2TCz8eLkDBpgVxoa/5gngsNM7Pi2TM1Ht1e46Cg9hKWAOoLvERTCpSdGgWQAkpEri
QiXlqR6y+dTQo0eD2lagS8RvdBlAfk8rbSWygL+EEIO3ZEn5fDcNG+SNhJSAlxSPArTe6LZ67WXK
Tt5mi6C/o/2J6P8gDWhFNmI2E1v2CJrfCCzk6noY71mYI4aIS/15kwHzZ2jiAo9clfIoFZv96nMj
FglHYZWdvArRmLPlE1uAjs+bKKvCDGGr0ifWkREMVIHSJ0JfKIevJccXQRsQjiHldQ4J/7rgOEz5
h2U3D4YWbWzbZQQ3/3o1JDCf2iCUj/dipfE5I6OPrz+Jp5aVn0Wf+9UA/8IZlPkvp26zzMzmerCX
xQ+Qa8vVwTNbgagQDJIKmZWdYzi+6QAfTJ5TnM64rQnvYGqK305GRnr5IN7BiezROlNZbCYVS6qs
YZF4pE4G/bqElCcGHOvDc3UkNF9CvzBfdXQUZSf+OPSx6KZD2tyMEYHlyEijNJ8D0LBjcaFqcWsu
dmtFf1rUx0VGHjlvUFHYCcRz17/5aTSYsp8jOoFO8y5QfuAbwQnTsf6x9MTGOkP02d9yNhHu7DF4
luBYCQhqDF8iQqIzra9Kq5O2F8k3W6f4OmikRQpMYOad6DBpe5Oe8ccuj79XYySKCbk9dRCRw/rz
xPAAeme9yPnTSoJDDvcSEXdQ3GP0JHS9mM0Lw7hKfT2wDZVm3NSqCta2JiWPTWUPEN12zmGNd6F5
kemPmc+FgKxbjQnaNVk1JO3fqT4FJcnJVpIIv1eLKy+u5DoDIXSfH1mVAMNe4YKml+CGL3guS4IS
lxn6Ia8VZaycSvgoaLkD1qnwg26NoCXQOVQajd67Ez1yM+dsr8/blhQETJLwMx11B4Q9HdDI++CR
kvOj0Mup5w4iCEsbQuFrP5AzyoZOfm5jSrLnR0+2e7ORlJ2J0EdlVuOXiH+7Vhzx9dKxFdpvB6c+
PuE16anuJHmKNZE+QOh+W3IRns9n3eaEgqKjx1sQbRTtmz3c9NZmU691AoPhWE9X0tNBEpFPy3lT
2v/sbqEInjSop25kcGFrNC+ztYN0Yg5dhcj1+bWrv6eXFtaInbkGGiHZEVczWKZQ2zQND6bjb+8a
hs66x4fx4bpIFIzp8UIZYX4dA5j6/mPNhQeb5RLKvaURkVhGpGatpxmsPL8iuJvkvgOmFvWYlLOn
XJUPUKGFoQ/SRaV1/3JqzBNgO1QyhTzRt+V/8aBQe478vIZDIboU/ahWZh7dq+Fl6fcZG1tlJIO+
1h7UNPBVdPyG5+w5J2fa1LwRV/6Gybon5MeXfvnDpO/mQIf7DGYJvKs6FOMUbytZCXJZ3yuIAH/t
ndvtu3Wz6Kdw98IjKQJqIw1cGQUYdhC4pxryoCufmt+ThZG3os4qRh3pn6I/pk0/Uy5gMK+t58Pw
Gb3dmOHxtgZYfI9nesJFaLaCudgaqTX5l3sA/DejohqhmYw15CFcCrS/z18wBCTPivfWClxLNJn/
sVOdGK5/PX86eDjFub63Lm6v9DOGhk0GLaEQJUkmMa+8wakwWMnkQda8lBwPabNy6is9a8SXtJMe
YB0CrF4y3VIroWlXoRqlZX62kTXAITDftet4rNjodOKFPyIEshbQUG5VSZ0ZBv99eEGu6K40RrW2
PS0KnkYJLxltWxZxysnH0erwsnqdahEi7YexGlS0QekJ3lrKeCi+3hk8j3/6VE4D1E0i7eowkm6V
dCGtbK7wW3RZuIyKr6QVbFYY1ZlkR/8OkQeFebuYx9njLSFCX0xTDMu1KWqBuKlj5+aJJXMHeOD4
7GLVYWf5jC0M2ad2ubhyto8YAb4d8H5gEz0o1F4H4irPlpwY2CbZJH/QEkb4eVvqi08s6GGTsi93
hoKmN4Fh23LBo6w8fE258RVDMe+vd/xxMeucMkU3+sU7dFzXSleDp1uWdybUUtYkspG5vj6z+yZe
R8Z4wedNaPgDKMgARMTkgglkb5YNozZdKkxRfZSBTwl4r4I0d5hd5p4JBLlc7dMCWPYuIYkdTXSs
3o+SOxr/+zNEYKh/FdOLl1ZrDoq3WwZA3pCLw23wcuin79Gk+RSeqgnxFfRDvD56eGc+lczICrPw
VGX20NPjYuxbX/fEcmPNxsvAP47vl+96TZErNOe1y4zpNiKYenRKKXYhNjYChNaxUvxAWrSUugfE
f9kNY9rqUJG0TfS+QGhQm3Zduw+W09xfp941wj/tZjz4bRSy1aSIbaSoyx3sMDkrCvWHHc/rP7ag
4C6htOUeeBnvPvXP/eGO4YetB0S/dhlisxordx6Pf1f+KhdETkD0A5jFGcdMbUHlbJKLzApjndkJ
AtCySUcuFn23qK7y7Wyr8RS1do+qVvmmUmBU4yjTRtwvn0M2kJOcLdcWZ/lSK+fWIqPR79zpcTIe
v/i0MqU8En6pefHLvvs31zHvTKM17JQHJA/nZUEp79fSeGIfhw2BWoQqaFmX7NFvzUwCUHgFt7Uc
kIfma4NveJPuARcN3/C8B703mdATIIsopbH+nSdRffGHscVIqvjzKCYW4nKbWeGVy+wnuCGiDqaU
e0Uov4lFXbxu6ohYl3VXxwT6k5VKzv5WyeJGBvWjIyhmh8sWDzUNtyUtpKGEbTN6+nzyORcSZinj
gsaxpCntlJotc+1lj+BVi9TxWtUR+byRq8/FBQQJ7r3StwoHu/FmltIsfaPbSfuz/eB5tCKWyCJl
dvhQ+eiGSjNtxYF3Cl38+RXBB7/rD6oOIXb83tp1mugNV1S0fvohPBNsXWN5Aa6TLmtmMCR9fqmd
cD/i0DES7vRTu+iHkBPLphy4XbfFRP0rG1SvG2THKI6BmZ4Gfkui1AsX5vUCR4VoWLfiD9uREQoI
uL4GgImWBWzyebj43Oaw93+M6zkkb3xNyzP77Bv608Zl0oEv30BGK3gUgmkO6xdyZnsEv7FwkYrf
EuAAI7kj+2FT86uzTf2UewVro7nYK8tmplDKbCgiFgeLye5xL7Jou/yALLjjWHEAU3YpdPl3AuGp
iZ3RPl0F56IYZJkWKy/9QG9wW0T6BLoFA5juutcZyAF0MbfEGo80Xxp5bdlzITB9smIdJD95+qRC
0XE4L/UkZJFKD0n4M53Ysc92PqqexB95ShOXcCF/SQpuAQNApm8m03h3VyG6/aX2kYoyuV6f00Ed
rUzCEl+Sc1uewHxDF5D2IFpoPcTzGLPa34KjV7cfOstos7aXnzlWaopBy4rBTimc/ygYAR+tH/8X
vzHnbubBY5ES+xyZuB1TBqQl17O+SeCCc34ef9a2N7jxOeJrEmV1ZU6oZVV/zTBzkv2caVIVVCpl
NO4KyzZ2E+ylrDiqWf6nt3WaWRRAkWazci0VsDHzG6hvAXf7v6s43UQ/hEenVZPzklaRTeGm0fkI
QccBVuUo05FNGMy0ox4Nyy7Dh3C5D7kvZwORNA++54Co489ZDx0RpvlECNa+7cj3xPAsVaNzYdlI
tnum7l/TbC0bDw3XlPW2RXtR+O1q8rF0rpHwrafHqzUiCPA8ei96jnzuBkYYN0GFoPMgnozgsuP6
DHWZj6EUgU3xjzBkxJo0EYOKjzpJ6C3Kql8zDJSe1xLmvausmMoMB8sFwEjRaSM/T9N7dot7DneN
RfXHAfVO4UVwsBOiUAatbQnj+j5BVktaOH7C79Kkj4xmnQsEnaCkNJfSyoPdRw0B9Cs8XpaXUewX
WHmGoUj09tdPmIDcV/6MGL4RD4PWxEgvvbJp/r/VKSQRl3xgLqxA/gC/1hP4bGGqahOUjFOBLGqO
L9LX1j6H6SxNYZ9UXQ4kwIAVuTr8yzL83n0Uoc/sx1EGJ9obs+T4sZpMIb24YxV96TWQcNLy51Fd
aSZTovR/tJHijTtVw3OkUfCRAvmq092QPjOl/1wkPQPDSutJX933FwVKeyWpEQW4re9N+ySSma1v
ISvKa47nKr2lQGXNpwTIP7P6f8gtIj3UNlkJChwslV1HCim+HITDOJtjZAfmGesjhPi20qZLJ7h/
gNLQ3w3c2TZFfn/69M0ubjqUAw32f5ep6HGMNkMmpmGSq77s7NWb9MfxjMHBPklaj2S4swRMAVSE
QTtCmZCRpoOKMu76g+6xEGKXpQ9uoIoIXO5uPQa1mKhYo3pGlb2tUnuJP9FrecP43UuyrJGY79pt
574plhuOngCu9TH6ISxxGbQAATsBMq1d9cOdhBUq7eLiYSxwJDBBYFNWEG6Xw0dOuSdRCJg/fx/+
p0I/sSWK5mkA91WYeApj4ifiy/GJtxATsJnIwaemW3FrucpKgmbNv7VIqtcJ6SZmoUmhYvFIUMPq
IFMeRiSVu37+k7DU+E9InOjaoN0CdoRXGqrskH59pphqa6cODI6ZcAmrr92yO8vKbEeFZdDi3oFK
BzJi6XLt/w2CskZtjbjZ86zEPc7LRF/Xwz9BTsTCmHpPkTTZRLFCrANE+4SNrafljcAXHq06AjXx
yGuDwqhGRH347NeBX9lzfshVQXJuzXtKCvcNQUkxn9FsZxrbcs0Su3THvSNiBwlvjs8LJupKLgNg
1qZc2h2jGsn2m0fE5QEoZozRxkEZUEdw5D7Z3fox4ChNF7LIfng9b4r2wvCHZobs4z2p75lMsvRT
19a23KUCeD02jOtAFJUh9ar+FRIqlkPN4P3J5WsfJRe49aVn5A/4/hDCYawZmk0d6bkHQtVFAETm
l/niRLP6ufOXAoo/UQAcv/DaKwxVrT+w8bp00pymRBkQgHrrNHw2Db79WQ/zGMhKoMTN93X5KIoq
EaGq4iUUz3gh/DzfKNnvm+yiNDwpxMfvLvUMS5A0bd3l/RtJAjCxlYcOgGAHyxOuBfDKTOAHwZJK
K5YbK1s0Wn82ImumVFdW2hWsgjpYcqFOFC2eLzgXKlSMLYaZ5GdKt4RC3RiHesjGdC7fadOsfwVB
ihFLYTrWL54p37l8FxF0iByAjm6IchYOSklfdGZkwThki9q630fcofIwEvgoGVIz4RtwOBS4PZzu
8mFJ5T364zA1+bHmTWOCy7UrD4Qsxc89H8DNMD5JPV7QXBN7K+PeQ2TSCt9UjpochowM94Z5l58q
CBqtwG9HfnPDiJGacFKOltLt2A7JsdGSZRopNm0Chh0Ij4SGA56n6mRGh9QmclKLYEOkWB5yaGqC
HWV6pM4uY7koyN/fFayPMLxbSQ67t0OcCfbBf8nuHCrPM5kHHk0ccquz6/fz97rOG/UFZWW9/Drj
0tbfrfF4yp738qYS7BOOp/uhgx87srq/+KB+DB6Wv1xlnFYn4/NhWdVo4nq/8DWaklsJ0JHQg3Fe
8HH+dcIx4MCzDMnxRS4hcjaDG1VOHtpzpxPytd+pjonUoAwCm1ysmG5WNzl1PGYYYW4du15sco0G
BEDRUJKtQ4XwYFiw7/tYYVFIFZeE6eRAnNikiAK4i9sBS9XQ2ZFaNtU0lFg8jr/w3yV8IIazN8BM
Rz3VgwCCWVMW+DJs45Ek5/4/ORnOOBFSMDT58vAS4PgJXzUkqx5OKjkh3R/rxckvN2IgxPyA8gma
LkHo5BI6sj7XRhvb6fTqRD0Ex68mAUsiFoCgQf1iQ1iwR27+nHsYHw39gKiHrlaO+Fqb3bu0Thib
wCv9+r9bhbjzm/BKExobZDL9q+MIZTrYpaSLkPEaTrykTOTFBzIUF7ZjFBcqBK76bWsbd+rX+MtG
db4AUWU7dBlvAFMku4XMifS3LmFvMcg1j3mFtSXwr3IPY4UWOkX0vbO/nhbRZoerorg6lc/oIMfM
ALQSa3VTjBqIeAwQLRYAdrZwwNd53BYzKRNwx45mqKY8MxntBtXhGZYyaHX+Y6W9CnhLNOXnFqiG
Jai6acr3DJq2zZk0IPGqSjupBoWxxujyKWcNq9HGldu+Unod9QxBLm7oJYLy5Jr+rxCQpt49EUhq
wa6STF0ssGN23AvmRqm+Y4kXJ4vcbAjc09mCfvcbdCk5aBZJI/Rq/Xk8GgcP8ZU+Jf2Vrv8F6CSh
6ZrwYw3+c9gxYoecMwcPanCwGKsg3BSiprITyyk6Al8ipKrb2q9srO8awLTRpv4txW6kH9qsHT3k
iJNvwPkr78IJ1264Pj2QhEB8hRxdbDOhAsBnDqXvYHTKKI6oFI2lJTbvptqZRo5kVfhtJNycfu0c
I478o1yjhd6EOzYry0flQRmNeKP3uXyZ8oH3wI81KDqR06JMmb6KxnSY6bayO91/SquHp+LtpB9S
aapUEWgXHhC/m4IJK+dmuYLiLHdDBrCeTa3iAV13jpAW9wggiHvrj0b2l/ZYNMENbLjb1HhkhlPa
skpzf7DyMOq2usx6CW44pEefazWX4VyGRLO4WgEbkRHtn4PCm6c14TLs4qK623hJYAmxD7hvNR4u
BoHa364spyijHZ3jDaO/um1+NHZPBgQu7Uwy2WW5IFoW25A+FQ5Vxm09ftNsmSJdmObXDvvkp6IZ
gdDBlaRWYc+IHNT4PSO08PHcqNpHIiHiDVRjnk4rjZ4857Hqk2lxzDzWoKYmUOdtzTmrkhP/LR2x
OwKIHao/XUMTmRq7ZdoM4FBDP0fi47QEZoHssqshznav4iUmsxYJrb2XsSyYDyMI9T/XcIPoMIln
aheR/iF8tE2cPqPNDtWOlLwl/utJBqA6rFBptum9Qi757jgxdzExzqHE3HD7LLzjmJoGUdWwtZdK
tFlwDOjrjE1AxC5dqcicxaSG8JGC2+ajpwJdZVqkuiQTHZN5BB3WWBFGCTwcChcsAy0SW5ErZd6X
p185s2gDRLJhnKa/sorQBFPLQqC3vi9YcnGROQtRzLxJnVum36UmHfgjBmHuKpH+fRCwnuX57ydp
baqypqTATZ8iLoxda5V4MskzJnqNnCJBWHwMTJjzyMt2KfT+LSSWq6IOIarjCQjQBjZZ78qyhAFC
VqniDOoTVsJh9lryzmVciYr3eMPVCq/V+bMogklXW3HVmaWvU7XOOMoZec6tmHOcpDE0HvQghUwF
ikaFRYajMXy1YvXDs8Zzl5stulsv6rnXITqKml2r/L4D60x8lUs68ryuwnB5GDmNjIn0rFb9P7k2
s/Os3BSvKRDhk/OJjo3LbV/8XWFHkjFi7IyqKJC6P/4RR6ivt2lf5Lk+x5X34pog5sSmBvyWMkhr
MQIKGyHLTgZs10I0JMCVbzuUWpf67kwrYNCyWthWsPvpa8Di85fNnwMtNWFuwkRMvbFwiuwRzgqy
9OascYkfm+46gHe3o3jJocSx4KvVrH34yQsCn3t3bh8+3TX5d8i3M1azeU//th8xa3Zk4mzW4Z/l
NtmOf1fRw6KOrrpPBoEKonMMzH4J/aF8GgBsaxdYeVzd+nneop1Jhy0kbisO5HFkLUiiNhR2x/so
acHEgGQ4ZfGTr2XtujOnUdLbtqfTvHsXiorEwlFh3S07N7cK3+KhRwagq6+0V3PSBZLnHiCTSZ4/
Dh/RsJxtR3Ra0Ca0+o23cTyXIHFZ1RzoQoBqzS2pD3hEd81/iWK9VHVA931Nc5xz/dKGQOnnONut
bdhSJIspVc5uETi+ZESOZtaWhcDI8xxqK9bpyybEmRjPrNm1KGDiNopOkArJRHk41Hx1nBbNAp6L
g0mBzXc4xjWC228FjeRu5EhEV6CqR2/nuLytSaSptznBvOFi1FgHtBIZMk5V9UAZcpzXyAzANGN5
TMoGwKA/C5vFjAc+qxotEOMZxCuXTSz1SlntczakVh+PjbFEODgWUyczNt7qRRbX7zm3TrPRV1wg
C3hX7M9HCwGWLEeXVKow+Uauqq8orUn3l9+rBmxPMX2P86dgsypuh/Is2nBiT84T6BgxBKm7ZjtM
UWIjluJ22euwSIiWdGLW/amgp3NL7PP6kg3GTLiQvw3PCwz7Aabobjcm/KNcuigY28K76kOeRcKl
LD2YLb0xK997dw3IhulLtTwMLqFVEE63zp0o6pLtMsucNcnE5d5oTkkngYrbUl9hbxAxeYrMuUjB
INGWsNNTQ4FdVIIz8HXDMcqHIZHxttEC7pm+RZbpEeDHdsNPJqvQuLyPghzoxgbTsCL/InpTFk0z
gAadOwHtxBP47DqYUCgy9REzCKWLHU4WOvA/cE8nFdp9LTQligZOxl5bgD+bNrb8KTMfR/SGA3JO
VqCW5X0FBDg0w5M1wCfSUg/imRHiwLnWisenZT00Nz4QoDJSWJbI8WXt8HBmKEgqjmjy7KRNeQVO
RRy4GFBiNF4AtzC6JAe6fl7IvKhsW6ijqNMBlFidLpyTOLGr50wXyN//6wXf3uF0L+4rIwf6VXpr
91SxAZapTXy9F6BW+VJl7WWnvCIFdzZRxl+mvnkFNKPOlUznUEmYhclwj18Ocl5vjm1lLht+g96q
nhrkWkOc+rwISjIm3Gq5W2lanWJkmHtbmPBTtR4NRE0TPC5Wuih7Jtp+Y+wAEQ+9b069JvIhFy/K
hjnJzVi1vVOuAg0+enQErAe4OC/tLkNZqLFjK8xG5BkWt6OjUQBLXtSvKnZqblpIKptzEr//M+ku
iIifXORAzfPvdR/fKL/2V/3gJJB+AYuVsNDKjHnkPMzqyWV9iMgD2p0zcRqOrnhxtCFzNrrN6ccl
/f9OhXIzI7/8J/vMJLmRq4XKkG6IkXSqirAGYUf9VP5ibHOMybncaatSPYpj/3Yxe9cK9hZehNlU
b3nQ6hFjFxrpjqAUv2sWdMlOdTYx4X3O6faiSjlVb2sOZcU82QRzFqAq7PPsiF4a+4Z2cz6XjIEt
jUJlNufuSIox4w7Em5OHNH6Enp4AfHjVDP+rJvQaC/d9WmOlzTe0H2yVYmPzCj6+cPZkfLtlPL8s
k24fCGBnNB8feIhvdV8IP+zYAFl7ugp1JrhG6pfPq9P2lRcQb+xcyTWbn5B3TH4yytJ97R0u/Xl/
dUJo7Af3IVoLCQ31lZSFj6uiwylLErpHDH803BILV7DuMQch6s2Q55dM5tPKE0GT8bedl2vCap25
ayadDF3pOaO1BaZYfHq2hG51JbEgG/G90cb9qoY+aTzNqx4rDqSAtfwmjdKWq50rH644RFEjyX/J
3NRjc3OzfF5cuXideZ6YcytEDBwLZXiUSm4LcmraEevC43ye8OYquv0xp1ZKocjMD7o4zYJKUZTk
z4/z+jZpQ74eRgIfN1PoQssSqw7JFuJ5CqkeD5dTolPMRu5JXBfuCuUrdDELc+34foA83yBKyprk
Y6KBLaHCAUnPPPUHbvr8FpBDl5ktu2ymqEBEvv6KWQWOuHXPCXESEsCchpicPseRWeeFhW/etD8X
5Pt96bjwaLw7RXBJ1NgqY0XJ5bKAX8v0sI/UV4dXIdsXmLB75IoF2bS0h4UQPdCSi6XtniOHLFQA
InUNKGquvpG7/xD2YA651M6r+A5DSFW+Kw6a+4DYS/aira484FBu/u8HWwr4waBUoOwyLpsnvjsu
QLwutWd/3926YQQHRr4sKMsLLJjl2oIkxa42UgJthY/tfQeqe25XMiHeMMBB7Nx5696JJTDaFedm
4Bs4hsljdLYi8pNiI6SB0f2U8aRMskYnVljkUjx7EZQyCioHmknyDV0WMwZplX7E9pM3kh27sZjP
AJwza5wGtsCPfXAkn84lyqCj/qCwDPQ8m5S8futwOriN96Ag6M1mjARcLjFBH03/q81t73woG7lH
fPABhL5G2G+hisrXVwe5yB4fFO9aifUMgVKZhzhEKjGQHOVnWvS18urUSPMER9AD4hbhMbPTdxkA
VOfNOZBc+qJWga0fh2DAO+9IY3jbrLr5xzkXXwnGNitWdXaZK0UQldTeRoMq62B3YvNs7WXhC4+Z
ZaNaXQ+9atYk1b8nJCBW/4/7LXLgcgs03AFiWARC0AgmxbhMUkcpBbTuus69viW3hRaiR5xq83pB
lFf2iqjm967puVol/rExNKaSDS0rHn/y38OyHksaCBEkxlB65xZ8DGjgg2JMSH/61DXcYjiXfI21
95iOnQgRJmWic+lvMBLGrVofhGfXvRKnPNi30ifbktTGR3Ad12XxiRAQXq6m/v6hFhdO7W4B/zSr
6jk5zY6Tur646GktQNL9/ZJEpuyfps7JVO1rQEzFCYeQX039yvfmXYNPZXfGdAD/j61zfZ3rm3uz
Rv641fFFaxCIVsAwztLVwrARJKKyi4F+keVeYB/0+CTGbsNhOenJ7AKojnDrFV3VNF6O4BcoI0W7
pezx7wKCyYtQ5NkdJC8IupUEl5zz4IGcIfok0f787NS3ZSBLZxCOcBTxAL4EwuT3tFnxxMttU1il
TfeCzP2bWu45torKcbvFAihSLL5WlYtc0yvBS3MLSJWZVkwrVZ3cETPdyUcdWMGcyAManC/aS39o
/I/nntO6RACNRHvk1dAMF90qDU+L0lED030EBquZzFvNEUWW2Ogvk3oTqReqIX89wl00AvWzSx0X
JFNCiUgWdUTxieLubONlaAWGwK7uMH1Z0Uu8FTlv0OJaJb1WtFOA2m7Plojk2mlQ56T3ry+6VrgC
PeDyCbQJba/MF0dGNcYzAZd5Lv9cqmTYeJUf2hxDIoT+TNgHoWncIJ8ksgZaEkgtddARohB8RNvV
C3vcP+3tN+p7+SKMizGsu9ZDquotLjtf8QZ5cAEsN7GM8uYWj8XuDfRyv/HNJ+ebveaMA1YzDUUN
7O19wxSTFsGfEFIo/Svr1jLtkDcY25GgmX/dGIsKE85DWhAj5AONxDtSMqrH+YvDheGs14aoS4dc
t0iwzsADkEb9nbGnfeV4iJtKCGzBX0VSZVZApJAnoyJ9PWp0lQ7C6FRx3/OYwyEsd0uxkMnL+ZAG
gz8+mO5PYGUg61ZoRFRzHCyJoNpU4EqVXGdAktxyeiV9rTmTiv5vcFzu4fZD/mPePpIfJtCZxc4w
ONOILrHEPaRxic2JGt3fsIW5tDmw95u1FXmxG83D3cnlzuzR9PN8V+DLpOOQER5kdRmW2v4yS63V
VDW+N4Hnvxxzkqo/9uQwo8XHNapTlTYMhguCfE55TyVskAktjUmlCK9fNPmh6uPWgZWgEVAC+tt+
5/+abIGyw3hzX3gqM2YFFpXfe2d+0BSd5FiWE3wzEInGSDj7Klvf0xQR5VnPhfljXNsawLR8hQw1
YK00j2S0vS5KyAye9KxKGMCsQZC6ILhwYGdXxUAk3POEtjck021EUSpLQrfzhWaPX+sYgh955GvY
uTJEkd53peHA3OCOj+5lPDqNu8x+M14uT0eLqO+rW1mDbUNWFMcJTOcPGdWzd6dJ4jw2kX0Py9gk
+mUy96BFG1UiSFvp05Yc7C8tcSlQDCT5Aymk104piGWkOZiZAMVWau/y4B4zf64eda0U07H5eR9Z
z6wmTnQGHzY1Sc4fkwgyQH76wFGwaAxpup/ZCJyRhz5NSglQa/ycNEDF2vJQLS7zJGugE0iRSof/
UGKRyr5MP5z1FLlxMyaPzdJH4fuk6ocET4Nz9XAv8ASGxI1PaH+9tB9m91F4rCIEAMbtiNnp65ZC
PhUj1iQsQMfOL88DI78hRQzP9n5ONQi8OFY65cmZ7ssdEcPLAfqE6cwReXkL3ZutpDJxcCdxOdL9
gRB3mqqzmGKbp7WorkbyE8fEQ/2ykUqw+GQPWF/J+QX7XtEF8mbD3/iUiw5swaCzIuotIe0gDYdi
bkupL4qpKix7z0z6QY2I/Tqx0i8qBeAaeClsi0SjRftR7PdWi8bdig5X9gDlNl2rMIke9w4ZJ0Zc
AdmLvin9e2xXaMg9LHdZDwQ+80FQKkUV9omP9T6uPiCSOc59Vr93/xivLbZe6krszLai+AIzprLj
Gfdz4hcFSMf8haUHh+KbfBa2PowsnASu71UB30MLcDnIs9UtnZMej3XZbnXoqRv89d09nTUwOyPF
6EsZBN6EHpR1/77oY4+3L/uyQEh2eFbbifDImHY43tR8gGjjpV6YlucHnXGoiIcSeg6+uZ929jAl
slXNP81K1HKqF6TwC60XHLuE5TfEAWgrlY0/FQRaq8Q79W9LjtsGAK6d2uBzdSfqVclxoHmg2SVu
YovswA+nz14eJabGC+/Jnlk1Hpmwf1eS9Ztc/nFnIDUQjeTmeBP7pGo4Sa+Fj8qelPOEYxLg94/Y
hiG9o/LIE3ED1h0mIWPkA30wxxTrNhcBfmuzLIlcMzG7F+cr94SPWJsNlMNiEZzxyiMsBrwhTf91
LVXmXgz2YwQxbVsYIUKQiJMDig37R3yMbngHSKMX4i+JM4LCvulmtx8/F3+LEakW2aItZqxO8ODK
3+03pFWNj0RHnfVro+tHvE77oGqEYZ6VRFOF7OJuZCFSjHUdPjmkno1UiawbOFLMkRHlDnzuNLvv
4dVcltfFgkFEYqgZ8vxyhZfcYWmfLSTIHajAFKXBRvp5rT3zybjlRaw3ijM/B2Gnk2BmVIncMLQJ
xuKFMAapV8rlQW3oIiwLz1XhE+s7JrrT/WYlLDnhbsV+SnE0T/pUoucQ/vI+puMgv/RNvYX4hFh3
TBVmTJq1Tsr30Yw0LLI+UR2aDv1Wk+Sp1PTTheYdjnVRkXVZMuQgjvsjeuXPQFKE3zyUKU8ZxEVd
vCO88ywY/SVx/MIqQlsIu+6IynCis6fhHkJcsxXjgAXgRq+MYoYk7w7vAvrKQaB3lFkEgg4trXZR
tjjYWT1WglUL2Pkgco9PPJLjGn070XA3s1e28n6Uahj/OS3uu4GTrzz+1fXxrL5bU/LnxhQivURJ
2yELL6nPI6dsV2uzRr4JxTM17wJPuLN2Jw18Tqp0hEGE8pMZNTAYpvfuQs9U71Y1fCzMD1U2/9WV
U8AsHnrfQKYSiKbftMKs44JXgoa1VLhJm8Pdsz3D/NHiel56PuTKdDTM3QJ1fkzcucg6bF2Lz8Es
5M5IQrcZWc5KbYiHskYNsDVWxjwcqgtZrN3cVbwCFE5feBkleyn430+vh2IC2Cr+D/wWkyytnT1k
xGq1oZdkbhRBPBftI/nQ48gWASnpqe+52dNpXBJlqGele+M8Xx7DVDj6pwruGGbq8kn0yIJ5lHUR
EQhOc4fwogFgd6WCndg/EKwWol3mX3C+kTIIdBwwNzCeLWMqS6Dx8JboZwyMWdJb2+6eHijRUfrr
ENsLI2ftHPwTCGmpqPi8G1hG+e7lrUDcVxIiKQKpKBeC0ouNEdjW6AwhLpZckZcsu5ucI1Y8ObuR
V6wZWOQayGGWO+A/boC2guzc3t/QcaVQpOSVVvTqYhppVx9OI1nY3SrA/r4kk8ANS2uj+gg35Z5j
xWCMHBsidI6dFunTfCowjdNrzBzA2LSPZvQOtGFSHUMgFSWl0t0IXVaYIb9+ZsuZsK+dhY3yS+bW
GSntOEDJgJW5KcFy+bSRQaqlY9mnxiloqoM6IIaHOqrKRFFNiidyxSh2EWJlFSrjpi+YjB6egJYd
6tPMVO3nyv8bw0nQqfFlkfTrVpLoTOutgbXhdXo93N4xYfamIyZgF3ddbvho9PxfiIy5N7gU4ajx
flz5zfFK0oGcfLQr8BAUdAtIAb+FKZLtUQTeLGTTAr1QBx1+kFbPULrnJS5eFKwzovIFJHls+F0u
hEGHdJvahRrq6aQr9gnr7MrUHfsrgJ57nKU3h0zGVp3SdyYHjmqfVFxLiCMltS5t7T9diKp3lDS+
RYN0f4SmdGG4BMGqtsUQEDtfqlnd2kcrz99rw4k2RQrC+mDJrDvw8n9ImY1tIqFSGyDUvy+lyl3K
B0YFU/feBIXo2oIybJ6I9n3SBULzWA4qELUOiwK7IosXIFlaVQ9fMhzAlhoxdix6Ie7Pfx7BHNPp
12grtxeczvVCSE/yhEgXsuLwOWHbMbtzyNvX0FAbv4o7rXHk7FVb12VYKv8QEOYDh9rN8kQ828kB
fjrBbgcwimvnJk40ZZkrbAcdStNfIZ8ThcfeD9KYFB25YDo4mYCqt6rceyZcJDvN8y5nZQd4K0rF
Qz4ZtBJXXm1MYus+G3aZxzTVCXX1kb+KP2IrkZmJTUrdUW7vg8sV34vTQYkJw7tKscz2BdVYC3HX
eIAi9t0DF5ggOjsxDCS58Nlmy0sJmH8b3XyObfSi1W/rBa2ec3vAhiYe/MuezeVrD/NlWEQXBiiP
isBRx5PscPbs1Y27cYka5kdVKYQnRhiAfIoFnOpQJbLnwq61QTMwzGCB9HqLwfcKdhXZ1VdCQWlY
mk2ozQbC2DxWqnPOiba8LxJZuF40U0kP1LToHzgJ3pAHswhcnv8JegjdTJHI8MO4Q+ID2qLkDdqm
NaV/mMb6wnlbl/nn0GT0A9uFsKvQDKW1Mf0wWT5G6Oiy1mnMg5OFNmb/mqoU4e2MGfUI6Y6v06wC
/JaPhZRokf6jHuYn+pc1Exi2Fdl/XR/Ldy6ZvK8tRMu6j23oFxr/B+owXE1tRsWQxNU0JnoXsNAn
7xdklupXsUIn+pAv9jWDLtq67lv3Nwz9Q+vn8J43xc2efIrbVR88Dzu6eRgKNhTtAQ0QeJITs50P
nbRpEBIdAuhEihztcqGGeXfRKTd8NTQv7pWDcST530hyrJeHU+oyXQroX3EEMqpaRyF9yYx8EXzW
Y9SD7RliRno6AnCiPce00Y7lM69u/7a4pXOHZVbIFk98LwWCpzE8SZ6G6NnanYxP90SrE+q1P8yt
6TP/EcDKjRjCni/i5v36ArU4SYl4xsAb0UaHQv4iWQYlwwxrxv2vZbLcWVTWVACdAw9bHDIV4Slj
oAZDYT8k+mH+0FFszTjZ2xSy9LWdFb1Y3FfkbWmdz228/arPnl27m38+altXRZaDJn8IoyOseAgF
NOqHMLA76uGSI673rwnssrFHqWTYt6CHo1s/G+59tp0QcY2HbzDHcsJJdyi8PuA1vOItQi9mCNgc
EAJ2nyJspunfdEbpwUf4UFp5av0M9PvrgrQ2HHt9+20wJo2DwKr4q2S3EljRDmjBDMNoKiBZz0LN
iscMn3QQHFbDTa7IggVjvsJmS5IWTEDO1b1hr1xbEvceCgkFictmhxPXBZA1xwdthqpPz0pbLrBi
QLlmAI41KdOGAX0aQ/TRNdXNhqleaseXGH/NLpkboFii/evxugwtm/4gl5C7RDiybKDoVBcZwlgJ
FHFm/1C7GzcM0KwUW4oL0zcSVmMCjhbID96AfEqsIAOB041+iaBy8aVdkfQOWvSgv4PgCLS8lW29
F6kCvm6CB8DbVZTI4koIJQrsS28YkgiTcMOA/mJnA3JkJmp99DWMRqekzL+syAwTnXn67wOH6ISo
s5WGIkjHSDeii1bGqXH5Plav8kJBzHGxfYxJkBpw8d4DfvUL/xP982HgL7VtkJ0aXNBzdJe0hjTL
wnOXLF43qZMTAhLzilYS27v9MiAWXBdToX8zwC9uf94GcV7qETKkl3TGPSwbeDdhbZewFbJ4IEX/
F4Xeom63gC4G9YmShYCwboqxRU7EiZmFfGEIFiy29p1TIAWwQ6is+1TdoZCyQWMOCL/fcxUeQdx6
5SGP1hciEeavq48LATUsDrPBG3YkN6jI7tHCbwzXcEnhoc8/tUcdQRYinkCLLPkIl7GBo1oaXT67
gh1iW8VVbap8LD+3b1bPSUGYEfLwWuuxbPwoBHk46TUil2vxu3/8I8MVGn7ouYCHs+ROLUIv2zoU
775+lgBeKOA4eloxKGDuHyBPWySbCKJeUOcvUuyW21rwmTmUpkoWXfEN80Vg6H35o3WkXBdrLGdx
RTuHb7LHO5BwvaYg5au4f+n7QSOxSJHKCqrGQqqxRJWzr4qTVygirpw/fORpSDOWUBL//n8X++wT
+M3m9zagmCpPgueokkkgXUMpR2TsbFKghEWJRVOGG+0bcPDEsPoabNeefPmA+s2utkKBPPR2EzKW
huK4VBDxCFC20PL3evmL+5o5YZzC81PHbLFifCLVLl3oLj+hvV/mRLri2FPKi8JBWuUtLAV0Vf03
Y05GvB+Vm7FSu2JOjZzmHghEb+1UO2YHiDA+vG/2DPsRYbmRISoYZui8R5hp+kV0eAolivuL0es7
n35x/ibEp8fHmrS6whNHwi1LEdzup2yMUygZR2OnX8B17Gr+99UbN0WLW+BZ8a9JVFy+8GmMNLZN
dmt4oXWDuakuW92E8BnT2woK9bOjl/ypxDHJliEv6W1T9CHOr+6JbcnZpghwKoc1gFztNNAG/0MM
682yMls3F13IVyTk0giParg5KBwOPF0A8gFdk13SvzRwtZFXabv5j66tQ3dgbGfO/DMS12SeF0gs
mN6WOeTjg9dAJpPYEtDL69NQzoeSjasw/Bc9VlykC5He5qMhfBh8LVsbOuZVdIcjh9WsP54X3uxe
MA+JJzltZOZLF269MryJgXCksKBB928uQY32PqKo2uXyEVhqWDp/bZb7nJSoi88ccKw9j4YMI5DX
IxmQV/1dohtuG91WKTZet2eX3gtGXS4QW7vuCCPXKdOnV5wARmAY5QljpInVri9X8OQRmd7fw2vE
rEjH58IQUeRPl5fIGFOU/kRiSplg0U5eOLh37FU809aIegSc55hgsKEGmsyqFJSQ6dycQpcwI55K
a6OvTXDsZTFnYjlI/K97STdjzWqrW4dRYoRxKUcPOA+ycq0jGS+BJAMdSLiR2p4p2IKn+Hwd8hM4
j6rGFA/5Q/4OYwvxlF4ryWjUmMz5i1+YGkgmdhIHP0XmNLohZxvKzKGshkleB6UVcZ3iNSxNoOvz
VPZmNEk2p2D08QEo3BcFMfFjpdeIK8N5ChyEtsnDHWVdeDxo+d3EnbIWyw/tCklXbTtPT9Wuht26
ljnlhPo2cO1Fttl+gKho8XhHaDQJ/cR9XaPO7xu1Q4lCB+xpqR4YK9bk60Wyfn0r+WFTL2o2VEwR
QYJVosjy7Av2K0jUlRekwy0vP2chYpcrTQVJigAyKAFBmLQE5KBkTPAd4HNN5n3ohQw3Xy68HIh3
TmVHuotDUMXBvxlATXcR/1cfOO2reelPCj8nN5v+Z5gjo9CkVR6yGHAXBWLH6ai5i+nrnZSGwbbB
md70ei70WUuMwbVGufdiZfbZJv/BzdHLvZnI+8fEVdJGDD6/gwMjSGF4cdtX+6f5wzOJebFeKfxP
gVnYdlpVvUxc5jFszgCExyFExtRDLTqU3ElDm3ymHdDCLXbcvybj/W8mWqZhC40p2r7grBXRXWmk
HcxlyoFjzd/V037L7osA4enb8lX4t/BFqWGEmmat0dZdL8D42VKBHBKebM4/EBAmYLm7NW1CgNqT
M34OIhKE5UtWIuzkA39PiBeevjGpN0XDZpbIkPM+pSOBcFlKuPdSUYA+YNxe8dpdIfljPw8RvIsb
pFOa8yiAVhtv2rALPJOsniTqzyI0w5jlwoVbrwmSA5w8NgfH99GL0fyUpN5qLDHOiaZj/jNS8JlG
+HCpMLRDAIJqs6eXk+70JNeSvk5c6cNyO96j2B34mD4GKA/9FsGrAWXjMq+i3M4jfjvkhFrk84Qg
ntqHWHSmgfgYca9qsqaSYAllauoWj+DmRoYnV6SrYD8hBlAqNfuQi6RWuyKziWKlv8oZ+uazyl8i
Dk0+58iz+Mg+RgogQBXA8nhyvRMfrAqYCrMR3Hi93MELEDQUtku0UtHBZFZ5UcAVRYiEkrGl7nOX
7Slf3pQ856LL5VUstXnd8bI47H/WC7ynTAj7a/APtxzNXIyxD8QHSZKatRFjiBoA+lZY7EMYp/Eh
vc6sBauzLrjraiC7ikEHSXKYpBnfDuwqNqWQMvxkGQBovSPMXicSOi5Kyw2pwEy5LSNMXq0LTi5q
LFZsP0wHGQs0M3JL+6PEI6sFmX+ii8q5iFCZLmkhvrK3mjl9a/oQLFUvE92u9cBfAzd9q+SRLZ0D
Gs2UcXHvf/47kp3pZNrwflOgBV9tjHHMF21WGNMjPmq+5lXlZS1rPjIRzR8xwbnWAg+3FnlG3stQ
pOHQQjMg6aR3FZaRjsw+GJfIRriTsgusXT97VAf6R3UXYgYY35/8KbmLq3Zy8BBT5y1zI4fl5x6j
WUCOob25iVms3dWtenvMNvbBJWmr9SLwpf1BZoasaxLrbsmXQkQxX850MD9bC6F06YbHYkGL1f9Z
dScXOWt0vh9ztyq991bVowuSF/ANDSV3cei2On4L7lOAAPEqc1IJGNzc/XoR0A9v1E6hi39PSIY6
HZqJ9sjhbppN67l6PLO05T6ZFfG/5zKmOXeXvXGNyemFiuDqaROfgq/cHzCD1K7GCz1Jbt0M9xMS
rOtJ13M4756gWO31IxmZHDMleAvO7W2i43lXP0D/rpdDcWRMKC/EBLA3EC20WwEBF8nEtloPhfEO
yUhffD3tm8fcgqnUSMFNWImQE7YHBCx1+qWHBiLW9gl3BqNjgAKQx8eWblWKSZayu+zWHOlfnmo+
rY2OWad3AXsyXuTQGgRHFosbeFY6EF+3vzYSkKjtstddkI5Mm7qw2a/hZXSQ/fEo7RKtqXRAuCCx
2aRzUXvpWIQ/OvbLWmkTNHPZHrcIkfh7Ui1etTV/tPpascKs6VCokqiVSrUJI77gLRQ98tp0SOSL
JmHWUK9krJ/9v5tN2NoERbJDXeP4X1bXRPOSOAJppSjmFj1qeZeUmc7kHe+tL6wd7NYtqqTVf+zd
D8sLVnHTY7SLccWELpQN5L+F9rk+t3rDWR7EG8CdLR63b6WJE7MR6epVjMD01TlhSQEl+RrsZOYL
OR4jW/yXxsnOUxnoxaCsx8ywhAZG3PZmcwYxu+XNnj5/NQMU9m7+ViF0xhDlyhbZt+CU9ttazV5M
M+XJyW3OPzp0639KQOdt97wdXK9s5tnIsp91zzFelr9yH96NNmms7o9qm8GU9ktxEU92nJCAYuRz
Tm8Sf0Y5DmaKj2DbU2ZD6tgrfhjNqkEm5hyz9W95eMGC+7/HfsI/VJDAGXe9RHmVnKFe5U4Qi2Th
YgbiGdzgQJ804F8GurQj1zKAHsWPaajvSZ1pDbZ+RBB+vfsqg5/RGFp2OfVPBJglBvszK5Qs+Nnr
S7JrCYIeduJ+e/EgUKQwBdJNfkP9+2MwZlgzBba7RI2E5Ks51bVtP2X7pfdVN5U6+62Gf/3pd/xT
1PfZwbVRG0MZ8Yrkp1H/4jkQFIb3NVVx6NYQVT69urFaVkOxJCc4uivO9PIIQ7dMSkZsEEhQEabt
DQtpZn6DBFOyubu32rB5lwutKt4nEHkUqvDDLIvPDcNaWfWfGa30+waeYBgZud1GVu7BvWpgNUHg
7lmj0+FG2LUYes2UrSt2T75FyCVGjO9Rmt9lLII9t5I97Kr08N64IY7QHMC8q+s+phFe5tmpvzTb
tK99vYPq1Mn/XfMgFi4q13pJVBPaK+RDjSXT7BA+ZT0efS6oGzqVs2y0D6SbD+FC8iuTfxOqWUAw
nPXcx0iAFguivkV46C7T+oD1eUtICKO3qg8sKU18KHqirrfIlUTdMCatyx8FocXUYWtrRli9jaEj
R0na0E58B3mePKc+nJ4+qI7ka+DtLCNCcmUSmzWF2oJ7t3FFQjqXDan+NXsmyhvNaVmPDaeS2+Ua
dZw+hFfBlFZMxjOtxf/fOq/E+p344twrstoi7wbjdlDHJz8TJGG4Eh4J+TBNL3x9hAMhlAh5Hlel
HAFwe4ojlxrKEDNbNkCWUogQj9cRqoOazNGdzSK8QsT8IdbZBHasYCA/iXXdSzoB0z8YHJr53Hkx
Itg2OAKkgUEhAkkoyRICCQvSLHcUvF5V3QF7zodSF9xZ2Mk79Hz9H+oGIfbmUC87zvW3j0Th4qIL
pnOrl5sJgv4+UDgP8OFrxtsdTNl3mB3q/UbRXrPLzgLX+rdNVlMj5eZkTzjCX69bVwCfyFQ8g2s+
VP4AozWnGKHxBq715ElSmCmqgNQ24OfdeHolKmhQqOlAl7BKteLQqghalO3ViLAI+ZPxlAJ1cO27
jUkka1Ex+6sZ6wvWqE6AppNF+sVG+2tBMulF8WCuVe9yPYVgM/G/U9AdZzatZF3VBi16iu1g+bE+
dMg9QPiquRlF+NRTRfGVs+yvupvTdCCEYtd1ZajFJ1jkSM97ICvjwVRQJOSzzi6wmhIvvA6OcLtW
YEWIdJw8LvP6HAuTuuVzsPhNmB/ncIAMrxK6Mh2gs5OzUJzb1iY4M0K5FihXOikix71g7P6CZTZ5
ok7c1kt80mS3EITmwIZ5vheB22Ydr4z5A+CNNHFS2XfxddZMu6wWlknGt5c3crcx7H8q3UY9UAHR
qXaraOX835udBfIxfCQfUWOglsDPSBhi+Uq9iRZhMAVmc4Jrf5NuQFKqtPgiEFStGwgDLcJCIWVr
LdO5Y+ow6P899BIS2kONFTQLSx60G6TcuNqWgEYyiJzxz85iq6vF9fcFQ9j0mdwEeGkbyfEXzEKI
GOrD82EnFf05W8CsR3hJxDuSRTRODyyEo1MX7+ZiYBbASYaV/xA5rSrge+/yCEorMVCruNpv0BbN
ntPLJ7lhVOkm9ORvryH1k1V/V6FYVEBkc+weeOOW9JloUzgstqtuK8QpwId18MPcIBwqxAfKfLF+
LN30fMzABJXnIoLqMX6DE+r/Z6a+5TS/87JPgpyzOpbXzc/0sraH4JP/Vtw9Hh6vBftAD7DrjnHq
bIi+qzvYFM/W2LCnufLvL5v3YU2GeeG4uvY7mV9TpSR2JCTTdqo4nuJL+z2BNoqE3xjl7mFZX1qe
hpGvEgmqkTTaMTzdNc551NmqhrOF43gkF1QhDoEsyh2PRcA9GETeoyP7g9DU9Ub4dMSq9dklpkRH
Nluo0gzTqOQOtzOxHu41zaplZi+O5p+75UeoQJCZMrAn8pvJzqIJb7r2qNNgTixAIHSqCQF4d17U
uZgW3LgEbUi+W+waEE+PgQ7XGRCvXLrBOwAGhvX+sjaUAdJzQq8YXZCy6jKxYEXdY5VwB8BipM95
bt82XhtlEdYn3+PGx00lFV9LHu04NfKshnEWIqxrAKmASV6dfREIPlw+NMwZTohS7A3pDSjR65oD
t5VPNYnKTZ9EzCQ1jd1QsuhWqsGxG/5/mqHwa3Rk+M15fKUQKEw8hfqiAwyVqGi88eIlUVdO5Kqx
lshek/9xLKTczf9yOAY9BozqlkipRJuuq049KNqSLlMkylTwg21BTa08UncEqEMUd0tSBJ0bPavV
VlEB5V7oFgIBM96v4qEQl3NhH8nvSh6Zl9U9b1heI3fNszfLdAqQ/N+RH5gOXrVgEoD6SDhsZaNw
Lj1z+OhHgbqw74z891k1O3PbjSO/2Dd05oZBC2wLYyAgfyOlsK7mPvyusMp7txjJN4IFm136R2kn
IhEZfMnYV0KeEX99Xp9TkvZ/vcPewi0h5JZ07kMZ8zp3C1iYPmF8Hr2sqzTtxDx2ANoMbGYVeswG
4ZChDVSVd7FcU9sVXcUFowsQ61sNZxeCzHTHY7M1jD+ieFVxOFBJP1Facw8shFVR1tGRKz5T5ouq
dXnRmOdLGUdDFaZWdmeQKCy6cbpgeLGrOpmASUxKZAeE1npgCkwiFsDvKg0F8+893eonC5mzZWYI
UuWyl/ItR3QwYqYPBdEoNgiA6yOnm/lUNT/HgyHugdmm9Qg+sVDuABu3/uV1ts6OEPCWUaYwWXw5
3iCoCHcQwlTyRtls3ZendK+pM+G5U4PXLnyFSFpjINB+OnBw5Sc8zZilFncWSqZAsFz4srDH4mmo
x3mhW/sZpH6NCl+HYcVAVCqwSnbSbb6HnCJD4uaptNTyyONyqcb3nRZ9ULCLFnQVEvjun6xNv9Qw
Z8Dpj20n/RMp0pkNUxG4RZIWePGWYdfaeXBxrVgHJMx+tjIjiY8Jw84DB/3qRW8GZ5hq0tXWXdQy
eiKOO5IWyFUYNvUvK9vOQdmUW8wKQWURs0ABLBRehJE6ZStEXRD4YePOEjXN0IzkkTamnu+XTETc
PVkHZ4KMxwiewDSMTHxCdWuHvRsFje5ZIYFNr7RT6qVoZhcoKA2egBK6CfG2lFY98iyv4OZclAhA
hnq0qc8WNTVhjpbznXA+358JBY/2wtyCWRdLoYntNJJS9xf15ePkiDVFbBNpV7ax3VVa8XVqwn0j
a73cVfTLUBWcA1jy1ESwbkmierMOSd7frsEeQ5qrAILVWjsek5oEImaa0IqRG6Xkm1RS++UQEbgE
GTc3u9leq4/yy8KWuR3JjZI2wMLRhA1ckQE08wligNzyLVndIrPhFjiKpsWf5LFUjYdTAqM0mXOn
C8eIlcgSWVFdsSdyaFf0EkYmcvnh+IPsX3DElzLQGmWLpcj6GpAdIAtxYdnXrPMNTMZfVCIMKnIR
U/Y0szS57lezv5+p7KS5d9xJIzSv6qyedn23vyRHVcOYlAL/VO2jvFFqKl2i7ZmR1jfE/itb9SAk
b1tWBdDkaPQgR97YSWA/7Ioi+aQPeSU7U4CRfVjMHUHlhn6SBPGZJIf070P5ZNgdylReXvstPht7
T7O2Yw7t8TMiid/cxusez0ccwX5+UIhRZpFR1Lm29bzfRYjWnSKc2tIm3xRmaZNmq8lBSFHxRymq
qEpEGHHjp/rH6n/z3sFaMlOZ0bMsxesUpKLhnEVKyBqS03SexZlQ9Qos+BS2Oqr12p+MbC76W0Xb
A6XuV9Y/bZNX3a+XUZlqMMCTHovD1AnN1ufgndPx4crX3WEmRUatW1wiBMa6WYrIJI7bDW1/PxQR
n1OAYNY0YXzfgznvYF2WJlW8esT/MdTg+UXiMWBkTbP3bCFaQLmshj1phWxf2f8uopJFFbcVUDYu
UXrqDkBVfBEsA1XRd20cEIGDJBhDCb6bPr39pOUPD/WfQuAa19Cxukkyf4vrUQfVXWlZ91HexkOG
wAzkVPqEltCCaNxGZRO5Xi7DGjMIeSFsZjhGxx/ebS+HNx748NbJOFV+02RUUivhqKLPUo1uuCwQ
8J/7HJhC9CRzg3SLeP7VbEo0FN2yvXm3JhuRhw60TEHFiOf8S/D+t+B96lekGW04JHGIVGopTgkX
HiOAPkhiPn8yy2A20Sz8zGolFPseVYQ7oqXbF/oroRnUgc6S4SfcFycOlqZfiTCI//07TGVpTgC9
ea0CeljBD03yhIWW5aajvblGE26NlMyk/9qAJjbH3JbVVX9dFj0m0jz4qbWEInRSVKtDE7AsdUD4
lAUpcOmPs2tPmtPQBTaTzeJkQZHS0bIx/xFrBYu4+wYHd7PjNDjLO2Ybxvgd+hgIYy1INQdRRrw1
KbewGl0uRfNi4k/wDiSOn2Cu04ymYe//K6+ZEPw/02CiAYZYMDVii+cb7IHifxJYymFvZ9BLB0zf
tRw1gjK8Igj6mFKI53qa8qTWK+fyeXZ45KLiOO9/D6E42Y9HBDxvSiZU/0cWlX2sKDlWlMeTlNOz
IrswqW6zzwmfAMDPY842cvKzg6w31GyQxts0DVCpr4wabhNwDsj1bilvhL0nqOwZ99xijfJzG5RU
jdeCQL8NdsQPMs6LMdykAM1ZDt4HBeQTutTNYw42fa9Dz3diPZoZN5ORC918LCQyCx8fxl9dTJU9
xa7wptKmmY9cRYThhUT60TfVFEnPmyurZshvxjRlnVvSm2BSgjeIEjhlwRrUbYrTgjofddO6Z91q
1oix+342s3X5EtT14MZLe564MM8QHrVfWovfWVJxOYtojAADFegMm6O+D+9aSJW1GjPxYLJnVWR0
rv85Tbup48mNbrq9YtlIujtCqn1k9kI+4Ct0SubYs7t5wdsmQqUCtkpl3dZWBOHJQQgdyUoybJfZ
KAtce71pPjDkg4gv/9ksdaz3ZkoTNHy7uQIC0ur2vo/nwY4eAZ5CHwmIkLuQ6O/Fld4Avw/Z7uYz
gWOXtC/ko00/NXcJ/HMzrwbLHjke3CqC0zctm+SD8IIpzGLoaaNMk23DDiG6YHtQ25ui1CjSUrpp
tz50dibERePSukOV9MEhj74pfoPJdg50sJXZTWjdfIJOAT8UkmbKvYALJfeGlY0LMhHPRgcfpFL0
V7arcXF1pKggbv0YcVNY2DpxmQHIp68gCK553FySdJqWeXNEvT6olG7JKvdW1dZPYBFZV4+Fj55J
o6igDAmuCALhR0Yd1aqxO3PsjrNFomTiTVGdCTezQ5tt1tgSwG80tItaooYgRYBrFrj0ptoeiGu/
zYc5nvFVtrBXe4Rr1bW5pJV3hp6zflBEpJJYWL/cBYQBaWwN7aGPhcaEUKqU271gb3XmDZcmWVj9
QOjjculNj5qphccGVt1j0KzdVpOiRNX0s68pgJXaQeow9WpWmOf+kA/0lIc0QCp/FLKIV+zC88w5
DBSCz2ag+RHzoKwSnMs5LlOPtI2001R+QC9sQqhM4knYyL43mvSyA+UWzuSPjJWiKOqbSV8ISHXm
h5EOvPZiLRATeBOahenbSZpe/prQCK7qp6vNQpZYVib6AlJhbMGo+43+vJs+cDx4tPuBIeqEGUM8
mfTGMiYxA4pO9JCv/KkBGK1wmTXef2Ddkfe7agvILozv1+qkCymcZb/HXIoED+GYdxRq8jWzmX3t
hQBHcHEEmANdDLORMJbpxq89PUetgkxdPH3a9qK08L4pek8Vyobb5iZVmIdkpag7bJ64vOvIM673
W/3dRRDmYkOAnGpdcjU90kUlgvbt9pXcruA7f0ar94S5PJNnZfaf15aFT0q3KVgNFcT64eCp0OXt
xiYJzyu4wwEectYuGRaTceSKGYXaqFupJDL0o4OgZbnAodtAHzgYOhtm/7TvgiYyN1lTyA23UntI
p1F/95eW7Aa25LjuBrDR2cWKkWfa9I9iO5xHvfsmwHTT9GTY9LOKmYGQu6KjCDBwZeu60oUou2se
avHAm2CE8BQdPXGMQtVj0x6lnokH4CKqfM5w9rly9BZ0mXJbB9Z5s1SW6Y3MzqVQ1JlRMklbuCQz
KFk5b6Eudy03s5MkU4BSBo7/KElssH8osAjfKd+e2YXQjO2wYsy/AbDTRnQkd6sGO1Kk6ZsX/QH+
GHY6ivEMHgOnQPxKxJQfHeuv98jR9oUq0n2I2wQkoE3GkYxGB29cbgptETpPTl9XwinwRmxTdXGF
s1Vl02UsT+PE83dIDzCVfLtaZxXcKBY8DdDw0ZSjO8a2t1nF2e5Gaa1kyOGts1wvecBJf+eOf4NO
5BNudKxtlNPen7AUUSxXVczYIIOk0cF0yafQ26lrTuEuMm65U4UuHdJLyrrt7J6OKNkh4hqhM7Vg
q336oyywggywlVrgRwgHZLs8L1OtfRf2U40Td8/6GKhe3uaV1vW8s/4cjb0VPCOoabpgN+lemDoB
JSycE/aDve7mTEuUayJHQrvoRjtr9SA/i+vwQM3VFOId+ZT4fIgxnvd1JDG60oIOEZSqvgf5wvga
bu2EqsNRnD/f2I7vGIZEY/RuCO9sXZVo2DpB9+z/hygYbs5qhgU+54VY5nBI4vWQbqxxOPFv7v26
sFSdi258BzGERvoJYTHITA3pLtPCSOn3yFhRFCNCP5nq3kDvIRO+FzlqAcq+s2TdUqUuUBqdjl46
S25oerkSotOP5S2T1NnTmUfzOv2eLGu2F30/yz+82kXZw7+PRbFRu28dZjlTRgSHlzvpdhFSuUEM
ncI8qE3z1KARQQUNRGMPopyH5JOPZMSsz381zJx856xzzec52oDo6pBS5JA+vmBGWhpvXdYBk81B
dT5Hm4VVkqIu+ZAMB53XNRuvKY5ukVsGZPUtKnNfb+qtcJLb1sslf89O92NwNPd4Pe9/qkm/5n9y
tprI6dZ3f7K8yrPB/+bbLE3N61jhCKJN/Hj95y5EE2+kR6/qp9zPri6mNJ0/MDF2Ue2EeTwnPMo6
Tmu9CcW9oYxLs6Hj+MzqIgOKVwmQkEOKE+EstswkUyMANJACFhNXzxvP84/ZL1qCq8MS8CSvlb69
2Gpbl7DHj9QXbXsfsULPwbLBa5l3GhxFn3JyzWqM63giIKR/2nv7QSE15qjwv/XdrqBDu5XlSEJ7
xfPj6fOgbQG8+p+IiAQY6MC0x0nixwfzghzR3uiOO5UAaCacVuHQRXt6urVo9lrS8peIztCpn3qq
qHmDyLlTT299XRlCa6vzrIWJN3Ipt3LAZjqEI6GMJ98qmQ0HLavtIx2cD2MDAAsmISHDvOKBAi2h
Mf/1jsgZ2IYZEPUPlAvpQ9ZwDSYwLW22KVvgN3qMheq+MeczpGiFMBtAcTqAorgekdx+YV+2ZBIS
1BHaZqHGFQhrf7VToLDukXmvyGCLNWv/OB4hWfd8fJlfM0a/kPTk0C5V0GskqFrYVuC50MQo9w4b
VqL1Eui1ZkswJGxYXGT8UDa714VClxO04on37/D4dMTxdrJqJtYfk3sBjfdsX0w3+dpEw3zc2Uk9
+BQcCOknsZrvX64g1CxMxG0fru5t4NgGrRYxnRUyZdkpFPUTphAEni6uppoSMB/2/UC1yG5PCCBx
wsgUboRLYTa6OJV2/NxQOiwGQ6AWR21SkBd+6yUapHDJQ9qjwM+Le57HXMQsYruRiKuR3sAOX88D
mGCJ/6ht9pwmT5Z1g373P3rnEQ9wJRwYaHjEmj6s1ingXOSxHgHM4QUkyy15dhE2vu2GJgEpU0Tr
hLRvvCJHqgZzpE6Ij7YRGvvhyp9M8xYQjZmBDgQ5kv2Ki7Emp3tZu3dfRXcTHKo1qncdaeKC5Gr/
UEmdvwe2AeJqXNgXzYngjZ9r/s8dv8yvE+CjcErd21BUkRF74bZEAl/opwf5gRAifzgQ5TIVNaZ4
XM7c8YDQA5puJW1wl8fEYtANRU5CoyoWN/QL1myX/sa/6cHUFjmRUZK8CxKC/D3Y0hBvT19f+L2P
9UB++fmZ8+LC3MZJbM/lU9QMCT+rnquX/vCn16L6dKjem56yCBCpu/dsGWuYscB3lalzoKE5whan
Qt1dPNthUow8eM+caDtrscyqSDqkAp6Iz59ZTSvWdmX7BWVvqUNNoFhOJ3lIE1QoXCHFQu7mvQ0K
4W+Cl+wwLtcYah4YCqQ/h80tNDJeoJl87fPb5ByhcfF18SePSR5Kvyv9ZOnPhEWlL151lZfl3Sqz
1EWTZaAbbUo0M5R5/PMx7ch3WPRnI6huqZ03QEJlGx+dNohJ1yfzloYV31ebsdhQLAG2FcycBx0m
+XQC8Hw58B4fG2nyEo3wzXGJocrH/vNAn79PGXWEKRFK/Tf2OfzEZQXXwZZSshFVKGa1twp6tR2I
sAmSQUaYUCiJ2ZwNlCNYmvHeqBHr38NraDZnFWdli1UJyvuZAfAxyCC4OKiPBOoUQJ1N7/F8mrs0
NGIwHOiWhCJMC+BehVId7OQ7+uBCf+X+ISA5nObSb8TxCe5tLzcvo8QjxKS/FBxQzzqv/fhj95bb
XYvaiOJ+d8nJw7NGa4ceg1J5b0V5XVPzvPr8WeSLw0JzSrYPe8b+TkXUxWFNCr/hsj8qt/PBeIbi
kn78hYOZ7hp8Tcfqn8AAmKJpBd/Gt0CLaUjvgkQPBlGA+BH5vsVweUSb7alsqi8yqcm8FP8zzU7Q
79txulrfEPSPuTsIZXxhmnSlBSXDk5iMd1FP66ETHZVfNomgj4RArmAT4xCHqOC8kauCCYep9yda
DS+b4G/ShCdl+ce6wC29HL18yzUeYgwNpWHlTMGoPNCAqIULZ0TrW8BfZGHg5o07ijhlbdLW7LJ1
4O/t37DBNZ/yLT/Noax/ctM/LuX/F9N3wnIhP53xdTeE5yD6TZSFPeMaxpyr+1PpqmtPGAnzgkCb
TGeHXxWJ/C43Jwnq4x3HwRh33tSV0pnracAQx+MZtX32fji788z3TUgebPcV718jLAdue+1ovJxX
cS4OO5QnSjq496WLiEq5GqUC4GrXEyGRQQ4g25mWU4gnPPmKROkeIHKR4IXd0iFrNaw3CV7VzjUA
ZHaK1eVdHtMr8kIGO/7PMkGtya9ZeZI2D5V+AqS5Gm2qDpXmd0is3BxpEf1oN/4En0wQeH2I2opl
yCdmUFgHh8dapK03V0M+a6IjJu5uBPz7bIJMGiApEf4pWh82Wmo8YPt0DPu7nHPxeYChf755KV8g
2y3ir6QaOJhxtQQpWrwET0hCLbwyPGFS4tScZujNdGBGkhM5ELX+2Z6GUtdAIy3gXIbd8TrjXFb0
riox5sdaqWJIa7yFOZrcwcfHucgGDR11+PLMXALlqUPRJem+2q2KzGFjihJFxHgoJ1xUPzhTO0mF
h3FZ6GXRB2fIMTNNEx06NoH58LcNN5FAnSj+wQ/EzKoQNu9e+7eOq5wnZ6SzJhbFDYr/ywCqBJlz
aMUA4yRt1EPAx0nfnhkdjYyY4Ybfj+8FGGqj/MyuvI1Owzi9Gv2eBYJMuy9bU+iF5bY5rWjxO8sA
FGmEWi9TKmqc+TSeidiGMjMDAjD1H89aCWFaFAx1/7od+GlRNlXtXCl/RdD5xvY7keYOtnLuiiEt
nOq5XTUwVj0F/VWr9utw+ia6U1lIAfY1SH2382O3cr0FqfN4JIMqwXmyypOhkvaVbAS/CvnmW6W5
KsBKtjqMmCN+AYXi8WUiLl0rLdkU3zXadfYe3a0H1PW8uaL5vG9GvJNb5AcOZIeBMFvtexpyXHjU
QxfXapeSJyg3tsij+5f4nHSMxM1YlNdUxBbGhtYLF/043fyAIxkofoV7OA2C3wXWTbyq5rgknj0p
aqjZIVIJVd2jXFqEE9Osj6kRAHXcQlUq6AFIYoXtRteO8esj1mp9SV6U6gisnVJtV56Oq16Oz/WQ
lhxJF4n4vviVF753tfAHBsCMlISGLJDnaG/4NMwEzEoQnZPbWoZFSq1f7VuPChyEjwDK6tbH20L7
/CMhI0SvvvA+6FIGj0OjHYjaj3P+lwd7cSHUG+5vWCSCbtX/v7BnYO8esqgMaAPcmsxNIi2Bnsky
VUMTt8CQTPKmFEufgN66eYwbJ5OHKA4UuOgtdRxUMnKbT7UpplOlPOlk/GQiMILfs6BQBlam9htn
YIxTmoBv8RNBDbn6ekjF1wUkR62yvlATcXWR4dP4UmOWvagEZsFoQbuz1FMq5B6/iRwuzrxss/ZZ
o2AcJNQzMVTmEfeEY2BazNJ/lfhVe9WlqT4jh5CS2l/CfnsANoaTs85SeOy0uOBAzORopRe77yWm
CwpJ9Zl7UyTPJ3kPjAF+/roByo+PPts7hqbXG9qWHZvTBQCBxAQ9S2vdA7JgqyUaB2tusVftV/yL
J2bKKj1Dw74To90ynDjoAqYl+TlRU5vCTLswoRLnXuvNsOE0Y3HRBvVYjXNPipfw6py+uqvtyjVT
/ncw6qIvdkjqi9f4HNaq0Rz+7P010WzKWOHPkuqkmOq1jLi4zdyF/L8Mas1vNZSFlqMS5R1A+plo
K45Awi4hfUEc1Sh6vj2a3hMfEawdNkiapMTBB6AZ8n50UhBo+eYNGNaWPYZLdlK4OtMjAClBybsR
25mzG5ai8E4niJ5x0UbQFdXg+ByDe20sjcO9cqzIjoZrOztj7RgoVfyjQ8wZhaF3t1cpQqiOTVGE
hgHtpZ3PzHUmejJBjadvnKovbC0VhC6QQYTmed8WK26/QslJ+HymLSmLbs7UGzuv+quSHwvFBZdI
KR5/QGAGNaIR7z9HqdJ/PKxwjnp0e5t1EQIzZsB/4FuH3Hz1C2EkuymURTwYDeISbgbjmrG+oGRI
UPXRVL4OP1DsTHCFBhGO91HPzPuY0i0Eh0X6EMjmAXVsLyoX7RJKBFEhhIE3hjlhffVIqR+lEaYD
JA4gzbHtAvriz92zEsMGMpx+tbtbYaYrm9cEJvbL6HbepgrFfhwu6Uri5EN94yxB6gWk93LHgil1
bk28UTa0czgmML2IuH+xbK5c1R92EbE4EHdd4w8DflQQa/mZDHQtlL40iik5sp/NHFrTrCw1xomh
WlcqWQqw4TdXp8aUMSbHk0IeMIaMqBEzjtIH/phAdl0jtYE3xDEmuEqzJprL0noQImZCLrwErxwU
l6hYwvytgjSKrw2BIisSUrP3vcbolV5Laic15bNbFB3DUQp+xTb7F2JD5J3R7PHx4h9LrE8263hf
FLXNyZCRmRV6v554OyNOaqGj4QAv6r6bFXVtstknnPty3DizclNF4j7LR31qRkpjJKFagfDT56MF
ooNa/EITofARUikcZ2eGOTXoHsjBbtq2FMWv/MhkoaSNzqxewzEC1yhIqoSODePOzUEolinklHG2
U4J0uPu/CDoUXAj0E4Gel/M6KVQSQE4FP1XByMnGRiydv1bl64V3vzQxJGgBqWikVLi6LBndZIAf
BG+LF10d4uuqI1gaLH539X2kUu+ZbvJ6PnxjBfqNjgLFdqt1YJcLzynRFct0gFt6QL+jc5Xon3yq
XKTduHI4jsZHCESG3+KsRfhmjNMlnyQiVoncr90dOkfFqlK60xGFwvRaRiV4uTbjFJBo46PQXJ0U
l+cweCPom6IgRdbrynw90zxvh5rgQO3F131nCIQrSoCZ4nNYtYU8Y7IuBAzsCew++ip+HGip1JLQ
7gUu4ADkaGIqxS0MlLsPoCUB9XFIVuKVXTfYkzf+WYI9pnA/XB4RJH3Lj2JUeNN9SHtbKU1GFPP4
gItAML2DepJc8F7+CxKIOLcd/W/ERXBqb8Utg3XduFzov4BhKadmm7obHftontOY9+PuZnXF0FC+
gDyVUPn1KDRAIdGc5mXQ82ucm3Gyby2MuJ4CBG8LBDA6Yv+Su+gvdzYNEqjcdUbwrzlFPmFkF1M/
tVHzj9S+iqGU3NgYBlcCnHzdcw1ZU3X0WYAgU6rPaTJrG2w/ziHpDzOZLro7pkXFjUC9pbGVvJK2
uimpvn3KiT+mdkHYtZuX7gSCmZ1RSMQDtAsqE1t7CTesMZu9alcOAZxauEZ41zZLQ2TAhBhT8pgF
PZLk9cNHUpSh5uNXo4kQojC4muANghHYuZpL6Y/J2GAwutnDKxLU/rfsucSVo3Hwu+j63xn0znJF
FbrGJNKAqbceiGVDlSb2hompQco9sawOzlrciGn6eJeP439IYu4QvB9C8d4QqDJbdJU8L962+rJD
Epo/j44bLliB4WN9qNyOPYnun8Gec+cgDemrOhjQVtK73BEGoan+vvqB8hqrRnLg6SJ/FH0Qdf9/
AvNtmdCoY90HSjFMpS0lJfsyj54dNssPAuFV5rHId6qlXtO/JmLOShqd5VaoKTAr8U19cN3TZBMq
HSnSSIStxSosPgr0XgEj4NXghuwisHNIaFmSozbwxsaZ7e8luPsozJFMCabb9ZUBFU0c0yZDoYHb
7XFsaUiaRaFgm1zofdXH2ZeLFs9A6/e2343WcSBrGAREloP8mdXqGEqMv4JKuc11IuS80iEpvRrk
XviXHNdtCw4g3kZtMnyS8q+0ZfefYGOQ2HvSaf8VyI7t8hAk9lFT2qTEegKuiwl3mHKDTNzk37pM
ID/0z3MbfG/cWvvc8vf14kadWy7yXU7ltFVyebs/y9wTOSsX56pdV08VTMRAJL2NTC6nSk5vVJXp
oN8lbzDd/ruARx3s5xc/+0KefVV4lB4A8ddfVVmGx6aeXeJSfKc0uooMCBO5ijmjp8vaCE2hWgiY
XyhqUcVqWb6w5jKNi35FMX+IvKFel/Niz8lh3QPiyKoJ4W65HhL1RNSWtoBfV9RhyB7ANZOw8bzo
LiNFmY6dY4/Ul0k16f13V72UbmqryEz76a32olXw3nCA65i8YkxJMnF4fmcD9qt14Z698hU5OsjF
aroh4yyrhrYkLbtWmlxhefYyV0URXSpMiNM4Df+W8mHTLzgX7aeTGFSagscazOXfaJrFFMx3XWV5
9aI+txrzQI3+2aiISp5cAP1OKt9KezK6nIylxMJz8kr9jEYV4ceVqT0a1POkCjHlPfkU8Lv/jcdx
SGeImZsh1IqOIFdeaX8r+osWLmldMerbj/N72IZ2/LEMe3Nu1NW54UY9UE3UcKUudX3OXjqbtQWW
d2+IteEgeK5FHRA92jxfGcZ7n8vK6EBFCkInLOeiu53/7dcLWuqFZGdttkuw5lj5R6Hd/yjaz8CB
7TjFYp746qtTu9wnrXDNvrlz2yHtW/xFW01bJF606mbP28tVeyQB5SsFq9xhMy4onKuQo97VtY/U
9WvNc/zJM/vu/H4no3eNJsjdRJfhCasO10412TAtlHt+UBlcWJ0QBBbK77w+w+wqCnx3YaahiaIv
4qEv7eJiUspHgY8U1zsc/ykAJf5N62dRFvpYYZE5nmvY0QLG7UYb9N1aWH0Lv7dWTVGrK77lat9f
V9TGa3iZEuR6vYJbB1XC4/QBPN9mChd6nhMEYsJqK+NrkkGg/TlLkru2Tsou0Oefd3pNth19Bz16
7X99Qkb7X0oHLd5h/QkmXKfm7/V0yawFwqgqL7J8UN4Cd65fSF3gfXlvxb/o+Y0MT5NJtjqQPKDO
RY6bHLZl1/WX9Fb/HYInN5qkA9aY4BVRz22A+JkYl1b27XZqVlFiX33uzSLZR/R5f8H9J/Hossi+
pcjcHykZl5Vg+AVi4xGyE09a45nrw5SeeQN5TKerZURN/W7iW4X8pTeNNphy76HK/LIMKyiljspv
fB2uOniIZwa10++rwqzfg5dPqaptR8FX+xziOkuRrkUgRwvSug/LgS6VacSr86g8p/LiwQYuVAZL
Gfj5jmfxPmcVekEAsRurROTsXIUgDrd1q31Y9jQdKJE5rSjBnpova4gkRBpyb9CeEyku2FEPSBSf
3sdC4ZAlpEZNyCLQELGIJGueBvbKy+ubi+YKkesfP0pPChcc8VbIN22nNVlkKBqbSy4hu816aQRu
t3p38A6M9dp+XaSmShE1KI99HWK4c+iF/O2vR1PbEG6jFrJbRM/a9RIYG9tIhyIHuzwWl4RDcIU5
7j7EzsWeLlbmPzH6/d7sHl8f3pLLYwM2pZiu7WWQXfMzjB7CqdABbpciCJ0MUjQWbf1jO5voDO4S
zUPrfATnemOaptbC5BtsdT/4/MZeNlQ02lkJgc/WOS+iykqAyX51EGq87RjipLbpaAnLuWd+59xJ
AcF6G39wQ56sMat0sLIs9xyyOEI/25GeP/ux0/I7xrbUNV36CD/RhTMT6Dk0BCRg4pdv/3kQHcQc
jnUJRbtJMdZpJti6G0y2mp6M9kNXFcW203kEPvqcRyY7UuOrSi4FKHjmYVE1oE4KBCRXJGrZ+EKI
Q4ChsXu5SU/JQNnwcx8+1P5zS0vd1NCtpDJQl8z8T8Wxw3xPz/79yPQImxJQwzKpCnrWrrWI9xxG
Q6EmrVze3v4yEKkIUGjLnKl4iBQbIV31yAqONA46hBUFkrIVonFUBEL/NtvFyMf1njMoVF2MkX5C
js7PUflrPQPSps8jNSQ7alNVtYe/foVQ6OpqGkLp/KkAUrYn7ZPtOxkkvJ7bjAoyTVLXaFNd+yXT
ccDCwPbiG1e6emdR/vttdkhCp5R/alHm6s+lW3Jbsh44oD/HO1MASsutzscYS9lYpif2RVF1P2zc
IpqFRcAYZQJ8UTa9YXI2BkUpx0VPOHI+IgF0wAV83ar+dmOBm6un/5Va1LHg/SbGDxTHeozbi+bc
qRAbioPEpAgccnrVN0wAv2tMlm17m4/FY899zzj0WBmNq2qsURKooSAv+/zQS4b5rU5fMx3UYjD8
Dff9GFDkGBOzyy27T2xHgm0DrBMaFm4yL+odO8T4+D/HcbpecKIWbOe3u5VJjM7bWzFC2r7lxpi5
FDBM2YyQWZ+YOcucBWwr8MWBNnaUPH6cOtw8prIci3VARrWEdezu5TuEfsAJ4h36w9GziTz/R2Xx
Rcy3XJ4LH9pMLH+Iv7xTPt7t1I8jfOMGXBmqPp92eRm4Uy/oFUwQCs+g3KTrYhttVtLv3XwMRiJe
ENfAYDitIbiPAE1HlqqdpzpCNFZg2W0gHK3OswEpdh9etgFofX5deLS0mU025FrLOPC64FIjG9Du
6SzF9wgz6s4WDNQULTavQqOU7LXi3u07K94rKHTNIfXX/6BLgB/0TvF1Yo8yCzggHqm+KnQlCK1l
S7n4ljqcrnmtTAcc/B7qfgWKrQ2OlqV+7MERNA+Ua7E/3WeRpH8Cfyl957Lja11m3C3bgzshXXI9
3xF37CflA6AXAXvDHTqUeSI4q4pepWTzcf+8DGFBXda5CA7xwak7almop+Bv0eLTsgfmVuz26ncX
eJDQD2FzmeUFw0qvtw7zwiBKjn9a0cpR7wk1t4eyvuKywMnyGydnltQqldFx1tTZANIzv0+kCk9A
KlNho75paQBAaxHRcPPb1k0fUmuSebWaC7umv39V58hbr3cNw4fj1REpyS8uR+BnQFwYrhQ1bcq9
fNes0QuqPTnxmqQZC2kNzCVRSaRGMZP2Ca7hqmvaVNLqrfsD2zFfFTxFVFog3t1vIIUWIIznfI2N
iMSBh8tTV2jxxWNdMIL0/E4g1NBt5qPwrRuasJ9R/P3PoBwWON/8dcYEmgOR/bYsH1+ajkBjU6tM
OtK7c3tZ4wMfAo1An/4o4iLrw5R0UAHBU1zOUF4VWnUn7lsKTWxFxeA3COYxQs69CS5laPH7S+EX
8wAgvtMxfhzi3OZG/dAkKok8VuNxt5hwl9M5lwYwBNeH+jEd9p//BzevI5XglU/y7aGpp2mTTQrK
ERCaPUlWv0KRDNkHQtQf9ILslESv5nJcgZvXaPiVl+r63ytll5NLn0XKxmX2CHN5C9cqnCySIf1k
aKguZmKvRHOYUFBIdZCw7f+qtm21K/cj9CQYhUC6ipD9qqQXqSOlzuhpsYOTZ9jAvkqG4/fGHEZK
Lm7o7BFeK5fMA1kRQgTah5owFZormouBFaZ+bA3XwqwGP1OiYTja5N5wfNNkfbwSrGrCZX5GWG+s
jsKzrjOTvuGdcBiN7Fu520+jvtEuZrTtIhsM3cVKYAJwLpHv+Bf0SHLWqWPG7q8nLYwbRHQkEAeD
+MTznOpPdsJ7nqEFmSHO2JzdL/EQQ14+J0WBmeSx4EuV/4ylroCRpklhsJF0R7aRK49nx1IOlTLt
geqEdRQkj69eCem5HCaGPNd010JEY/l1a1VcW3hwsODix6gm42gu+bR6I/l36o4aTqEbVVtl/GKa
Zv/wA+wrzjjQmHWqepBPjckivqYiaYMSwbf3Goz8dBZBTzFt1Ez+HeNBcD3JRysbsTQXMPz4cAIr
ZHVLfTXM4rCsZEfuJri5ml7cXFhsRel2UC4GZfX5zalrTYZ6k89unHr2+/MWUHMSaee6q8DkLdS7
C19kQfhoQBHqtNSfbtQcktp0ngRCS3rh6y6uLt7jDbeonYWoK9QyZ+5JKv6urA14bOShkFfdX1Hh
DlZb9W8BMavqkT4nbPDOjEiO4L97Cr5bMfRagOMao0ewVItsu1F5dv29oOPs9YKCHh/4reXuto48
uF/lxr3uMmsfbYxIPocKKSQ68fsQ+4BIVOnukU5MiEG7MJuUJ/WVy+GJTk5CTf3BcTlj+L00R1id
vi/1jfBlXzKJn7c/LsZ+eGi28xHg6a+y+/IzyypLS+UQRdzfL0mVuRN2tTnVz7x1pkfuHJuM1Vou
S1u1RciWQUY1WazLkxM5ymyZ+QvIo0f8nZL5zrPxnMvwOLP7da6LOJwCcHQJBoQu0nVMo4jX0s+R
yqRbfv7G/jGoGAIH04D15r9oF41yENwfk96sU9TocM2AtNXVLSPvsJrSgp2+hZRePlERQko3R2Nt
zyMQQbhwsrzqH+0a6+lcLVCGOFMP3En3RpdVGMhyXD7/pu3OLYSo3RDOL8USttS7rnSESDV+mUvB
w4UhM7xphPIQPcsli+EbWYlJ5VTWb9GlY7QSI+PJYrzbsiB07iXg4eMR9bWGGktkgHAI+3mFtUAK
m7PUdG0zN8H9J3lJxQTs+xPKUrtEbSOcCTLqC3iAqamzwqIehXv1eg9Q3oK0Q7xX7qztSossJveX
yhpbFu3wGeLzwDP0Cno/60Mgq6pqdWrLXq6ky69py4FlATlw6giGgKvrgZvVdCm8Dn5R0oDmuLzl
4pclqJYNXFXPtXgFnC+0G+NAUAhnZxFZPq5v7rWLTURT/VMkKi+XFHb8xpHtIb/p7Sa6Tqf/xt1X
uvd46LnLcX4aeNhwg27oWaQHryD9lZc2IrH1A87PWDUi2Z4p4DqtZanMTESXomfW6+wQPkrhtSP4
bQQRC3aMfy7JOeZ/1a+Y6WGFhyq9bkcKMZkt+3vBKD1ViDxcbx5aqYnwbCpTrQgT+sxrSbYczdCt
16JQtcOtpg9zXsiuZ2rotFFXZA2tFfslmU0IUdMOMjcvA98qjZHo+xokUcbl4eyTaU2icqTaf9kT
BgG4EapBwE+FV83Oi32uEBF0fvYpwohqcKtiOMiq3QwTJ0uytVNcQWJe+bQnX8/ER+PIlRXXkqfW
OFYWXkhAejnz8qBRDO0qBEi9YB9zEYLBjOKAKH+Wp/4MSQMq2735E9/K3pUaBvuBMFHPOzz8w1Sr
yjy40kl3WyalgbeeF0aUh1EHXTctuaddSXkj7OkwuUHR21Mf4+L4DgFNXNMQpZ3vEisaHKGHXAXf
GYlg6cQG4megHbnLcHAp25zQaMAUWrjhA0T1mugg5dLywTy1+gnrYmX6knsjnDTTp7gUqaf8Twh9
xC2TGQ6fx0y6ox8ybFsAVoklvz73WtxTaXZOsYag7WzmisXphU5H9qtgIGXZQKgHunGnbQpn9/KD
o7XyiFfvrpavdWqMmNTF6TvY7I+RB36J+kG3/L6HxWe805uJNiAno4aYL7BGCAeWarE/yKKE89Ou
0fsZo6o3WEnzvwMC5+TyfXpBTIJ6ohghw7zT5leJ4Ouc6yTTRkp1vBkSFv0W+aS+Eq1MQO3v6nIV
YasEBFf2t1ZMpB6itAVJKvMchIuyjYpoLvt+ZHGoncfKlNYrEJgjsDnuYdn6mfN+/3JpNx09Q6Xx
97CA1RKHF2AJK+DA9NFaOwxD9wGzIEojNFESkL3oggchIK2+GPlAy6narNgRsnCHNHEdaLl2nftB
sL+ktSImBQKvEzPu2NGl+waqm3ITsuDSiwiAkQg9CKYKJeUOh9fMsMjV8k81kexGeaEHV5v/sbH4
lJq4wwspWxmEG5SLcDm1a0uDlVIXOaRGWZqjyHf3D42ZmrXr0C3P6PCHhqu53xXGWHVXCDYgv5Sg
YK0N2ktePMey974ydOyhmNYhLmRT+vwc4AV+QGhnzgv/BWNsh60g7eDkzpBsNRqyxYhEQWbOZW2V
Pi9U0z3w2Qzl1LyB5A8yjRzpJscGweoCX3/S6vF6DWuIIEewRksilK8hcSKaSDmMqvqZUrEGSXCd
aJEyXQZfSWImD1xQKpuWZA+Rxvx+M49BpetQgb/AWyZyynZW6eS+KyOa/flS9nhxp6v/Gae2ak3O
TJSFxghUrK5TKkJYfgVOpH5Kqkw98jNxeMp9VknYM32v6GY50Y1/kkzguzrXtegg5qVNpVvbdQ53
va/sptdUqDhPfgROGD6gc77WFl+KJXFM2oFWgkn7Wy/TJsuYEVL44ZihZMy1qh1D9cv9p8RyKE0A
BtSH+eGqAbe9oYLZAAUK0aBUU/cFOBO6ANzLc6Gf4VmeTxs6IRZCqZ2ykBSw/0VpdK5Q4/X61Uoi
0VGHFgTBd7FT9ADRw73pwVOpU2brxZLFAoX+z9YRQA5nDwIexe5MUYb2WoAaATjKfzkCTWy9a84I
afYyG2PCT17eSWTDqgeqgA2Jnul37tgLh101beX3mwJCTlKGPddzYYlAH5jLgaIXRkaglHeBVAPC
tnV9JN2R8VHS7Mp3UxVzqpnO2QHERXnOozSWWb3xXYkKZK0R2aVK6YA8d5y0fa7BhkO/rjptu5Ya
YTgcVvG+FmxhNPmB3RJrJZxQ5jjG/snloslv3tyo4Hwx00FMCBtR9kFNfooXlzOGBLw5q3ojDrJv
Vzhhj8K7CZWSNI6fTQR83b0ezWoHAyrXULGYVLJiOTV9x+E00BDN3MBdGaPPzzt6AqyszJM70YI9
AC5I2QQdqqZxr1jd3hc5PAnICQRjHOFriLoBwgYkrTh0LmAuJDofabFDmSvCgzvaYmR6383PjbVe
MAeEmbuzGUm9++8pu87oRtsRaj2AAr8gLnjFWXvcLE4/HVT8Bxwy2V7kFk+GJwwlZ/5xRmxf+jz5
LhXhKe88gP1qpgmHNwq3bVr0yu2TXNFsVyKN/DgXm5Rt8bfGVlv2Bo5lJfUkazqZj/Rt+iamFJzy
PwDSZUHH7DL1HgnsRVpSE6i7jJNkL67FU/nlCKiPDXAC4Zbw0X04cVKR3XYwFiP4yDKWeyvBUmI6
uPk0/0T5/kZf8Us+lH2ehNgp2nYJpC0O63Vb4vKVRSCRYdeKlC+9a+myLNv46Lp2kqd7Ir3rc9O3
vdOEpedoaNjMWFhZTXIBzH9Xpq30Gx0NUkVZikRwCh+imREUU1oTwfLWggwTMaWubneoMWE6W72K
ws+f7gV5G67RapoeqNBnBvBhf80ULl03a6xqFknlVdh23wJTTgf07Z4cEtgUPsVoR4r9rPeDGVfm
ERz1OPzTyriwkL/xfsE1PI6TNjSlc1VIUtJc2ypLzaLKK5HpStQYTWK3SJWhOZ0VaYh6AAYnBU+3
zDeVlvUMtOJO61Jg7u6EcTlAf+6jhfqM1KKBmPuLwNtbxXoE2n0NPqMVSHt7JwBibJPS0KrTP7xF
QCZMjcCBwGuv3q/L2jgF9uQsmjMcLvgas096dk4oWPTwTxOsNnFvyCWpIX+Xnee50hbOv7dvQ+2O
CYTBW/Xe+qHPKV7mO7bERhNwT6blW7XE3Vu7JKLfZU54mkqiGlYOQChziNHDCMCLmzE9D4WDU+VO
dRmXMEGdqqshGJ8ukUApHA0PkBv8oSHAWOv12ZUfrztlr31ocUBDqcWNaScVAzoWX5QdbU7CG9vP
+upbyPla5XCNxZ7vbBgTXiJxmarikndkD6GJbitanRk67JnQjtcM0J4rct51XevE5wUn60dH1c9n
hXY2CALaXSkviHrBaWRi7aaJwVn8FQ++bS0zgw84wV/ZWhQ6hP63K0FCLeFK6Gv90J+VZ+XV/Kle
eWKmJZbusUkhkKqn3ikVWM1c/oQeVJkuQcjfJ4xPYZqk+XBPL6p11bZgvm9gse5gXbQklnqMIYA9
D6g8SWwW7/ET1bMzGOnswjnHcjPOci4iIupa/9Y+ykTwaREfJAKCPG2rOQUm4HbK+3a64+543yX5
J4oqEbSDHXTQcvITqR4xKIOvhnoeeabNds/3DsGLpRaAPWyaSU2YBsMqSoNUNLc5/0FKMaRtPRYZ
bk7EpGwMCx+E4GVkRepsuWLUv2GukW0aCTvg/2lsIafXaBmOPYLpdYOg0dAG658tiPa8HG1ak556
N+Wpw74eCQ0NbEMaKY2NDpCo6qGNTcp7ykIO1Tm8rmJQxt4xhDxuZ8CYRshcaRbYYzoWGF91dpZn
3kYwaWrWGnfe6/4PfvIld1h/KlFdAHICSQC1d16Z1dWVggmhHrQgG00RRk+GoNcTCpxUCeSkWRHw
aLDF+Nlf/WzgcFMQD0MzvdMHVxQxhIK/qVe/kLFGJwPlo5nTMOIMmqTrL/jKLwpzEvbWu1eX0d7w
ve3Uo0IUzRTypglPefIBSnm3iv9Pm+RV6Dj0lqcGGTfEDjf+GADPl2cpiuYHGKCpfIT+a8CnS7an
YIpwGi8jrw/3iZeC3Md1L416OLzI5AAsumQ6WEKzfQ40TRHMMGa5KyQTtcxbRawrvYsSHkS0uR0+
AE45KXumUxrbKuW6YVEY1Wy5z2z5k12ujIOU0hqtTCbWf6gFlxrHUX/Kf6QfQ4VeCp3iI0lLxUNl
CDv6BGslL9v7S3Pr8bEspgcoEPa7+xnJX9tz2VeCNtUZ99QBb+bIZVEdEpKYVAdeWJ8kzebby6J3
j0CMCSz1ODZYiRkqXxkZ+Rizj3xFRl2R8j8HNpPdD7yPEAvvBQ12XMibzkCS/x6cVXYFQWxzSVGz
5/TpauQoHY9KEtg81N+6b0cS032CBW1VhqAhTmtSsCuJZJQ7SxvgV2JWrqVSF0rhYDgVR6Zf4KfN
vHZSoOvJteYftH5SDzj8vCNvPpB13XoP7RGQuryVjCQ2vMVeBdTt4iOtLBCVsQwtAzze+dQw+ZAi
0N2BjBk2eI8JAtshFS4MR4hLcZqkWs3ArGIntWbQPdrBE2A6tVPqt8lLo4yizKexIYYyKGnUZtKN
BpgUwSz/y3Empw0e/cTtZFl89OzXqUk89xJ2WKXgHrftFB4LpVIgaPAz6xOwz8nPzqntwp2aPqBG
3rXjZaanvLIswmQiwc2kMO/AieIP6JgmHrGG62Yz4nJDtNLPl35kz4IWh2KgsWFSMpXUrXXiMJU2
sOKF5JVB10J4oXs6Nn4yuuFRqp3c6V7chubr3kKnT0Z2oGSI0N6Zj6ZATOQrFVDFLuDr8lUBBadK
XqVulcblvt73F//KjtcXu/At5O4PRxNrktHRTCrOZl0CFHbW3M7Olh7eIT7JwEA80tbRgKqpsnKt
5qzM0Sjy/axIpc9xDZVayS49kxurfmylwZh433nu2VEEu/vBtM451z34kKRbgPG/yOYOwFYPKbmB
No+DzhJi59pgmjxyLAqyhL+V8aJUmC0uvm8sPwuuOLAHbLi0hu/6bH0kAQIJYPsqoZDC26sYzLrH
NW0iUYLOPbtBfx/UpHdmoQoNpnKeqICISRzlaIv0lrJMp4Lu9sp78JICPJgE9Xhw7qAhnWq+fFwL
8tZMYLkFsxw3oKkMlmwlzFLSJfSVn5UN/dtYjJJFASRjDrd2/86IOg1ENDJADVsWqc0sB1uu96qe
m9cGn9CWxBdGHyt+k4K6F3PiliSLInWYKelOgw6JWeklh7IpkgTOFW/Ib9HHcDldjLJLrSYfEy0A
GEdVfPL7yxRWILnOSoahBjpKql4N8jLZ4Vxd+DV4TmD9RJRIhjs1+i+uYp2U1++ZRbdTUxaLmczM
MigGM/MjIhV2wUnbRAC6c6TYh7k3OEB86UO9X3jaut/A3TpFAGDIIsCSBHiivVLYB04ws2Al0Mnz
v6VvqJueqIwxfjAAZuWFTLcN2n6SxSjHInneAUYV80DT5GuJgLGy/nED5/yQKk5ehk/JCgeKnDgz
D64LgBpzwFUu20hmGJhQdM7myQkosHIH5934+fiqJCAcrYaEx7wkm0t7DcMSjZfxMRDTSO8VpIQC
DXZUlDLvobQ+bavM2al0fO4JxEKN1VAuSEqdiRp1vn2qRkjnNcrLnsZdmWzoRj9FVakTi2OTz/aT
CJGrWT2mQID9W92afeHyMzdPHeFGfu4ZkI0skDAswqU15/xDVmpVGHSJC+uMErd6Lxez2sOGjvCZ
jBZSLO45ziE62f0WqPiPLyoLzDB38Vb3/B9F55+QkosrSXbQ82pNyUljswQBTXgT/8x2O9GMaRHb
QyNUr1i4ZqSuBGRlOVKu92XmoqAsdTiiYVpmi5yyNyrqNN64XIengH/qRnnp0PF+IL6OBDyGRes6
zo4bbMMGNiv0XAR/3VVRXArtgFvG7rudMz6t0uPBKH2iB4zyvS+1JaRFuVPxvUR9lF1bpUAMufId
+bnnETXD/OIOSANjzmtLQXfDy+q5ZckkZXICzyN3LpRgKlKeizQfDoM37SRvDnqDHAl+tZTG2YdO
KECIvAKnSVVfBCS5gLb3yVITurN90TcAHM1yvYs+vvCqnZHx+EgRh+uDr8FgUuQoxV5KDQuCkQiq
JB7aalgPzGF8oCVqXf4lkpkY4OkswArh2CITjAIX0PkZfgwLfyCSSAabHNrbkZDGQ5wfLw9ezg88
pnsXn2dtNsDSPu18/YguSJ9E6U4Tcayy+jB0lkWTQN8D3oC//TAogLj8Hwi96hIKuVtmgiUeIaMi
TSwS2psf/zhqEUwegQSWu1enKgdPWUpWpj6LJ+6uG7wbrjHfJKeBRzNPMX+QhitSU+OTfGdftL7i
oHDpozET0f9lfOYsVnNy6GeRktGqwnoCXuUcp63uEOIQ6YaokklNpAlkFiryndUgWga37gA+Upob
uHZB7OK2V37L8pFYSTA0EooUoWTpKbpXcwzQ0Q5CzIhYaNsldqvdW535IsWEPjCd9j8qPly/CLqu
2qI2NcN3xH3xakytl70teFStsEOJd2C59QC8h6TnN6QsjKKDDB2I8NxzctnuF8vV7c+MAL1gENCT
wQG9GtUpaI+nJMcGu5bqexiHSvkbTUftPWEZNIPjcOprGOR8EJ7lGdziBI6B+QzqCGeTPfu/Y+vu
4Q2J1EzQuEVG0Cfpw93ZHP8a+DbG8XWoKq2pguSPzcvmoTMZ6G/DtUQIBjQXS4S4vxslj5Epp3wQ
RqwxQ6m+Z9YkPyrd4Oj65Ye0w/lIBsFOBFNG0rzcYgFGbmM3QMF/HomirM8TWKAoihJ0kg7qX//o
iXuve228weSYsCfoqElpFwroA3mYqANhIIhlvi+1F44qzJ5I9lMUxFnNIPndKkOgCKoJmjFCNo7B
9WuKodw4FqMsvU7M0Z6C5NySDs+vxfh9vsoAyJsgrHfDjnlQdxImeG2mjxebbXos4Kyjbjaq7jg5
XZtWx03G7WK9lFe4d4RrM/QCkQcgQX6GamsmeEsR93jxwolb4yPdQ8odjybGaSPYajaV4DoC7kE2
FbHnnUljfwp0wbNFYo9GEu/q6wkqn7/RstvSa7pfY2i6NBLosYXXq4xZ3n8cQaIgmMJTkM7dyuh0
eD1vVt7L0mWC0g6Vt/OFP/v6tSpvjIIn0/y7PcwrXXvxMN0JOvNYQfdRZn83mTlsmg4lc8mB3Vpm
5/TkjWQ1qsFnjkV8VwC984/vCM7BZGwC02VwBPEDG072EzvLgH976wcY49eRKC4HrHld2HZnMqCq
s2YW/5DTuC0J2ZRl5TXpSDEEFLRid4nInb5HoQgvG27xefjKi8mNLoV81eSC8M7gYLP4epgPwK8+
UinQ3M0NvIXvkKGigld9V7w5voO57qI8nEJU1tdhLPFcaJL/kgfZ0rTn5jRwXiL9qUaZy7l5+jfL
YYnHgUIbQFr+OmDPREXiLfElYdYlnuHQaSK976PvriVqbeBrT3kwrI0Ip904J9/atW3whFNzs7XO
9Lor87IT2TnpXZ4IPPLQZiAQY50gst5BTery4Et0lAICGXNVq0enYrPJ0WpP9RnwPDXTKv28bfmK
VBiWc99IrgHCYvE3Ltaa0fuuhilaX1nB5UYc/WsrAGPmCwLPpQ1Lg3Oi3rz/DGXWU75pkngAclLG
bogr3pdCwFPbcH/HBZ13edaUn+rbqM1yrrxAKtKD3BTtV/88vXsE+68b2y0PlEMYWkzpXC7avN/H
dQs6eb1ojwuRORAch0rsaGWE3YurAhbSwRFydlWrtPd05h/f9hnbAQYcdGQQmps4JN8e53NmBacm
PFve02IR1Xx4G29GPMHEA7hVXfARUNfjjUtWv9auGFqyWPdhFOH9dzTzRv9jNq8XjOei/tA57ejX
6IniXZ2fVnx9LgIVk6F95Rc//TkbUz7+BTEcHZ3KCs6AHZOLDSm1vqWe59agxa3DMzdIfMnwJLF7
I7vzxHmoG5/GwsJQf0cXoGuAYWNzy/iTyBbjniLtKlRs3EII5vYyen5WMeFo0vawznag0Q3JJkCe
rDrAa1TNMMWi7DaheszW9XSUEOb5xH3XF5TrBcxy02jM1802gCDO4cq7V8406/P6kqAWoVSmjX71
kd5xYm2ALZepsa3s+8isJcGh5SYHxXT/Gcm42OF4udni8JCTbFDRyXCnJeZf0Ohr9PUoRITweOpp
X+8hySTmCrb7Qs3BvsWK2BTeQKyavk9aUIgfVt1q/P3ZkWRFO6ZhPU9GX/zGRgQbjd7pF7iAkBPl
fS1epVGKTLPhp+gGFaw9n+y8n/KXyV3PkFlwnAevWEgMt/0liRrlyELbPlxfgphcmwKFpitmMEgu
GMgUzx/Iljd51D/WsHAIwUcRlqLna8yCitxu8+QYINGSM8ivSii1W/vIsFhMVqdnmgUd9m4V+eq3
/r80POKDDHAbi01sTmOF2/iYLMWaNFuyDE0kMl8F/IrZYeqz66BZfqje/202mzwb1ApqPFOjKyLJ
hYAYW98Cy9LDYkPvj/8Pkv92ZGHWmiUZW1+poEOOimLSDid2K2NWh/6UK1tAkqnfHKj0JwmlwbW7
d226dDqsF7bKjz1qKfEr83WtV9Us7LjqJqU5m9nWwpyx9zysBMdKGQConiDq7TzaqSV1dHVCz1rR
OVmBjFlnhYbN4zsXD4U5Wdru2yyPMQe0SCOOJ29nlF9cBhIHNOdOhgj+KZsl7hYjGMuAf97h7QjV
73DHeiDI9GvrqJMhNmDlvz1bQDIFYHrvweP5DBDW6zgOzfuuIhQqakCZnu3QeqK+V9ZyYF1fiM+Z
S8hpBkeiXRdjVx67N9ppDYMJba9FEnuFsZOPsLuQjRm/Nrs1ZHwFpUiDCLq7JwML9vLrOg3kOb0b
HN3zWk2/6z8Wq0GfG4qVtDZ4DfMoTEKzydZSSdtf7lAybgZpIyXGvgSVZm+Tbo1zl2Euw3UaQxWn
1R/X/jIBqH36TRUEoHQ1CDyte4vTk/pYo4Ajhk/YMr8XfudJgKKgjqHM4WUyM5gZo6A0H/qTbdpt
7Bp8ZCwP1m4Abq/lYBngR2VJWeO8VNIdg7SqCIwhZa2XD8ARd/9QFKPto1ldA5//6ONT9GNiS20A
wqNuBl8CfJJel1Yul21ocbAOljAt5fBLGJzck5A+nBCeBsS1HA+Vw9Oov2Sc2GANHKqqGrgxDP8E
KZRc552isVTsqcc9jPo96m4SJk6/d2PlLTg+du+zo543w71cBWE78N34a23Z/GTgxYy0btIJd3ud
or1PkNTZQFr6FwRvQikST61KYjq//S5zLUibecaDa8UO2io4d+dTPkuc2yhZloeEBAHZafECGxr2
Jakwy0H2LajpEn/CJApHwvioF6thaCvjJdZfnk9g8Gsxjf7CamvOxM8ZDi4tDAbCm7J5GU1jYd1w
3SeuzOTb/CYGtbV6UkQnbsHAIKJKQC9opXkgWsN5ZO/rH+D3Uo7XWGq++XYAIIPptSN2nlAkGK7w
RKi2a0CU9JmDyGZuGIQxagPlgoQ1XblkLeqIy4ZWaQJ5P5Zuu2a3+KV/aZKdwKnn+9EWBPKC+p16
kK//LJCyVki33wKqdVOoyLye+guNxA+L+AMin9uMeXw+NTqA6YubJbxs94itMYGnFNFUrcyNwR60
pi0QPHvR4Ow1VCbKzDFvnLlHBvjj+nT03VC2uP+n+cH4XrSbKazouyjjxIkAg1PJGP1NkVyT/5+g
jRzGIZOugKz9j8O6sb3MNAOi/trxlwnvfBHFHAwGfhdeXuwocma2jYrVmVxPn4BjKVjb8gqzxbv1
wJfbxCDMuoDz46JE8yAVuk6obpunxpEhO3/Yu+itlQ+oyGeg1WskHtnIkrnmixaG2yeQ6fJRzJCe
IO4AjuPty6xh3sF9+b4SOd8LFRQv/rAXj4hQKyMvr/0hDBbS932IfpiZTf4e5nlwkFQ2FymGgqSw
jvioPxMCWkeWsPRk8Q4SwzkMcu8L4cZWrm5PJaqy9J+Sd+yxuI1iqoAREe9MfVQIoadwRrOTHlXS
b1sBI39/G0XkfSHssqJX7mLK/7xIOViAPQJvyVNPozZL1xthNOEvjlEBWdcO0I4vESU8dMaVz0Ex
AXPqu7T6hRwMJnuq5aAoYw6RpGIlU2uYLvK2UwuvVWksf75hHzv0cxQUs5lb8D+Lt4XSwneSHorq
tKKTzf9wmLQxyKVfLGjlrOeq2RoRxhmwgtI8Y8LvLI+6k6URnSuT1YxjkygRGeQooJWC5eEmI+gl
4HnGkOuP1L9HmXfVry0sCfZQfacbN0K9xQ0+2k9hqa45B74NTkeKrzatAmnwmcVXP6kiStLSjjB5
yB5OVCMOYbM0QI39qHY+I3casgu4VhzdFeSucPFyXkQygS9AVPe2vBkOYEIXVI5zENh7RDcSFf3z
2v5m7aPsCyTdfndF9hPIN+QL8mFv7LR86czsDyGBtwzD4rG38zKnfbUHda99pttR3o0OBtfGWQqv
Wq6kLI0VM+XCsabiy0pvHVqzXWJaSDA20tHTAeC7VDCcMGvIg1zUfGjkOtfizVIREFix0dofygkn
dyX0Wd7uQiMx5qu3ae02fn3uJ3HDXzubqMR2QyJr7mJJtcgK8P07BQOjcRp4ANzKqVI65wRMwj8M
YPfH/EHNysiraowBCaDRmSlItvUBLDOzR9D52iQHe6GpwICpALNjBhMcZ+mURixHYz+ZzeZpZrz4
sVYZDv+Z3gofpj0oxe8xQVhzeqZrqUu6G3ul8mEZG8cA9El3/OIfpzaPYsvzsJKB9xdnJpDBLzeF
H3XbhjgCVJBsJ0ZufYWwxtetYAhT5suKiaWoEsBM6+Brf6eXvFQdyjc60fOfZr/OpRYOikRxr7DA
F5Oeq1YqtG6nqDMgv3CrLSvq/uKJRO5jbaKcWNygOcSCRSE7AGCzGS41slz5itBfeX2tnplvZyIR
P5HkjCvKO0M/jUaiN3GNvYQ6qEUCySO5qKUI1K2/kiPeNdgC3bGdUphtd4Tqnx+LAFvBxKrAl3FK
ge8sl2yWNLh2KDk5uwOWtMmwJq1Y4ZvOVLSwjyNH0v3yT0hj6pirEDz6oYTHRYqi6O6e55TdVa8i
uVPbCAWvU9h0y7HRslTf1xoOT6CZ3l2tqK9xe/DLs6C6PUOlsDusyZTF5QcsHSjSUX8iQIwxZxsa
h9/EzKHFgU/cDQZi6L7knzOSM7F3O8V4gPa84v3rNJkTg7MuoycsSI0p6B1MKq1qAyHwKZp6gXkd
kQyIqw7mmShXPGZlJUoiblpytoS0a+XFGU+WA7n7mSq36IL8SgAC2xm6y1gSW6NLDJnEaCcEpck8
AtLo/NPtYmCF1m24nl6TLXq2UbaiSzZbBjsz2mjIuK9Y3cQqmtk+yn0hPqMb7REuuGl9IafkzcEP
1eApQvhKkvIi8oYFwZ+F13drls3lk5vpMrkg7re/gxo1RRv7H13DpYjNcl/Zr2EJCaNBRyz0kmNW
SFanXbU6Vl6NF7b4WH60Qgu1BIPii1Y51iSYxTvXC6if765DQIwFnFjqVeg6UG/6kCDqPAFnZ8Ng
fPt8817XMDx+iJOCLIY2wr306AbA36RX3RgDAtWTfqbG0DNPKLV5caiRbKAww/VCoBum54wa7HOw
5/9Pn3vTyKMmYd1fHU/aCS/BM8KCzSL4v+rOBGSgxTffTALBw9vxPpaDgeQgq7OOvyUPG6h0921S
6CL0EbfKOoCGjG0x73dlqMGWnszZLQZJ8wKH+QVIcjNn+Xv/Gj/H8tCl9bCJQ5TL+KcSuBM1v5+K
+iVjD5xzahMjCBgf1SePntBeS/K1WMmxpSY0VYX0U+nQbT2dRWsoDVx58XREWcD1+xMzQJKK60Yi
jH+Fy1DQTqtWASz3099BEY1FyW7OwkFP3k95UQL3bGK1+MXppaDeCQigttI59mPO99mHf1fdExGJ
Tp5dqzzG0X9eRxUIg4lCk3giAwUBmVXqjFJzb42GfjeT+raX6JJNtRzi586EoNfqJC+SDPj5HNl3
0GFKeIwvL/rl5W82d3z6Znb+yVpiMw41U0OMG+Jse/dLfIoBsqDz607edtdeN/e1mgfOgexvI46X
Z0QuOsoYHDU2PQVEsRGHgdiFu5k3/twwdmkffICDMdVHVWpExnWR2ABRVBOwwpwokmgquJBgNDyt
BFYX05kZChjXrSKaxivYPd0v0RRpd81fKihuzcWsJTVuAw6Iq+d9q7J3w1TrUyNoFUFpAIenXanL
qTjIOGMk+QRImPwPLPZccLiYlfNo23h5rZKSQkJNfxKoHx7gjjQtZXv6DivcoFV+lvw5ppHtaHTa
/tmCDeA8L1KDLLy0el+1OYaW2U373ckRS3LBnDoBO7s4gzzDxJT7GbafH4g4B1qKIE4q2sGri+SW
mSHF91iWJlzosEy/JATeLGvVqR+yBFi5+7klUfOKEDkrYbSZxaIhEb+AP8Wt3dg1vnDprz6Y22pD
s0FfSZ5PT4DfeeEDT4cn7xRwJToK3pYyyaoBc+LFoGU2q7i2bl2JfabEf+a3Ps3bQGKgXRVAKlFk
2VoOrsmgi5MXzuMWS+vAjXMEs2b3krk1FkhlvemMYyCAGMN8BsTK8nZhRi4G8l27VGfTwIRNz4Wr
sEEurZjiR94ehtYnZnLaIilb2M1SB1fzb3qlz62ifxsC6w++qgkX7FTSl+vs5urn+r95u9Zicc/T
UX8cQmhvJmYf8O4Up1jE7xMP1b3bsYe9E/KyQwCffTzkd/8V2P+vI8FcN4+VQl1caTWCTPab8ERR
GSYZAhbEuc48yroWKriM30hRsEdBXg+dQ3uvVvyENF47XPSyMjBap0y1j3i6A1bOnnGGYDX9xvTE
jkhAwP+zA1UhqChIk3cmJTGATeedj97IX9YTdNpzrX4UgSBLzBs+fvEv/8zybPk4DEv42Nd1NVPI
cOkoOpagXnlErI3HqBfk/K71pxKCkarG7fHR9Wj1ylEs3sUGtDH6LZI5euulRuJIesAg23L20X/C
a3uxEh0n2HlslMdNP/KBT2NG8AR82faCRZl7Ka5A7AmyrjNkNczJ/Vky1iAdNlqbPBRMj01pAos5
Oke3H9V/OJ+RBFxZ/e0XJbiCbuewatFJy8t9WWFvp8N1Z3U8StJR8P7GLIvrRxSHUy0+nkc8zAug
EG0bhnHIwNlkCDzkjht5OxCJXQQSIFFkxCK1B2QWcZ1sT9y0XZJH+9vn/h334gGfALu17I8Kw8vR
kleAeFTsQNZ8+HcgFP4GckNS20QFDpizBHen58ik8oDjFbKtWtCiRWmL8Aio160GmuUV1IFKDtwW
n/ymj6CgaYHOQs1rrFWXVtjUe29zOeo/3fimPc83ktql2EERiPGtrZtmGb+OgLJRsdWUuFrZm8yk
lf5z61GlyC73ScQniHiisRGSbKkN8/ojKnfOIAYUHIAkZbxlKwlzSbx7+O0VqwccFkvWQIXqKzL/
rMmm4M/KIfNjqjKXkS+sZWLU7gp9NsoWat7k/avX55Aqfe1QUgvPz5UfNW4z4Zl8S4mytpO8RK82
1T3XdDHI023zw4VGAJ7XGzxouEPQPX5BThEIvkPeJee/jmpHDBCAR2piJgVlydGTskTeO8FaxID4
52REY766HfhHFYPAv2HX7PFSfA8fah0W33nh5ih4LC3hWttPyKEfJybgVyE7RDPpWFp+KFfQFKNS
1rhnjSvGKLja5gn3XdFLpLZz1W2ikxFOVmJLVpL4Lx1oV+d7QbcD8hUn3KIeLCF1omexder7BbwK
wuzOXPJxZ2e5U9plqs2GnNCfmGmyo1zQlLI7KkdYJpdLyseoZDIp7tdUDUXm0YJuPgaTzKSJAshA
LMyr48btkVodekOZLDoZ8gVcd0MmevC9bgnvcWtoz7IRFB/CfbW43WYlwu8aQdhJD1XOS1KN4t5L
gM3msG2rrrUzUUNnC3WUL15GxtOtzuazu8wwtEjukzbVoI0kSPdbzdpWrH4AZy5CrtROFd3dCibI
pIoNqmWKq+aZD/7Ueju6c/4WnSZ2rdmWqO8SqCrk2mLzm3/X7ibZrcrFdofpyMSnIPq0yQ0jqPh3
raQyj5AIY+4l/cufsAq/bR+GQVqLlnetBz3dqVmmGwh1zga32qR0sfj8zhhl/X9qbn4rmJOnLsem
3/ACRE0hgjKbxPjdLjIV0rgAa2qVZh1vMwkgiOXgn+y7qHsPF9Ex0YxeVcq9kBoBFZwcXPH27sMe
nRqcJBo8tR/jSWWAwClxNrzmTVZwS0em04E6tH+B4NFw7i15IjunJaOVopkit3f1dJQRmNecDEGv
syAdyHpX5zQPE8VEqCEFA6nsoXhCMIAZRSqAmMOPQv5OyA15ZRsfU5fszRR0Kwo/h5Em1J+vLG1+
ETwcrLkU4GhEdlf0vubkdnprvf9Efz+PYWjJNOKnsWdLGVDrvj8u7wnFe6e1nqDkx/vmj6f3c5aX
3aeZJdNO8eMyYmq4F83tF1kuIeOhq/eCQvz6Liq1w/EaekdT9N8EDISWZhzh9QbuPJqceiwhoxkD
n3snW2WnsJxlGzV3jIgogn018JdemJKhisBATvcU5KMn+VyqWuKPXDQ6UF3v4vEUo3XpdnpzSWII
syEdl0cUHFAroBppoMfpQAo1SZyl5nlsuVP6oUpe/Nfym3G61wMmgNLWImZgyBf/bSAG7UAYLFUo
u0FTjyQlVC22T83w4E1YQUT6Ylz7QmsUztqEmL0WTBuHDYZiYeXxDi69jtUEQJD6+tHYNnzMzzT1
/YeW3rVfU7KKMrrQ6X2LQXbEL11D8mabYtZqbIxiaUA8I1jTPapYKGVdaTUBdNWmE8uF+3SZES22
ugzdi9KRoPyLLE2L9YwnRK00XRtDgEHzyoKZ3XgAxgLGD37mJXGy7i8WM/XqVPwbEOgXTxyIjOk0
DdDwjEBftNrvCgR3xERIM3sG51cyz44F8dZDdeoGklRMjiEIAlZtCbNwTID/mQfwr1j5Wo31Adi/
n7KfJyKTarTcttlYspnTGF3R5NY6tIYag6nDFWJ8hqYmgDE1hSUlTZcRrAxwVaWaGE4izk6Kijls
ZXcasbCM884oHrcnDIff3IVKoIlVIwKGHQ0My6Q7JVW/vgc2zAfqx6DRqCOF55eirWAbN1ICiZZy
aBKZzXiLx8Te+n5NVqPWJdmt3hiTVWt2/B2tgjlQFZZ2LrcsNsfH1Gdm5quc+6+L0uSPngzMG9Qb
rjMyi/tRJiQK19PMHK/SUFIEQ0SZcocZyIpEtBsk5do6ZP2V+40BQBJnakqMniFo8fWzeoDGhUyO
QpHcrD6ikG2wgrJAkMBPGVcqxqEAzZbFdyyqek45wrHcfNeFA5JkNHTfVK/vsnG+sQ1VNLVMWF0e
Gfq6nkZiI2IwRfAoFhkHPrrY5c3QQ0D5mXECyLr5EG40D7+ncySj3Ua19wX19gGrsKHuLgUkU5W3
wBGg7+9ecnfWclQa/4vTAPDbEQtQ2eojGezCH74HQZoAEOiMLMW7/GCgoy6QE8LPquUlwL2zWtvJ
UEWQT3RpBFGrw8hACXNxgWmqxOb167AibFYeLi5ELB0AC30M/aVRAPsmgaWDteP6bJUkQ/ADYtTz
q0lgJOddujt8sa2mKeEM+n6N/tIXF+v8Le8brcXc7lp18yC15dHN6BetSyyPD6x2XDJNJh8AGYim
ck1iRJUpKEBBRHvxz7WTO+l48GkBkK33kbVwXaI1v8odxhN5Ms2R/Z7yasXvzwxyHfJchOJTvDJ2
lFM7AsxRZPoYHk//oNiwCNpksleAQfPQ5mLgua6nnalgeY+ARQi6QbwWwdnbWHL3EAqFNJrP1HYS
zAvyyVibmwkJfBogOMcDkN32qhTfukhQROCycFXUTj/tIkNB0CsGnrqi+imRJB+2NKIbFmKfCMHT
VXDVUyZx6Q+wLRRcqEEZxRAXx8+urIfdS6an42+yCrWO8XXMcFO+kpG9Qu+l//DZeV4Jt/wH+iu2
XhV2I3VyDkOMJER4FNhOcj6udFd0wnFWU1JAou10fdYl9Yby38h00DRTe7wS3Mn4otXB6IZ3yMwD
lic+8yoRPjBO9Y5K2PVG2XbZ8ZWdr5BOCpiu8t+KW3Ua8qFBTu7leNN6NWQ2kaMjDLRxh0z1qAXV
i8pfAycydNGb2eqwei8qWjDuLqDEAX6MdvSoBsKdtPu6LeTeo5upk13NYLkHRWAndpWMY2kRUgFK
UTucYh5dSH7fKHFRrHJaWSIDAI5aopGMgj3r2lJcJ7nXPF8SgUuxahhiriis9ED8VrkqGttgvGXW
YYGvip/aDsl1HboQPJXaEoWsKM/1DuZExa9Y4R2A8U5cfyDgq3pKbdu/y9HSmP4ThHxl0CNXL7gT
EkU58Pxsb0C6y48+jJBV83DIp6I5EYRs4ctFFM5aXDoHsNqBcdJj7lVPrO9h1l4SNEoycrkgOOxb
Hq2LAqWPxsg+gzWerp5jQNzMD1EmdLcpOTHW2ogRYioQZODGj1GMVoPw92SKwUhbnF2NQUbnA7IM
NN65S7Ei1xYtBGvp/3I8P4E5Tm3ZT0WwqkAFAS1qIP3ynoAZZkNt5qK0/dleP90s0TnrHF/FeSR6
SKzd5qAT+C38yn5yYInDxpN6iOVuGtp4fgHwO2M/x8SMS5daz/aNVzTHMw7so3usECydc47j3Vdw
EFXBtUS/Ab6WMv6YOW1oywoztZIjPnDjnoEHUlj2lM0aJjkTb3bXuMxm2nSCqoltSgAfGwqAYTUL
bHq2c3f+ubuPkGoT71fhHcn7mdI9C+EMz2V5WtycICtMWOz1sk1uUOvLVSJOUnIHWnGw26NzAvkB
kIPdtuRNFvB2tPhcD6HBnyWOqEB/folcWBrt+VzKk7kk9lJZqZQ8fpX0EKBQxfybz/9XtyOIO/qc
7AQdqYxzlHJXdv1W4ksuL95Q1pcUkQsxBniimXSKJFE/FB+5cW1DevLnTfFQcImNgE64NJL/MxjV
LjxvuVizJ0URMY/X5ly1wHDo3dOJ2Tz/tDlcK9cZkFzaoSkhykKj8Hr5mS2TU0UgsG6E9pe+bjsY
iI6k1H1IawE1klFeDhaA28s2sa9u20CgXMge4fc0Pt7K9+IjUX7QlPE2CaW2RtFC+P0cD3oE8SC6
KXtH9WPGcw31ffDgtDM1gCvgumNeK1Q8jbruXDPggmGi2k6qRJOXvrtilO6/zzFbTfhzl9L2460n
DTE9vIiqVec3ocXyLRiu3yslmeQKsrtL1oCl+DGejrHRFBIDEPQ56pKBjCKzVRcs+2DgJDw56F+o
7nhjNlUORgB3L8S2v4gBMzUYzPiLRx77lZA6gXofDNTDqVsaViMbWlyg9ovoq5kHeZVA36knIid8
uTe2QquHchKaB5zeVVI1dO6dUrR1CJMXnAX6Hve9JCLsecteL8l1kkraiSv64dn7EZjCl/wx2CJg
JNHqBCPLnwCix8TczK/tOZUb3XjnHzAK2KDOygMGaHWPgAc4pvsQ84DoOxKxwh9IhpaDSaIE0AGs
EAuTK7rTCTtOIHeIk70t5itBcT4FMg+RNtCFA1FYskWJdQBFCWy2w5AgbnQmQSQp05i5Ok3WUKv9
XhV2gLBZW1i1CnO/a5vMMIb/0UHCzZouMPbGDKQq/LhQPKwZPElVnTQ8YyGVPg7QicSaUxbiA2k9
xLTX91qXNu5M23/koKAeQlWQmKPQyMqS6IIQAUkxYnJVxHOhNQ4AH0wmbC4DRheBhYcWy97jM/6E
H+980z5GwGq9wp/OlIUgMYeTPkdqZreNw9KZI8EPYlvoCteTiP5ivp4KW6NRL40xRL5EiYuJN042
ckWEw5zWB9ycXeBG7SQuUm8H4eG7mokQ91wgI9bl83292eHW7zbJtUTHMHupSkfMzvJhjJPr6e/6
Mbyt3VXEVuMJyEXl51+94JwN0Y1f+HhP1k8UuS++5k92sr/QqBUiZfr1Bammh1PLktnCMLU/jZLn
bPdLd4Qr5n3UmzFJcwG4MNkNLVi9/oxN5+y5lx15gHr+5ZQPZKCjFh0rjv+HG4/mKEIrv8WSi+a7
BU+Gqsqdp9Mi/g83fLSRahqSWZen3oSYvbVhwdslPf8fpTgSyAPKLJ6vkuHN/3ZqXlKsMIgD7cfY
m4B4FVd8l3yMt28GsspButCn4rVeESToP+MEzLBihhy3xTg0gUDEPFKpkS/i7T3CeXp3l7EkiuR3
0TyYhUWh9de0YdNbXn7ZlSlrlr8TpztiXEkCP1UcyJ3XkOe23FQR2TbONz80Q5ABPIzS+pOcM7/g
XE+JL08CkLC0vV57NFig4il8FON66TRBCJXTtFbfTf0+HJ9dP+DyMmQsItLMxVtN4/qaN3lT4q8B
dJkmG+KPUVmtybNIRTdVDQ6Cfc3bHrOGzoFV8vodu/Qs9VFf9KpiikwYkJ2zFDQGkk597JkbrA3I
V6W9bk/T8E8sdhaTih9xLMQZt4hoD+ATT8hxH5+i9ljEqzasuQVKxw6dADC0c7gQHdsBDhfxNjEJ
b4ATpdk1O0Sy+hzbSdoCH0JJkAsWySOBLmEWgV51yG9HdhFJZZOvRhETV3h5ps3Fp07CRbDo0wpj
+Kgy7VRwjFFPwkjuUdh6ghIkR7oy+MxOFg9kYYNlzN2d7/sHzCf0V9mPhhs0YVyzLzPFkqdd/9We
JJDsW1G5uX9YN9BaqRQCuxcYrRnkGSrS/dmeskCERVABOVUs1qe0iU2gludJK1ZPnU6eRsNczbA1
cVOicPCHaFxTfjT7vC9RFiJ1kJ4fPYYT0HzxjRehzOBvwDfNCx5dZ3UK+kcI7Z6bIdt59CFCyfyA
7ao0OSGewkg8PDfRyQVDPLUrLrMKpC82M2MHYlN04sbU7FE7HRUo+4bw4UHOtz2pStnyvCIMAGQc
NqF5efi+/tZhPp9fxRi0xhwugvWQivBuln/wMKlvumKsKCWoxAp0CDu5wMvUBoDJyFMkfeYKPnVy
v3XaLo7Dub6lD22n26bFKzNdcqqgNLE+CJ8kUArChEU8sJRtvVWzIip+Av+KCa2MhKAzqhsY4hpH
GT/epVgqIi3jTFds1UVeWv6DcoyxNVbdeoqMlDPdoskaLHwrMeRQkAESI25eLSSw0D7qbM3kfC2N
8Mm4hAQTFU6yJDK8RQvxCPCSk/10oYK+rac1itYu1ZVJ1v1ZOm9yz0+BM/TqTDXtUGPQPvBUV8mb
1zgasnzMDkGV3ja22RxcRAaK4Rfaq/7kwbeYcOjkeCdFOKNN2k42a2ieJCJS7zHVulZjU103JzAh
dHuRDRlM6Hps87ZFvoIWGfkd2wn9q+am44s/1zqKNEOAnaS8kUgTMuZN+ORhJbe3qof1jylPLZVc
GRpxWQRphXQAqP1sB+MBQ+wuwTTxZhCpvi5GxH/mDSGKfjkZGRbHQO0y0ivs6sLHVY45AeZY9dKC
ggEaIqxzSWLAqykWXdcbg3gBu8PhL/0MrdWxNGmL/6aBjXOnfp/t4OsmF8HxzYfTp8DeDefdyayn
ZVq/yCfjm5MMQolH4TTW45sT5l5Kq4MxOYDyGTTsyf2K2XhmcLOLUnUDNHnDQhWtHuMgJNHH0nHO
DQgBPYvgM/DUA96DEOTar5O4kJyWI3HXADdy/ozuHKfvdKVm/QJwgk13kMj5fPQvzUddXaFZFmc9
NiNE8VIqg9y5+NJ96WGikXzp7s/gbYTrHoVfxVz1wA0Ir5ZveX0jl2nCJ8Hgdo/SBGkqmv0M59FL
SgpxCzlcEUnIu3kRwHbFIosb1+btwW6eUvRNyyjxiExkgFDYh0BDIhEDvSMoKaZEfRF3MaMTtm86
dF758TphVxoQ6eSoVJYUsBdZd26ilSGP8cZZu20wDdkzBZ+Net9gNaevIIiUWQCZSNMTcVM4deyN
elmEtmEXZI6TFyDDewN58kGSW5O5Oez33Vg3+e+5/AAI94GinBurAsIdfmUwWN1bEQfLEAIfrtaF
Gxiwd3lp7IC5F033VoRLmQnrMpAf9ITpHwJedpUvJluMeAwyV0oZmfx8Zsx+PGvilRZppsN/Fi+J
rnWisMNj4IwyoecNqW9iZ9/qOTzxz9FTn3YvUGjf8pMUQRBJVt5TO4n7eeqL27FUJqPBJXlLvH7I
T5MyYen0g370LJHaFkYsKvKcXCaI8upxUHAglVzwHqeylEns9DwNSn4ytJh7a+Z1gWHUinRYoKoi
1H4XK8C56DBe5d6h6ki6ZMZ7Cv8Hs4s3R8zo44DD5iVgs4/pUNgDdrpRuUtroZ5zr9xBBAXFVb5x
nMyXlIu+O/zafLbV1R19rAOsi9dTstw3KdFo3t3IfTfAaqOx1JhQdhjWezYpiandqVsJOnwXX9nz
bkfYsFOV5usCqs9Vn5481IuhgLIqs6ozjIMWyqgpMo6aClZt5frLp13LjfErD6M9cv1SzlUjlfUT
xPGmnh2/d9Njnn2Q0Mbr4EZn8Kgrc6cebjcOz2FJ5jfqWP3d84zlWM8YN81SikCifyNoM56cyBI4
gm0mcg5gFVM9b79dZZrPShiZ+nDRPb0TQ9S7Jxu9nC2YAbioC7sHG77HAMujZfrbc0ddnDhiL0GC
c0noGoKrNC53245w4WLsJ/Ep2O5qFtYMMPqRuXVnWGAgQiJJDaDk8WLBZXTo3szIOt5zsAbDPdpH
R+PwbWkvGRnnlnns+Fg4HdOJNGzAhFpj9Aiqao/7WDL3qpwl8v2umOGu7HhRIY8fRh+V70EoUuDQ
Da2G3ptaRNVVMCN2ZESpMIB9ieYeeervPD3KQz1Q5o7tsphDUP3talb6cnHAgiAecBQEi1725t/g
qPtP84gSPagyGdYcjelfO+HLs72v459X5V8SE0v59dGKa4zNKWICMx5wkm799xc4JPO+Cea7EQD0
ZomnAhJdswt22y11pQupwUtAGFPPCabZke5trwGCcRA7qsZ9XLlQP7gi3c55Pq1Ka72t5Fah5+n/
4sI8bdO/H4atokgz+QgXHH7dkN1SfEmo+MoI+URhh63bCVU/XLkaQdwUiVZSPePEAM1AzbJkOO4i
aW2+Z5hzYJqWeJDn1NdRsKXoXAgcpht7CrBInPWyLKQX74GyTZf9PJpD/YoSd4dN0CU7XuDLZ4hh
ftyY0t4VDVBiy9ApkESUV7mRhW7MvWONbN6GVovZxYxLs0O7nCio4Zne1Kv3aAVHLl4R3uIPUBeA
oANvZ5mptQ7o4P0UxeV/ULbDnT6bKDLO2v9NmrDcqLvF9S3DK8gswwG/OdqZ3al+AG7ecZ7Ja61h
SKTptjWe05EkDlv2xK1phSzQHymFBfjzBJaNkaDX+zvaYvqXQFxckx1SM0aA2vqvbzAZVbmNcS/Q
AOkNqcocptiVlchJox5xwRny4qYeKWqb7NULqYy3Qdz8io//t7mtgRMxfc8YpSxO2QHA57FJM89B
U/bDSwIgpOcNM4R51buoHLZNzNV68eRjH0O4UDBA6Ar/C8uG1BYcEkd+HYK3XHfoIqrp5pVvqhbC
qrPEwFFp4UaN2tG9fJGW8jfadW+EG8auO6wNT65KNHJMGS9fOQ0IV+Ua2nHjZUNBOoRxztT8LhA8
NFZ1tcfI4ndxZsCCc58Ur4cyEc3xSLYlqdoT1WXzRxq1eAvWVWPH4H3+d3vcYNIsTckR0Q8Bc3So
+jAstBSYLiP2qthmXwgYcP90g0CGkq9WQJqEV1Mg0M67BZeQQy2Rkxa1XCCruwZ0NI8P4qrauMlo
Og6OnYIAlwzoDyeKI6VWseX2akh9/J+/ZgYD85DxMKQfP6Z1jLGOp/N+0g58DPMF97dsjjmDMs41
Iuybi22RbGlP4GmlX624vnnCV9i3c+F5/BBIGWhrnvZI36sUzO0XavmAhdbSNeEzwDtxgqdV3b+B
fw0BTi+HZyp5Syl+Zccg5EDA/0U6SF686xQxkEMM+g65AD5wvMRRJIRjp2/Me2+En8XGUqTbZsUw
DPUEicF42Vw1iJeYUloOexGRUYcVl0bebZrgyVwxKXnlUkM3lNloDC8xxJ1UTXx0sVn62OPe8wnm
4ko0b6aSDxF5cqZsJrAhlQRJkg8gIxPTUY7vH7yuhtN9e9FwChB+3hKXP6LCGgUIhrBmVPNQvz+m
vIPLc3Xw3ZH7QcwM4hIu6EJekQz1grNU5tuksUHhJbyM1/lRA8N/vTKd45K4j3msLU2TFLyxqSVM
c4LE8TAYKLbBLfl91VtGC0msYdr6dWSU3AXNgRCbok9H50l7niWwZ/HKLre/sQkeGo4sxqnZmxjb
3Dk4RHnanTIcpxAbq6r2MhMD5apqw5WScHyB7m2VLaNrrliSp6r9POpr3mhsIeUFERyciR7r9iuE
VyzwIv+ZbTn4YbZA16wblFDR/fTFavAVkXGY+1seZhkxu3otZ5KOqcCNFcAdP41ppWD4bfmpLcWC
r4iUInzeOSpzaM2zQvBJDXjLd9Qf7q13woBs8JHSoHwacernigmlPyrE0EqLkjpCKO92t1AnNZc5
tt+XSeHrhRNcF0KEzAnR1V/R5dRWa4H13A3JuHi+DIVfzTFCojzRYDlBB6aZ12wFm38dtuzDgBow
PGtFLYOi4FK+wLnJPYg2GUnKVYjeMHRfKvJfhfbwhUv3Vy3ImqlYGWTuGM6qyLBwiP/GhcD4qQO1
RhBUBuSLmxqM9LH3MSerBqj4vqKsrvQZj/+r4ytuUdJ4OKgBlojZhY3wIToB4DzldtZsLcnvukX+
6FPOWVtxK/YY6qCcwt/XdGT+K0P+mDo3J48MErhbwYW8IDMbYYthDHxs6Yftcf9lQFLS4SyJheV7
DYXURBNlY8PGwbXjWti6gC0E8OPgdMSCWyNBCTv54D6PKj0MQO0VWdJ5WkHaYf56HTd9uyq7laMx
5ES/iW5k0sTlCeX+5quEnS44DXJ/gi4BawQtqRimHloOy3MjqxBGpdw52EycAQuDpXBG5YETpXAj
O6GP2K8fIIfd588tvXRe/YikhUcf90z5Bh0X8hLShIzYbCHLNnzV3uN4oPElhjn3GlayQ9kbsd8d
vGpxw4izs4BQb4nRYhC1UMDwm96l3yTC/++ouOb8DpdmarAQcx6lAg1aRET27XqVc47fam4SAESm
PSxqfG+JbKqrGhjVMt2vqhY0iklxr+UkI+WqXBU4xWOWPadzHI1U5uK23XBkIfrVPrY0Vlzsfv2B
tw6GtQORioc+ADI3PsGgiI7PsJaOIpnqKT3NyB+LqLeN76QTQQfhM3nyPaBsjZTo8zG5iWnYe8zt
W6+wK4YZomgQl+Cdg9B6rf0GQZUzUwfJ9Y6IszqEdGTbzznITMmFlTOYbekwy8ifPYcgrqaFdlFt
KftMi/OW+wsAkSy4BXLadOjS2JVPkOt5xST9OLAd1vxPo+DGBKPKunR7NG5SaTTLy1QL1rTj5ef8
LUH+cy5OLiBRNJvtR8CLb8K40akyrXPkkis5xMfJG5/bGgP2Aa5RQVcqGJA+O3uucZarfDCFcTZj
cyHlqhGWt2rDKOSQAxlQwCsfODJ3SR3vMeSSv9xtulq+XgyH57aBNAvbCSYXEeY6PvYgFWqsgd+8
wOVBjgs2IphVm75zhmV/t2/0dvvCEeupim1wanT1yRxfZ10E3YCEeQUxbcxvQ2xAzkBLx33xONcQ
kAF1Pl3LcgQu9Fo+R/L9RH7qLSO1l1CRgzINjUj1OhA/0Yg832t7W+jpLTyLAy5+kcNDCKxRWQxJ
QWJS8DV9KgM6g0D/tFd0EKKsLv+tQIi7RMOjgAH3qiQsFEzYV3OcYi09iJbvDmaRpszo71toVY6L
9N0sfZyCbOZZIPM/ZNSku6lqxzsTzSjF17Ovmg9hadTHWmM6fEAWSzbO1LxrNJdPBqXM0+klI1ug
WZ1GNkHtMqcATHdNCRlilAcW8T5gviGjXMCnTuUA4jFwd2WBHZ99j/m8+GU99Jk7fsICqAiJlJjz
MXfrY8MJ2AcvrjAW2OCXwUq40qwXRtKrfyoaX/irUSPPWcJIC7S/hTA9kZvtD6quncxbB2dkwVwf
JU9+KEcpJ/XB0nF4KJY3oMXwuCGh4HS3h/Wb7Yl5AQPHgPc802IztkBEDNYPMmIdnmdhMUehpdCR
3q6A7zq3G17m0BWclKtJYZmUYP6w09Ls2rLHAS3/0SBi1Aou+lgCz4PwMhtxSS/Rb+8JHZGePHgy
NRCd6z1qp9i3IEOh3m5bKEwwzZUgzVhVy3xbBs/F6OChsTBI9SAbxN7H82V0wi89gDfh8ov25Tzn
NG5Q8w/GRnwWn8oYe0AneOdC4VCYVL2ozYAV3mQ65m4H92VOU00Nix5hY7IiW49WeL3neWVSfpEC
T310sU4pnaiaih64Pw6NpzokpF2iX1SxNoTFdN7HSwe/3GeFzRS4Uf4cxnkp7lou+ECPQyV8JJqH
dud3MHX82Gje/LwYggUMAdWJ8gS2ikUmdQxIZ58pPdAOp+m7Jli2XujPJG5ZvDofTLu85DU4XwnJ
7/owoZYI8zV/U3c+j5k8ErlKIm+Psl1L7WW/7+iuENzWssrks/BkqeK2ENy5R7u+14oqKw2TZaP9
pAzIg+SxX+FDYdH4M38T3EqZdzAsSGKZww7JwxZnymT4uBxuwl5+wOwkFK0FA/1GlXVY6h7tQxRy
aqtncUdLCKqc8wlc0veZLB3c5pvjAPC1w+97ZS0udpX/w3ejwSp5OTpN9Uqk68RbLAQsUgtAV+R4
VLejUX+uYOKsJWvnx9PVQW8DqZbqoLuam3IgSiPj6+XbBj8678NYBWbtWW/mPS8zsHRVyzdYN4FX
MXoky0AaA0+yjjWyr1r5GtPUsccL4/NdgF0LI8QUYTGpcisTE/ofaVJTvAngwXCJH/QOmsaNMrc+
iJmRu6xGOYYqv8cB0rnO+F1oBoLr0dY2ZqE1STrZ2am+AnQbZaMo8su6cmTpyP5YMxEcDJfjmsYi
Ipdy/2nnrBbWZ2ORKuztz03b0Tb7M+YKliSe2VDXml7EkawfLi8t/Q7HEwBAmfdPwST36Fl1NAFS
e22EqnIWhhUfcFJLYJDWNN8Spx0wVgD2p/GIpcQzTlE9Q+S6r2hcZ5iDKWSk3uibHwIFzwUTL49l
oiO/d/L5g5sAnBB7AZsdDhQ5ctnbWrJcRe2UwiaL+kobipxAHsgykCgECnU45uJmGnwg6R06FWys
ge0c9IJ2f7p8tHixIA1kkDXqhcLZplr0CW2dYLdv89ag0x0DIiFvoOeun1DceujgtTtDf0biStrK
kgBRnsowNIm/5QiAo7OCHgXl+5kmhf3aI+iWqWYM8OyGzJriUaabIA7lG1+3p1q8hrPpLZcvsste
DDZ7WGSU3ggZF0jGFelTTYmfckaZPFnhp8JQeyU3+ar1afN1+pHfX2hrGyG0ijYLGFBiXQJE9Idu
WbsyK8Q2etp6hF7y4/I5FlWLi93/RFkUp7n1Vy2AQyawKjaFZQXguQo3/QmG9x9hE0wOho+kwYEY
8xp7pFyeNcKAG6KCvj8Z/fXz1xTi0cPX2NtrQXgNBGAAAUiDzeq4Y3yLHZK8bdiqTHpXc/bpulAB
I2zP+BssweivnyznpqfBU0LKrPhoGtKlDXbSSv3tzIxSPbE7a/YhsjYxQ6dLCwOzi/aGHpa9g/KI
iYvvOZc5XN6PKlNcxKvM+vLuxFPAuWlLAPSaIGFzxB1a/7oRh6s/87FzG8tVNT9fHQQG7GVKyCSR
Mi2967VrbBpfAefVYrD9P9FD9Wfv1bwVN48AgbJslNQm1P2hUVW9zRn2SZ3pg0+Ljl9MFAMy5V/Y
0827C/+0aykvRRspfzREYBur19hXGnJIZEsBkrTSLBU86/sEuyrgw9rI4VGiN1djZmZsBKV45n0H
6mtWfu4bbvD0HbqHowfu7Ku76NMQNL+eYmFk8AS9zOVaaCtRNucwWZUh1cONO+IL/FQYw4QG18r6
dHG7RHAAkvU4VG4kQ4/h6bg9EKN8mE4GVxjVJM4NW02FcOnin4si2+E1Eo9OCfssqTJg07LL0NAt
lKlaP5umpeXpiL85eAVsnGDePtky84zv5elYQoe94aXnv3SEqf49L6oGGxPr8dk37x0i/rJjyvlu
dsBhJ8yf4TQM+nhvxp8KKpnwOFqdwnhOPIu97Zm+uSGIWELSh6201rf2wYr9M1jxxPQtjKIOZJ7l
ZYHCWCNl9rVc83Px1+gDE3XN9PnqntL5FyyYk+Ue0/zCNLy+26NASDSaTGWnxmKsVl6udMvsetiR
Mjcl1AdlKAq1UPGRES+MxuHfKA3hFdJGSevHYjJKMf0QOPezESJUTbZJ55D4kwnKZeFDJy3FtBIc
xd0pfOxJnBpwaU+UJPHi6niecaiEu67W3AvwUNCsh7X4Tegn/RwhA7tcHhv1xOVORF9/ZOrYHM1p
fMKzFW4b/bodRy3MXylmVBI5O/yx5HioH7+O8JtWsYrkGDpCOWq9tFmdIEEgY/n/uHlShmyM3ivA
i3JhZaTsYVrDt3ku8ew/1IV5Ppl+vh749KpMCeDyrdJeZ6FO4KG0Zg3stkMQ9PuxRp0LZW17QwXj
HYntRwUPwU3LyT+R1vT3xFTBaiNduU4RjClkOLB0fp9nD5PsJ15RkguuX7mBQlvpgTwU54qtji6c
PxoZbCxtsjv8iRT9a7CIjVZtNXhHBTwqn7PZHtwux1/6zF4yFkDMNFbxMwV/IxZ4DzXHACTf+7M4
k5xMvUQjMWrJgl/QoArA0xXrzlIxFpSIiwgSU0PVog49+CWFhgiFgl1zCp4JdZCwGbzwx/DyqnOV
B9XkqVCC2DBgY94G8KQY+uN8GUecMhVKMglJ+E3L6j2NEihe2nUhIdGBti0TfyUILCZlPpQ2ROOv
NQkosNV6nBhI5HtR1MrDFKAwT/FcLw0ONHAGcqBpEjsdyDy8Ug1H90vIt0ZWLVFJOCD/06Fn3v28
TVhiR68qTnJ/E6cnoPB4UWoRKPOLnBFaFUv8EnWd45iANevZDuJkw0uWU0UyPYBpBhkWhq33H6aq
3z2ik1a4azemWmzxOq5VG3XOdXqqK/S4CBaFBuQFUaPjCXH531yJuyVE3QLoF90oS5rk41eaHlOx
Bk4szAMGKiuI6csUUcSTIHmQ5hTAYKqE4T/Sin76lgbafZycRMsexO/UB6MfOHode+fA2vUW8GwV
leOl9Hsz+LbSEIW7h/pu8Xnn9r6B4+kfULCdpqZunGc1wSbWHZdNOtxWnDWtio9S6h37/0eOP+WQ
onNaOb6Edq0Gc4nPJBqPFrCgD2B9dC41/ltd9zqhvLoERwkHRkzDi931Oqbs75yLfaqXNmnQVfyR
BrYHPg4yo2ZAnPnWdyWgjT/hv4fB0FJ2Q9TkAmlMVdztxuWJwNl/osaFqN00lp2HClyqTVFu29p+
kcOOEb+loxdKpyB3DDC2J2LgpsHxQfLk0or2QZ2IlxNzvG7ozARR+RaPfzbIZLCXPT2qoSOpZKKj
UuTbjSuVaj89kbKmHSabWUKjoozVn/uKSDXyCV4KVZLOsXbX3KSbI6AyIFR/CjaEWpyPQRk6VXXO
/UE3uKbqrnNrwm0gqNoAHIZED8iOIWRx4G0IDlELwHx/awErc+xi3OQC3VgyOvnMwy8Wkt75EWDZ
3gNDNWg7ptHOQRJS1lOGkIjUxdJyf0/tjXGbhaD3JkX8w3kLJRQ7fGFzD8bobEqd4733VkMT691Y
X/otFQmV/IgVjvS13EdM7A+9zIX601Sd3tdP6QjG/qKYlovgOKEjcP/QekTp0vEOPHLkYQnCSZpb
f6gB1TECkrEd3fiPfP3Nku1/EHDFb+IFiMaUt2+GaV0QusF8ndt2Cndzyugm7pkc2/r64oAOq9Bd
t+1SQLQSfawfuJucSAp7m7R78kU9bShC64OwxMHopHxA5bOgr0ASGwDkslIN0SL0yxC8+mGn/jc2
w0G5N8nbbwhpfC/HtM0Or41SUgPWuYaTIhuYa4uJxaZBxLML7gKCfAJkHYFRSgOZi669mJhF+y5E
jHWyfHWyQk0vbn2erW3lsETWq0oFclu22mHFfTbSExjOUQmTH6xbwO6jVSK0v0Lxs5IvmL2KrHAn
swIQORgNlNPk3R1z3Q5uH+ZaUNfdOBiPJ4p39bmBQwy9dzBvlyYxRT87yUXnGJK6qDRwBai1Dp+q
WfIDesT7JbOA3cUU+0UQcq7PgvsZLB21h+oUewzEg2AZheB2r5RiIMwAx5jo/9LgWbmvy3W0wcNE
Es+FaW0I+g6AwVTQkBcOzWFTGKbyBRV9eF9Xgut/xcVEed0iBe6WWGiL68lSsaGwfnnRGphYaaHE
zl1zMJSkSJOD0+SD188AHAQRizYhaqVxSHRPyz6tDg+6U/xIa1aPthnEykHz/p/aKAe6FZnetJfm
QzzWelSpxMvhlM0D5VTM7Qhc58E/avLGF3EqM77qcCdIUauhI/f8MhO5uiSLT1pPnAgL+cqHp27w
xpK5pI5kHHDmDJjK78RqTcMutRaMJoX7ZDLcqYgX15PWSik8wcuw4KnAoUt42bD6+y8FNSpPtR6x
puzL9qnZ2p49GhPfSNYs9aiMGoLyQ5y9/Fk6U6o/3LbVaNNzTRiJ1AXJmL9MgPMxQdmXV4HJnzJl
ELVGubs6Q7mTCbQBDcyTOUFYzoCSwOTp1FLG421Cr/khAQRT26rG9tfi1RdCZoZKeEY9pJd4sib8
+KP2DDvYqwEtIbbTIL44c/NsTkRgotCfBQuuQFGjpDYDZrduDnASi/JaFp0kYIzKOajh6aEcIGYb
QRpVMXLOLCMFLq4WOAfVWf/00I9/9uTPLuABHRCXtVAL9D0O75AJdFMzJGxCj9qS6/D/T1XzC84V
pgNn51wiQseRS1QYfOCR5f9Ui0DNkdIdnQ12aX9Epr1oD/K8DwYz199kczoHAbvzQFhnjMflNsc8
e55OrTXCyryqOOPuma8l9xkMBiqGl647PsPJceWu0Mi8n6W80iwULJ6fasUz+xBb4ZoHWmxPp8nz
5DI6y/dykLsXMVZvYwgAQt4mux4NnEMTsKhP2wiYqYmAMm7Cy/CXuINX2kYO3DHa+mYhF+X+/U8S
QoHPOMf7/uXydJj2jNEst3sDYD+YUFyKGPdcVcQf/3GXPUXoZ/6yQAzRGBRLkns+bDszUyjp5JGY
3Li4X1SFahRZSAUGAU6Ek2QAwN6MSMxMCQyv3tE3l5WnfH5f6fEbdUtkYCc/NUTGcQi2ag0oSXqX
LOy4xUve8/bHVBEEqtCPz6JwMUfkF1CcKTnmPo651rMB4ZVDW23KGDwk7tQovHL4KldmHp6UuMSP
HP5ufoLEOQnDAjgyePiNtsx7nD40cR6ynm6g4ZUP9hlfeCV24I95MYtX8TMcYMis0EBLRyvRoR8n
L84ZSM40nzkGxQ3omEL5IufeI/U4en+RejBisIBJ7VzQYKJZWfZpkvSpJ9cm5zstQV6A0Xv5IWZD
x2DpUrrhGCwakICVNxsS85lIVXZgUeDsT0UR3vNNme9+Xfb1Z7ZmlwJUpR4v6SHAmeBnq/xRI1Ay
Uh6itUcKosZlqEloAOK4ZXsMrUoztwfLY4QnJeR/6m8oFTZzfXTOdI1M9QctyF4jMNcglGaAfeWu
KqbW737WpxQ2triFIF87X8OJwL/oj67Bdvwg+CbY6bnGVR51eJMBoUWyGv68zz5fPJKyarPI+59G
NdSiiWz69E1yLmcedwKX1O1BwsVMQxn5D2WFiqG9TQerviOty5qfizTefMP6/IhyJygqmfubp/Vf
PKj8U1482XyaeltpzW8qGxSoohQGdVsfr07C686bMKehRvWADJjfHzN0vtz2zm+kodXAvI/iIUmp
NheZEdmSz4tzltra+PUKZ4JDxnHBNdhUiFvvc5ZNc5uVdQ6WMCcnpJ+JYRjuVEcQNfFCQ5LZL40i
bOFAnPGgU3m1obUfpvE14xNnGdOkdIWcK/E+E+4zUpao3zzEiQAk8mB7LAUXfVhF6FkXuGYwVglO
2VqtWZKOCXIzb0h+bPutLilw+3598UVSvrJRfvhdh0uuk5Kjb8f8cTAtUxVa068ddOKlI346enGV
cdrM/J9xeo4bMddDf/i2O0cRbfQteW4rHAQQH5y2wrao/ceU6FD6Be6ztJDbyo7ydLorE0f2WjZA
EkrxuMLfHwAnLkhUWo9TxCd7n9L5kG8EXnd3lt8X3NN+ZTeRZtiLpECk4nhRgoES6coMAtfZoZNy
5+Yc+8SNe9lE8guc+K1PfkL3bD0X2vjrG77zfnpzWNcyEsW81S5ik30KhUP69YKmLo3uwJWvNVrI
Uz3H7Zx89vWY8GWbsIWno5gfTItBlQsbA+NwL1Z/PEJvn5iUUBV/vSjOQ8tmLstnPktWi5rZgqYQ
C4wPECRggG9OOa0FiiSc3L2LGx302wU4f6wsuGS+RD2JI9JanQD8Td628wId8tH136pK2HgsygCr
LYtcuj3kKly5+YZF7yXP8K6jaaCRl83SAc8XT/3ux4M44zxUe+MIvdzHhc5duVaKG4LEQ0JghWxt
2YfPuDC/XKJdsRlaxJSpJHft+kOz8JxMiWPGWhtwgq/5PNlKcFYRb5/ZsKwAAw1GAdaDTaBL2ex3
nYcGtErwGXSyZWsXUPnIiIj/Jb17D9BDL8jJMsfMqw+lbiUB1zkMR+InU1nyvE4E9avMxqFvAAyp
5MGHsrkbfC7QYWwZVz47sfmgjXll1oP8urgjw2Qa4ry65VURHexa3nyQ9DcuE4e+2/Cg6bak4hxu
vXnawRkA88YQlJqbQDrD9J5frOJVuSxrnMhkiqdyNoBpWxcEzCePg08TtFR6P11+Wl5hGidBQXW6
B+jCDy3lc4B0EReGBpMw4WfQj/M1LHqk0ZEe5mskjx11QJFJpzc9RevhHPtYL4Enqd621oJNmDp0
djH5E2Vhc+jUJkyi6kZnZ8yjyaKHwZlSEtn76EDZfbMuq43AifdLp1ODybSaZDPV3FvFI1S9kjNJ
llTLLGAy5ajoXHXe8uRiP1m+jbn8vmv+PXLGG99SVPssMAKiYy1nwGgHbMZFqS81SkzHBphCdmD6
VlT0tELBg0gzfl4oTI+/LOQ/ahkmoB7IZE1UNHIaDNrIzmDrbZHbQm4BywhtqawyHXNe3sR829nF
WkQXm+1XV2mhbMkojkglF2DMaK804qBHVhMpJlVx+HWGl7krR+tQ+tTnTWT5bypaSEg0kUMgJMw2
Ow8R93DsmN0BlBWrb2SGpql0qs+LKjASeIhG+FBEzd093afuwlk+GbOptu1CnNl48x34jC0noXlf
rZKOLUlCeASOio0w7mmYTCUnHVme/voSFUzkLB5go/Qr2splxmASZ6m0M3Bo3tFiO8y3CAKuZNI9
r0s4E/VHV3FjzUtlFoUGbYU1Ioq4U4JZDWVNj+1RvR8R9LzKBojkF68sW/2mo+zeEDIIaJu35987
6+QUZn7GwgqRkpE8weRID/i0X5rdH4m3GkOcGYDpX9nOVNFlNxpdHV9dMeKIM5GVmQd5RJ6Ubati
KOT7dBHQFjsomolGMtrZ2ibeERufyAYShlJ1qG4pxtEp893j8GPw6Hgv5lVQLuBCUuY/Mf9R5ZtM
IJUV2MMqcT660p/pb/GOy2R8R5LvJDRlI2IK6i3QyjGL2+Ckq3xgn0LD1yJRX52TEzEf8pYSf11+
xY3qFQK7BMmIn54xWA6rzAx8awscpR1CUfiCTwtkvIoa3vfKGRVeb9O4FmLcTNEkXlOdvM9vr2mm
W4O6UWNd94z4dmnGQvrfirtdi0vdqepzogdB1juU+FICgsxLqJ5TA7f0F19T26/zOYawM+7zN8xq
JIp+eSSOhJn2DXXhxMwIowPmAU4Cl4fQXIto7ES8Rjj1atEwe5rwPwqmm5O/pSumNd6P/cEiYd5w
hN6o2MUVmDj3YI2oAdh9EyqUI/tR6XuMS7FFViPXFTrxjfCke8n942+REy2OxmV+CJ5T9MvN8Doy
/iJsQPfltIm6Xac1pSl7calICEwSeE562gtjp3NFwdFd7X3AqG0Q4kMopO4F4ZxH1OUuxia4wyqh
fwVPKAg/krs8qeJgVf5DQrw3GXFzVnXOS9XOkMRON02nbX2sodAKmVYki8BaoHHXrSV5SPt/ft+y
iOi0GdOfOwK/VADuNGVl+o7vp4f22o+RoLRbOn/IJ4IYTOikAbur/VVQ6IULQIb6W2vDeqKLUNpr
M7rpKJhJvSc1pAZpowLkI7hzSVVnC9R3rIi04Dgpt58X6l9rfa7D2WJ8IdSqVSuJuOBT+eFzP0MJ
kYIO16xsWuSr7S1xDvb9bDeBkMil72z1sjddMcFV9UQtZQ2TNJPG1mZ08+AUfbbx3W8nAV49dpLl
qN8inhMh+vIo1Rn9rJzPKDPepoXfHghjO1776vGbkxv6wR4CwdJwjbq5QnDsRiAPLhM2NK3AyyeQ
ifsz341dn5LrDFm9Wkl7sS3zEJzWxm8xGUOriOS93bjpPIqOaKR2ny2Akdp/SI7D4jP5QOsZ1+iS
/XS+iscBW9QBlfmaHadS2VYI4vbsJ8v9ioqTuB/g1xCKimFBHb5Rz9DJPAxDMIRkrIhTUf5EsHgy
xlPLjsIymkPFfU6SpT4XcTlyjGjB1MMEKSKAJODo7jRKyNauhQxyAH04Uoeu56RLE47ST6G2SLWj
DUmrdAKTUTt7EMhPvd9c9sWgdB/+4HiTsnau/T7C8FQhBKYhEUsfgFQqlV84nsh1Io1UJ3AGZguU
3tTvOc8z4abpxQjOmiszxFLw4gWgluXeoKUl7lHqKtZjLcSIDRL3cA/pj21ObSgyDnkMEvgFNvm4
H2f/OEj+K0PDkJeZy0Tihyfm2uFW3aPiyXLlz6e3lN8DYT3E+ybuF5Y0wbZA7JozBIm9t0NQM0wb
ulnwSe/WX8VhDLDt7gJ9TPi0ASsft1zJ28FS+rQUe62OhltyOLTF5PQU9/bGsJYil+WeKjLndWx/
AtNCrsAByX1cZLJVNdWERAEdk3LdKxJ7oyTLFz+qv4x53CtS7udivgkPoNIyr6Lw9QIAMBimx84k
9Y4f0ojjWbyIfiytQ6VRKzkE1SyTlsvLEl3433N9cuIdTY8BKkmbktAmBNZDv2ch2QALlGFE1gIc
bUcECibrowvnjZkEPhBoaxBUzy7InmNXY/Dq4rfjjMbI97NR52gCUQ8DFwmVuqFz8t5HQH4iI51l
k/X2zJNKkQX2Em7NPn6fY5NT30bQVZjmRHGL/zSQPN9VjK125EIOXt0UUXGKSOvpj1edVEx6PuN5
rP+sxOZX4gc6G0Durxuy7FqUCnCADgVWHp0GE5pe9KFw+TE1EBuEjZt+VkluU3JtJQrvh3K0DvpU
6eOAworr5qlX+UX6w4soId24o+jxSXr+LWREunjm3IzORTtBnSwe9LHjKzeJrcudOqkvqHBjoGiv
OPWW1r0kuvi5LIyi/WMJEmNd/12FGQcgYJyGpu3awh8TCsUxKItufscAt2kKQz1CDN4GdB2L+vAd
NVCRJxNyj4smdeNM961NIZc3OKO8+EDHJqoG79LVZTnI3xm7gknr6vrLDzlrNUC6uQI8xl5vrIdx
FztazDMWv0Knn3q54GgXexNVDjRd/0yRU69e2zXvI5ArTeaThpORvfjhWme2Js9GoZ2mfHXGbkzU
LjR7PIgFrj+VDocaoZiGjZgILnFwToRsvkKaKBiwxhAeI49DpG6hqr3OoTHSR7nUFkKBZs332QPx
97qN1ux5dAbPBxEWci6EkZ1bJ1JQh6PfawL6kNo+UfbPtKzGYiRXD6SwWWEMChFakSO/kfeOhHZx
QN9E3ILrwRW/U4tZdCVOfnvhmt5n936ezHLmYrHjbVHvGeBmbfz3Feq68Fn5LFzAQoYmG6YMMmrs
Xh/81fS9kEHKH7C7QMSTVlLsM+jXJX7Y6cBaW+nzVzJYTAl/SLmm8QwOI30V65GKacWbs+9J/Wou
G1toJq/fpoAB3ZWNoesvGtiJyXh/ypA4ePY3xTPWYGp4B7UMWGY6CUkUAmgZYWPEWn2rl4IlryZ4
zQZHvv90UkSGKpbP+y+bX3ly8Rg/GFWGxg9M5xgtsBw5yKEj6lZ4DB9iimOtrWpKixuZvPWxU7jz
NJuQChxYS3gZ5LzZ6LCWOzUXj+c6jqBNQ+4mXZyiEQnxe0nuvoT1tpeizD6SSIjvGrEgv6J+VL/8
HI45qEYskDOOozuqcnrcJ3gSYsxwUU8QSR0OtqoxxWKGCIBH5pWrppzC+/PcsrSUq4ywLXSgTKhV
/Ul+pq+hbhyPnGZHXuuUGQxygpdfArVnnfRfE8aMXfdnFU38ASjw+pKZnKCIu2h5VvMCF135yR/5
FaUHTkWzqnkvecJEcssEiRCrHLAZXZpuD4X+NyJwahnHJ7ut0kletKUXZlsEgkKxQSTIoKbK8SQU
dnBcZaAmctSTsrNWFlcxBvDKDeV42DlTQb9U97mXyIyxegMcSuBA7DdCVfBUcucRFg1iJ/a1vJr4
JzIPzzG7RwLJj5EIwcys2X9KOuxxXJF1b7/tDeDDwOC43a5EWwdR0vQsKDGC/rlc2q/5/z2qWQVr
MwDFMaYw7yMQFdJjC5fsh9//cmhB+3VfnrqjqDQqkE/4iK7N+Gh4tkJJAUr+p0sUeVy22q4qpcDy
Go8qWdUiN8cpMZ1f40u4xshjHP3eejGuiuFLqSDUavkwKIOEcMi2coIE5s3pdwi5pjnu7S7Ku455
fNDKyvbb9GXP/CCOt6AX3Z1osctYzaQjSoc+RNQlYM6MUZqSbL0JcdQmZ8TEVIBlyih6aMFzlTb0
lTglqdqPJbn4GH6yZVFJc/lHAjko5LU89fKK0NcXUOBu5HmkBscioEYr5Q7LQoCQjkKBbQKwnD47
JFw+WEn2dmS+6XPpUifQaWahv5ldTL53yxUx88LCv9/Trl4bIzYc7JyU/wM0KaLTM05tWYx5Si6N
hAoBVwjmymmBB/tO8XBLaSl6UXNf+hqZZWzWbQSRb/hxICgYdQ8JdB1KdDmRt8gGAPE4p9reSwk9
hGbUM3R8FSsy86+Nb4riWe8+mcOl8L3OalKOl4I/slJv2rmAEQssB4l5COeBR8zZKPo0VbZ51Kq8
RVRSjOMw9sDXKEvwKGcRq3Jv+tij8P9oJo1/pmQ3SseI5c1QstM37ShDxbtnhq43+4wQanT8Q+J1
Nsm3ipVCLSxGLaJx2GiBMrHbVPeUtMTHa6RjIdBwrVW66xLcea9Rik72KSGWx/pyuOTQ+r6RaqpG
dhpjSklKDXeWwPCG8eL5vCFW4+nceuK5HWF4jEEY2Cs+WBqNL2UDOPyJ9/VQU/gn71EEyY1m26wk
xyMILqlW8L5pBIP6iBTSLgr1VQMQXnwXqWyHoIQagdcWRH73OAm++FN/sxh7rBRDPVa2BsnKM0ss
Kz3bB1S7KHNDAcTffHRrwNpLNVHH+JcKDWjkZourH1OxukzcP9Fiqy9Yd1wzn1MbqyzDi2F5dcti
w4GHh6tXxd9t701jnOayRYwB2D8LVLca/BP32CpUGMXhCEXFXxIAILOv+u/2OD/53AIfa26NWh6R
HYMDZXcnvj3SNJqJ4MVMjh2RgDBmHTSw44WMlrT4ceIh+TWwqA6CnEUGl20+yqRvyuxkfjXcoh8O
o+WchSpMrJfmkd0BcEFtRgNomVhwtAU3L6erQ0v3/gX7XTMMJdN99Z/zCemvrlyyqL/ffp4Ujhcm
lgmx6Jleh/Y4/0qST67sniVWM2ikKZwoit00hRzW6mCWEUt/Nx2YVGBhqU6px4NEEFtjEBC3K7OE
1XBNvPfbXkgRdE8NSQoDuBrqJat8SiVtbPaQ36hWAEWp7GiJQpP7O7rIYaeNrGI0nl9Oq1oNfpRk
jxeEUnBGJ9ALe6o02n9UjS0dsrPOYamIrPi7DOKTTGgiw6lj4jtNJ5Eb0leJhbs6qSxkR9KvRZVe
jOW5Zz4/WFcSc4/maxeKAWAs9XLEe3+HXx6zAJtIbSxouqpQkovwbOmn0h3V4UGmaJPv0egE7z16
hNqcRE+0oVJMK5X/ckF0oJ25Z1+niaP1HYNtiKzPyMTs9k9vUsk0sHeNhD+xpUFwX92WRX7IbWU0
J6HhCoDb4MOd2JsusWkX+oK/aGudGoq4ivjLJtSQwW0WTut3pXPeOzJ5ul0ojJh22MeZvaIDpa2J
EUBszfjT/r+yIr1xFY87uJEp4njy0MjWlGDH/pLaz1E3+d+KtxG1B6U7xe0Q4ohRfFHy+ZZTdcRE
tbEDRlsvjsFtbQvYeQ01noqADgqCIpI+pV6ot9+GQIxka4F3LMSXGAF0sg7h4VaxB8+8kvvzUPIM
Lul2s/TGWx5YsqPnTwGrO2ZQ1Ofv/06IaUq/S+/WTt9y6pjRcAZFqYPjt6s4X7sM16AIyWMngPGb
zlklKP4NU+8UkvDGw/QSLmgnQ5RlbRclfrzs+GVffrMdc6RonpIq2F5BvdBF9/d+I+jfT3Hcmc6v
3ElNESnnwn5Q87fGeR0RYgu1nOk/nE/cpeaz24wBpmAR8YRsJEgtsgLNUVhigtEtbUmGRKsWgPGM
uSjmNutL8py7UzHMOoZsLvFbE4IOMZ2S9KkeuVNfnNeXCkrWyymxYQQbsLniTtNTsrN7L6UOTQUz
UoH3mHY7X3DbEVbguinRapqasLxflNzA6kK8XiZ6QwGLWuGKL2fm/SCyZiloTcI2bjRfZeocrqnd
OKGtjSI3XrRc1cH8bfLZF/JE98+TDbqyI9ijWGJo2AGFY4ky9tFIGx4ObMY+tJSQaS7CcvirKgFX
AgRTKODvcL0/zHDqU7a0jHHjD2LLU5JK798TizXLeBrG/pFwq3zOMQP4wl2gVrRFY83AbuNexHL8
4GukIhPOEJ9HSxAFC70C12wCG6w9UY6lY+WsXBYoksbBZQvwykgVRzgdmXBKGWRPuSrHTp7H7RcL
tXZEr6u1xQ+WrEFy04GM0HgYVqfvscutqGBEh/HIeInrT2e3tko84q8u1a253yDy9WppevnELCWb
jhztNXahzzNKme7odnUlnlwQzgO/EPsuw8N2y4ACn5Lyxv+8nghY0CNsEPiPSG4oSc5VbQ3sjFDO
NG8aIDhQMbQiBuX1mluKdFGYELc1zoAzd/qkNAkUxwh/bfe0Tz34owLbNVafzBDt0tTlX1QD0wTR
t2KAfztxZ9+lWBi+ybPB92v6nc1nDmDj8Ci4lDzXHGcp3GJRbu2nhyiQikHf3FxRgBrN0RWdFkpj
vy3vTTVZYzkJqaJ62jcuD5CdZifB5Mdy3xOlL5gExas6mGiDPfSIqy/4wNa0b3Je4X05FKjFkFqF
eASZs4wUv906dyzmnCS5UXl0myq6dO5VIO7AOwqWnxZA6fh8iW8K14njr3x+wZkctqkgOw0Ji6Ee
3wHMRsgES7yq9RYV0dSnEQK8C0ad3WXF7zLxsudHBDOGIjdzsGmv+jF8bcL0mDPO6jzOnrnDDG/k
weOndmqaKb34R0DgIf9EpkbPet3w98pX15tP6QQnAxUQc4lGcnZVlq8pDVywuzF3OVEFxcJ/xVEl
tRleeKa0U3ON+dasZD7stpJeuNALRejWh0j/cSxB7XT3cxcr4Tsv8adLDcIT1+GTkmXGoBrbtcLd
oLbb8XHgwILvL9ZsVSYDvaG2YgyBjnvUQSnnqxJmxe2p1A5swHohoN7GXRuAs/PW9GkCrtUojJwj
8RDAMh97ulOmn8YxH14eySOnWueIsG0Dpjv68ABS8X6t3Qv2avRJojRn4PMbJAeghsdlcWf12Txx
ZXumGyZu+1gd4FW4gRvgXsTJoRaorV2MloGyZivoVj16EYQxFxYvuwNQuG2xbQgCwZ79BQxyEQoq
/j2PlvvRLcI4f+FWx7+6KMTwCWupNel+pgpBG7BrbCZDsFdGIjawTuOyoArA3hiDbH8Qz3JwtSDb
ZMBMDZInqyZq26yhsuTifYWAiQ6/Hn/gFSmBbb6jxbo4BoTr/cEMmO3pgp/814+X4OfujuwG2cuH
T4aRTK6spMSaq2ptMu9pxq3ZvhDepx/lrpDrhIocPu9YIQvmdupLWYpmgkYOevM9pJExuFg0oR6F
MEjNj2/d2F65t7YfdaP420LkFBANqQUFo9Idx4EBV8K+t4IkPwzOTgyl2zDtEwRdRprzy2elNnX8
LhzaeEDzjkwHPFLaEKYg1opSvobGUmOIOfsV6zGQUKQBmFCCeXrjElI+jgBl3I9x3ZY5s2KJTwCW
17GnLRqLBWzzwNC+Qnkp8fABjasJ/KEQVCITIGp8/icAdgGdlpOv+8LUAiORWQIO9+9qkDaLeZFS
tsgIVcxULEjVWkBRmwXcmWxdjxva2XPFTiiDgYXDEds6Wg+I0KPum0+CeavLTRqFIRCY3Q8GxnZ4
vCeaOucY0D3TmT0/1Jpvc9r+GY+qX32KWjizopMuWzXJwKurhXMdRwlLyNDnQI8BumA19kTpeV3g
56NkH0BGlPu+asHiWK31JBzJ7ulAMRyRnPgfbrncJW12cRlJzI6wShsFNsuQk3EJ7/Xm4yDoJx86
Q8PwLnWESiZ4Gh7a7kwi4VqxKFzVJq8cSfQ4ESTqN8qk/ZliEVlGiHSsHOl8V41UZPHuUGv8/APq
Hr7ZhMjTmE9FDY6BIU49hOAJEOAKQxRsffZjpVl7AWtsrQY7YEgJGvw3rdlYbidJvFxqquYBQKck
5nccQweq8cdJn+wFNMpkVfx0BZWzI6hoe0ydbjdx1BJU53HsgYE7YPWF6FkD6DSFhWRMkeiunNqt
lfP/rizHZOJFikuGBrTd33bI5F9Tw7bTIwAxLC4AGLPyniacaWXZyRU5S9wDifxRfsGS90T/5CE7
LdPHoTRnh+LzY5vB2lWVlnACSF58/MHskmmpsncIbyd6kYNx2wbmTqxry2txZFXeAarniKTVfHAp
ARP5+7TzB67/0vBm/eN1iOjO1LutuE9fwbOWAPOy9ks8ChSSczRmIC/H8Vzc3Ojj6yRFACA+X/X1
7nhc0QTq7ZvCb0VfaDZePUf6g/7/5bf8uQ+loszZFkFU1G5I/KkPnuwULHW2yLRggghrtA2jSq4R
LGTjkAqIINWTxiBw878nHs8R9l5qUuSEBtsAWGXGtVi3hCd10NyBZ9xAcIR2gxZ8mB2MK7agZ8PE
GNl4TP2CCp+w+pjUl5H/523w7P6XUypHSHKoN2C4EU6MTFl9+EeITci7AeWhDSzj+HFFSgUl+N+2
L3o7I9jXdT6m7vwhQ9dMWTTrrasmiUwZy0aCEbOKyuPkqpM14YvUkbrTu5onKeWtGSjzyt7ngH5B
gJPyy5MikHLHK4jA+Tza0PozFeetp2HuLe76LbHANUgTCuvnBDs0BMFq0a5X+kYAv5hyzAUOMXp1
9a+PBUkBBnnf3bWakYc3m8LiyF+ao7Lu5GdEzmA/9FUTmFojj9R2NYj9F4bcFT1aT/61kGz6CgEG
4Cd8/K2Jtku6NbyX16PFCgYM4vtoJvC5OlCz0w+jVpVcsXoTloFJm3cElKM1SkYuC30eSK2wXCgx
d0Z7niJfABgtCbWBFOeix9hXLUGO/PuBCZZOdkK1rRUMlRhhgKsCYDrk78bg9NhAhD/S+cmI1Qza
b/eKN3ZPY83eZvzX4Dyiwt6WiJun1/Y/afCTv9GaK9rsafe33KimqY6474508Xcs2iCl2U9oK7J3
Q3Kmlp9OAN4/Qy56GOh3nRQRnyAbzF+WeN1aS8phsf37Gmq/H9xrQlOOGi4sNXEok9TJo3OdgdIo
tU+tL9TaipVOHd62FA3noO/Vo8RKk+bBe1IABzsTdJR2fsSWzIynlAzpBbpyT+wWTCfSMaesHhNv
F7b+hxVLoOLpRj9X+JOUyNbV3zc23VBgIw6ThUWisOuLdpLQdsfTMz4h7ZzSG/Qe2ydQw9J3380x
+Yu3LpZ7Z2dQ4f/fzdZ1pRE515/eEkjxvWYQmwszkB2MAZsTpU2rLn21IJ+7+/Ox/4omBzg1nxA1
BYmG53m+RgdCgQ/D5tknMEP9/jK+3ybwIb8MxdGRTKgJkXULJlHO5YBOiHH4D1VBFEVNXt7IArYo
ytEVD2lu59qD++8tJNlsYBmj4A7jsJhbZHjwBbAKHH6k9mHb45fM/hCXd9wE/mR+QroGVKWR2oxW
NueZLPCzPn8x1BiWEQriS+dyFLq3lNo37vUC8iZFHHoqVJrx0bzhs8OnmHhrUVVgKEaiuqNy7g3a
GIPan9xc9yYUJxzkyAU2L7zOwtZ89lC/zlsbM7t+q2+NH/kT0W5Gxm42nmVyar3LoBHoczcqW2v8
pOPUbym9JQPL6ucSnPGxX9weZFi2A+6eTrn6V86q7Kg5GpQWNhFjIyaZRZGRzJMMbOJQoAww3ij7
F4WNR0c8f+Rh1FDvxHy6jmf0LlRjN8vADZ9eohmgFrJ+1CqsJgAw5Ap6XEJJldqnM+mTiWo9XwU0
inPMPfMLGrqTCoVpHsFQrsYe9V1VFct1LdAC1OALSUKBxKNl7d5SqgTC9ostXO/CcfGdfl3rRbcc
yporwcKQyvufrkQBi4/GvQCOS/6tKtQaqywd7iQCymRMfOeFCUlpXMt/5GarU+BnFchbWIMVPl2x
MmTbaT3CmHSgKXMPGVCMS6UXuMSl66eW9Ya0YGXTMa1x+jDVsmC4QWZeDmn+IM8PeYILnGGUKK99
S7nagKFNSStVCcJUZcNwG6V2jVk2+8bSO3fWzm6JfCB5J+eIu0i16EHayQe8tUcMEd3i4pVactjn
FYUwyG7WK+m9O9Zt8I4vLMXGZNbVvock01N4AQE+aZkanF4+6wLp5ZJMsSegvGEH8S/9EStIK29g
Ojg2cCWuoZxx6I5fzpoAGoItMm99WqHD3kM+EaC+VMiDXmphtO3V8KUQpnns0hvv+0yUhN6BZr0V
DfU67u6ufNLbBOgYgEmnIyUp549WUGN4q/mweaFLGv6op+Qcs81U/Mw82A3KzJgGrRoC6cSzlDD9
SQRx4wxEokdpQ+bJpRx/7RSm2e7R9HgxIk+K6kuJjEfAGTOrn43lsRoDw49VNfjr5hDYiUzs2UzM
EG5fKBkvOLZ9EVaF2gMQox5R7KhuxxG6uBH92UEQtgWN948OOoQ9Ze9BafQCqHlvWXHz3/Uo5d31
hQ93Fc2jWLox7y8CG0tOIF0dwEfWfYhnNu5qHwr9BcM6EF/iRojkNYPSJcjYJd+lIRyBsmT+NiUa
Hp8DvP8kFVhcfMI2tRW0iFfqk2ZzQYMEkVmJUOd4f/j11GRBZpyT9XJ3HdhDbDjaLKV6cKCjqml9
GNh/JnJD8CcycInIckdRiqiHtrzQ9G0NjYPmnhC5nIpqla7wFJ12jYe7MIB2ZdPMe9jgse7LrLul
bOx5yEh3ez4vqVusMn9BIoSkiS1jYE2m1U8+4e6u/IWk0dsDkVcBhHAJtBpQhYUgR96WNOJHQUP5
hsXgHNLnwXKTNiKIbvdxfCTOT5TSpiOspZHEq2fCaFjGnUni0+L9S+qybca3Gq9EUBi+ixmSsvJ/
TIrlx/TDUgRR7JFuKOrv6/0pz6gr/sKqEUWe8I0Pf3GFdTAJp0VZXX172awxQ3ckdTG4ZvxtMGn4
/zKBfDC6CKZaMEmIH+GY822EWiF2KI32MgXnJKvLWDDAdTjqdSC89D0/mB6dqKCg9XG5H8t9kPL4
xiMFXU5++Nirl/I0JqemU87U9gN2mImY3jwTRuI5SDuRa/JUBEkWV+gRL9BJLGtHEj7J6vxTU29F
X6lhAH7kKXhOEbODggSfBm6boSsUTrR6yOrEZsDEg+VcaXXHOMSRlw+6AX5FaZiyCGWQhMhXEsxm
hF1ELRZ2gIWL+5t/TfCthphuo4gi1Md8X6Uex3a9IsKZ2wfK/Io2DKoOt5P5ITuslhvCO8vuoDSq
K/1Y5i91ia7bj+OnJc5YpFHxgf9vjuoG3AXIFeeEgqny5GMbCzBa5KKlB20/2votT7nAr57n3UGS
ah8KBgXvdpgeCs82n7VQz+kZfCuTsey7M/fZPWc9tbAcWnKmWcaTy2Yty0ARpm3EYCcnrj6f/ZJP
7xbbyHENduIRvxkiwGTDTGz4hnDmiRFkMkmiM5fhrLuOtlRQmkHPMu3g4mXTRpXwc0dIB6oA+XqD
JYi92M0/r8QRBn7SI3ENUHw585YRPkGDydGSVys4vWFLybFEiW+co+f5d6+HoJtTWb4/4WJkFIqB
HC7g1zoQy8TWrJIc/R+Gu68P7OrdMszOWxpR8f28dVCr/Zuhp44kaD1vlyMOm48OfuusrsNmN0GR
fRGHaqBkVv8UrhWzdHQjUWCYTJNae0R7Abydwj31KRh58s8trPNfgD4+LMnCA8UGlGr4yPXm6XVV
+aNcgNRzzmchUDQOSwaUUw4hG9bl/Eb8Ekt5reyOQ0QNLy/EJs1Z3ZRQuZI0HLXHhG2OFfi991fh
05SUM7aMq4dAvVudirrwgRRnmwNlyck5L4xs+LzgxZi0wEpodsSsioEKW1dVMi6f2tKKgJb7LzeL
3rQOkBB1gKj35WDX6PI+3jU7YrHNe4dBJckZFEmSxI6eVGo2Rz5I6ahxkMwrOHURYbC/6s5Z5kOI
aUejd185NktMIhdbr3fCvgc1J0YGeSQzQ4holmqhY+OyYbnefzCplIt1aivUz+1ickihcUle3S3/
0GZFPzvZUrcXhMkYTPqN+ozz31LH+ISEFjD5FNfOARBcTcNeMqEjmdzrBmYs5ZvpnUN2MMSfQa0O
BdSZ+NVu+AQ7nL/qoWc5giKezC2rCMVkgCavoNnxhJtt/AujlSkrz4EGsLMyVd69GTWJisiy3HH/
J0eSfZLBI1rrjbmtzsI9w2iUruap2xb+KgcC5KupJ/UsWrDK7oWpKgygfJZVw+l6fGx2b7vCsBdd
Ipt72d9UI3ZPgIy1Z5jF8Zp3tDCIY+EUgN4/8TI14G0+p5LGRsnhwUrYEI3LmjgxSsfHEso3z7U6
phEtlxsniC2v+1DtX3YBgST8dupopRUHqnprlsrkIXLMQovViTzHhq5j0z0gyITT6ATjtB4UOyUP
BEJbi2ralcrk3cPB1adTyvBCyx3y+S94pRszqEy789Z6DIvAkRdvu2fxf37EVE1MlspRddVXcFde
2PbkVouhKYrJMrE5hX4gOEja5Q8W+nkNRv4stQtTIkfHrS0WVO2qYZpMZlwAaE7GpIBAAgQGKor7
QdZpsiHnGFkwpjwhF4wwTuy3H4ztRqkYf0krTkt4ElrhkF/D0C/H1beYzeck3YV3fQUZ+OzdJGZl
P0Cm+Gstv7G0mwIQh93WATmDIrwRe/d6KrcxY2xjPdA2TCiQbOzuxCFyr56qZP65x6pOxbnJCN7a
J3JHH+dH2Ec7KqMwgL+iLuw4yoMTHv0oCJ0mG7AlojfMdWHupqPhKiSd7sIUHuZpgYPU84NdlnTX
28w67zgHtAri1G5SsGF0eWyo8/UOVyMi2j3VB80MRJJcWcYNkcMQSBar5vdgO6i180i76TTKnWxK
xrNyZU/ftlLHALu/NSq69FsI07z57xqnsSLb/FGTX7YfANmnVRKb7hTao/CA0qzHTZHTJBo3WloX
ssURx78MBK3+usyRHrs4jmKVdWavxoHiPIFZVxua9HLMmOUJc1x69jpmNFsuSd7biaX4aZbs+gV/
4huybtfvKW2iWnbwOFD5AzGJBHnViGg2zV2vDYO3N4KuEYjl3YIc5J77AP3FhvXkbj7CdPJeWpad
YZIa3gm0RHEe6jOHAXAIbZFBUCZXHm56/Vc9T6Hbc6XEBx71k8KwewzChbeSS09fXwX3WNtJl0ts
HvMr3CAIztfebBQuo8l61lOQ1xhFtjmDuFdIDYy8bZFbj1R9Y5w9DRd5jSNk/1gAf0c9Xel07rrC
i4h+3paQG3v2tdHu1EKvkfNpOqerbY3VqIfDY06dTt9AhlifHT3jCVe7CaAf3ZGdQogDdVGmJOEs
M8L/WfyiMfJu5NiuVECjvemcT0DOeWuiIj2MKr3D2Afoo3D2Defp/NPRxVeb+XYO3VCjfTO7WdW2
Jx2G7IAwMZmskS8D//vq082bmemj3tt5NnlTBgki9tQ2Nz2sVy4wQX3ztLJEAtaVW2QH0ZTstfHa
i5c6GZrWtQXplNxtDhGMbGx1XkZwcizfQSsReWmtAArSdVMExYYLaMhcR5SsMfMrgBWzCNriPuhJ
ZhFZDhUOeJCDLluOBJchs/p//wzIuIk+AJ+NegGegnjUslC/2nbOpDGlXS8er95hp2kOTcm5u/Uq
gBtzGiUpA7+BtRoE5QBxI2R9QgWZCXHNMRZHp8zRoNzc5FXEpxrLR/1XM9iG4FehFYRVuu0a49Nu
85mDfUUM5UOMqBZ0wG3owLTp/3aFEybgc9+8GOrRRVc5OxZVtD3rX+QBMwHwWBKNPrxoJpD6mexJ
FpECD3BLJSMAbYqGW8EeEJEfgQu+rWcn5IjlCE1bRiB1LEY2zMz4T2yd893ztH9nSiFgjUiLigmJ
QWo/xqOSKZyKgykIRQOKmi8g7Y5JJ+P5UVaiiQDc/bgVuC87h1P0IHMJz+1oh47oj268yD6/pv9A
HZ+SfDeYKtVEGYfoVciO4W4cIlttT9MzEMQRuMNRdqjF668vhY4I8qCOLDgM6oNDswQ94yJXz78W
Lt3FOWnBmpjO5mqvC4NaF3evkLwetC59geCYt94l5aGdpMMWShlixADLBz7vPWo5cEOK/yy4iG9+
MWeY5fxIVZpCG44Qx6NneaYVs+tAybdTpmCKEh92IM0Z9vXT0NQOAOeQ8zrS0GmpTgIJIkKHdjDX
gwF946ecHrF6oep3Hq/KdyTou8sE5M0OKa9jhm5NMY6CsMPCA3jgKd7A29+NF/yepBpSjqoG9P81
VKipbvC5KZ22gF6uKNMBFG4u2ic+Am51MF1VxTCUul/I0qDXNNkCno0A0LA+VsHMcSgwkJcSqRpM
Jp61xabgyg0xhSD0IH8T9hyH9cZ8t+C9OfeKDJKJQN8UDHo25VBgtzPuv0W67T9X1hqiUWg+Jmmb
kPNpl5TLamlgM26Xz43LG5qOCNagglaIWGJW/g5mQHE5SzITIIBRyMLMl8hA4V7AGd6niaHvmTeu
eCUNd8wcLbwFfboshRJbXrRTcJKjqC1aUVPdGLNQCFvIhfMDLO8U4otAipTKBeFal/C27qnHikNZ
+3p0kTQdq/sU+5PUMIvkyKeM+2DsSoWqhKDDW7srYSbdGNTYnEsAUgBK1A0jOUT2LfQ4SHSLT1aq
p+8vSsQso6uQIPKiAGQoaghDqEfnxSV+QXhb8GC6M2LzBAWC1adsGMj0R7PHbidm4okfIgPVj8J0
Mwj9xnNrDHOpMWPA1mr8gYLswqJWI3i5k86u94e8rLDuHR6NkCM72bt/CC05sXd2f31xSObCLuiF
7GKHr/WcXUEXcg==
`protect end_protected

