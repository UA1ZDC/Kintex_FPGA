

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
GWT/RJdN/UcIKTAhVxs3scTnM63xEPkso8NeqXOmx+sudHjUMJ/qSt5GFjdXAqexLlRND8lEfssX
Q8fYY8TuyA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
J+phMqmkYiPgvjvEjlpcdWdxzP+34SmYIPyc3dLXEqt+h9EhMcqfQg7r/svpEBV24DU6CyKyCXke
3gZaY85pXANGRT/lW2K8drptf9l9vYajWMSy/HjvETFYNanQN5XDicKd40/UNr4NV+8K3+zJSD2+
6HJJVC0iWa6RgWieT3M=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ZrkwjC6jJHChQhf/EDIYzNRopX0ckXH4NL9s7GZmKhZ5Xuu3xV3LqvLjlAq2T+/3AXtko4HEVfJk
jD8rEKHAwLnqMbikHpL2pup+LY4/a45y7duxNC07dpJvYX19IW6mqYLKEJTs330XVwBLE1KOyaGV
xhWwwqThGo1V39JpBwMcpzmL4YnxHaTlERiq7vaoQpYAMkwdoBVpG9MMAn3CbeZJI8pLk/zNkztm
rMeS9pshqNVtzdUse3pl3EDxWMB2hg/4/G9fk9okekAXBV0rv5NMqf0xPrBsTvRJGO21aW42nO++
dC8am+sI7nAhoG4w6z/WxE1BGkRuZGX4CGhIDg==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
iexpjlh7M7dlTcv5seskQPlqyHreGwsr94b5YKwilWQsfXW7U1V2aK3O1/+pXS09S+pTH0rKoHNi
ofASVdK1RB4/i9AYD0Ihai7zYaqt6eRX7azypmOnO0M/ZZIrM+63BHWcDodlNlh86PWfwaKQSqJW
hLVuOmY14GXZev020lRZWg+2UhI/Cl3c8nww44erkAvCrpxmrhaZg0s2YPKI/KBqZbZHwn0ufJSY
5EPF28uCCS1urKeejeaSBUmimEDyf29zU/xFd0fvevSdWXaFhwjT2mOL7DranIxEzj0yQrN0jiKy
Towa0uazE4xB+gMrElDuwpcw6ZUMyEBsaW08mA==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
DVPBxTgKjw13z3lZMl+QMKXV/uHfXNCgMoWbgQb15TKXtTCmkLiaCYkk+UNjnupib1FZuwkbZs4q
pFuDW3Z3x3poQoD+4+Z7IIYAmkcV2VNFgSXWGO5qpHWhRfkulPfZcRStTLiN9EUcwXJUsLi1Rwk0
oFaVSUr3p4Mr6zjC18beDCFomH1w+aZiTDmIDtnqdWVtxtresAhXiT6k51hdPESOpe/yPCGrgQj7
cckAkNk0Y7ums+FtMhs5xsfKLV6GQGr8vql+qoCmnMNbYofWKIq3pY2FrW6f7ZGbFhW+vgaVatOo
wR1vGhSucCD4x9efRbKZpd3HOhDW/vOAo1pd2Q==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
uIb1xi/b1sGS9N5+ge4ctTMaXcuHePw5wBb1FVa9aecf3hzk8F8+/rWvK4DX9IjVKEx0PLXI6xjb
IH/rGtJXdtbDJdBaXxCtQZnZ3bb8a74BAJHYm3BEextG398AX1ZCOiiun/unyz5EkREGrSg9f1qp
tvP1wCaUgYbP8iAi+ak=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qK9lK7oKxV9h/658uwPcMAAwYeLmnKNpsdduH0hJUA8HIiT0JfF3YHf9Z/+4sugCSI1ARr9LlbO/
o+J2NPNqOXlyDgJW0FGjeX+G4wdX5LlxdfSIcRGs2vzyXQiAWVbMq15jqJGV+qheK6QIsLI/qwOR
naZ46kfkwSE8kQXhF7WZE2kD7kLSTF5QPnmYFPP1wrSHpjD9hfcjmg2768Oxg74FqPuAHl6cX4Bj
Enf4+hzQMQ+IcGssYzesFwyeHIqJFbufwMH9hDnmz2bOveVtLUI33QRmIvvIjsEuvmQwCu/AC3gG
UyfxcM7HSiPQe9MbxhcS0KjoubQbTx7z04URRQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 504864)
`protect data_block
0CAib4nJVSnsovYW7B2gFJY8c77VzbfB381jlAzgqSXnk5E/S4U9CDr7kUeIPTtx7xwyJZ6MXgJb
PfXuXV4AVP+TsEgHB5/YOJUhPrHAiIo4t+ANddCgElrCGM0klWHhNzHFOz0yMXlAhteZVvxtSQxP
B/UeYhAlbhB+wPMYoiktgTUQgUcxg8QRgR8Skiu9q6Yl6d1syTmePYwZNQ6tVFH5XOGlFcSIkDJ8
kFtyfmkpaqX5mkdm79oTqEQWCyVIpaHA3XsOPXQDL70fLsJnfGzuLCugUiv79ilIrjmgGFJkI55R
mHwkSyMqK6mzIwBoCtIARV/RGXhR8X+N0vAlplNf1qozLUtfmZ0giGQUSfnX/0xM89PNtIwny6u3
cNK6LbQGogq4Akst9zcH+2Tt4AR+0M+o1bUCzbxTEmF+O7wFblHswv9JLqDCQV4vYNROFzugiaAu
RWFNoNm067sE9gkY4+VNsoFH1y7xEAK2C/Y9cRECYGf5XpvgZa01AAHcVN4LE1ctFCzW9bjHrsg3
xp7goJmY4x4zrku0q0LfpiXrAztmTyebwDxaBfiynWgfk57DqgTkUhipjoqjC+OXn8JEzEdaST1K
NQxrEr6LuJaOk7duW3z9fAMDqedQRUWdFAmCeCotaTlrawWHwUsweXXp+KLFE6+f6LFYQ06uSZ/S
u48urFMLS80+jV2bRhyRrVeVAc05MVTHGkrO4s0hZgGJoMMaQZC/gymIgtcySYRps33sOWlSHWIV
awNas9u91+Zvm4TgINanjF/J2CMj5lusjEBkMx+b2TGbJfjzki+xOdoyq+pTQqh2UTm/i6/2+oMq
f2DWjV0t48WXEIHFttRGJq+UFk13YOvOouPlQuzgmi/ana7bdSp6jSJ3bQ//wchtSwaL3XGspUK0
J52IINnNckqEPpHyQI3O2Lwiu+mwTi9AP28lHp879egTXwEiiiwGtHgSfopqnZa3lZhHBgDVCJR1
YYEugIxUCW7u8OdojjkskjZgySEFMfLX8FbDz3uh8f/IIN4JNSd5BplB2m0mKiPQZNf5nWGtZuzL
A3dOCbe4q0bDoK9iBeBcUllu1CzhQ3UxrpCw2ocONBiT3fwdapfuYAM9wYPhVg+DvrTHiY8lKKQK
lvoX+5XgMn2AamRvSmc8BHu1hz7nlKqRSVOhLrNUx9tzfbj0OX/XTZf/rwK8yA3C5YCZTMWltQ3Q
N7u3EV4v4PA64l3phHyrBMuY0sZnm8pEpC3DBmfz4VCU3zrnQXJYOL1dKbvwR7VzxZfNkpORlNks
Eed/G3An61azL3iywZiNwEIJwIo3HYiPKgRMtKwRE6y9P+qRd+Xe7o2G+f1dSQ2ueOJOTIbjxzr4
RDVnYwTitkWLbrveMxCJFP21gdLl35sSs/YKEqiIGrZ9R9do1LKqtHpvCOmnVblSznRAFv2soKXN
awhnis5x0VcOGKpsDJsoCZxZ5uS73mhblK96rXW0n5NZVAGv6i86qQBi4ZSbZjkxlLPCvwJVHyeY
fU01eUNM6ywOuCkjOHu/6DFfLYafV8VT6WdWtb84DgXONlnpOiLwFNLWAoO47Xack2GbIxnRl9kA
f8fKY7TBayKiFba/C90FKgrrtCij+UV13gztrcwovR1DBYDgXjxlJOxSGUbhQPE4D5VuvMX8dLNi
ii1dJvgKaLFDb3nvGYbdHjLMNzQZg0qSaU7Pk6rO6G14p8WvyBfbsF1mgQgytz+j/GVkNyD46EYy
Ymj05yEbkMwuwp8KeBBkjnwElioJqkfh7U3mMWWjOeFS1uL6OuIzx5+U3iSxoaU1O2wJoxYIqlBK
1uZB9fZ7uWhqyQ5J5gwnP9RLkXt5UF8+xBschYqPmXn61fgkL73IFSvC4UIXOuoMXTkfGQfSy9Wr
H5LFiY7iKZY7ytq36BI2OmAI4QDVMYDJB1IO3A2agCyuXW0+IDZQFgsjsODagwWJpt/gat3nkAlO
Q0w23nQxExA+EiGQZk2pfW16mQCBP36c/FHdUCeZ92b+sDueORYrPVp6xVLPKAVNpKCTLy/TXWB4
dmpJw9pZ/VPleS6RmHWS1bHYhaNsK12XM606sTVWNF4QkwRUu0DdLlHuNN/P+dTWVXl/+G5l0mhP
Hv/4OI88bpWiSxVqfaMOF6q7BWWMaFa96fT9/lvaYc6hbQu9Aez13LYt6OljYK5SnOSo+dx3Xx1j
/V5m+ekWOL9hFr5rZF2Crka2QeoHL8hlzQSk0oHAb79aRhz912+RcI8tCRxU0k5NKpmaqxLhS+Yn
mXIHBw4l2uKOq5m0PcaoWg9xtlw3xCvE2pIiM0RpTRDWajXnef6s6dfKeGee90jqu87pKOr8Nk/Q
8WMkz3RlIf8DSOYviX4BFwe5YpzcueMu9getVjNEvd5AOmpdVoHQjlA3EsmoABqTI1Cz+EvjJcKm
PqIoqNFKdr8d97g0sViNNLo8OTmCH9d7KPFFrt0GmevvNYyc38igqxHPfunn+1jZZRrGteCBA9sc
3wYHuQFHDmkFnQU9d8qtUoQ5T81fkwXMweJyJouUGekTvpjz8iA7U9+qEB1qF2zNPS5O4T4yjjHU
FOU1xvLgkunl+CR483LLUMFp7RMJrrXXrFLF0Wd+Zh0tO3Mn13FJTLG/chGeJdv8/lSXnOaFzyP8
52/rcKzl1irY9rYB860Q8yW6gursP98feNBFueDMamWxqeel4b1QVh4nqT1+S7G5j8xlizllDQZC
4VW0+bTfwga3poczX0DjPSH6gy+Jmgp4wSK0uodb1DXBKMQ/H5D8CfE4g2uiA2mZ9rdov8vy9YfC
15AlIXNi9oGoH6t3291LuA4rfBDq9ssht6uEq23gEgp6DVwCeqPuZ4c+dJERzMRMgrUWpkLiryJx
p0ZZmHb7B1tHuT/lSQWmIgdnV+KsMs8EiCdVH1PWfN5KN6c9ISwDRWgpOEycHqGk5X5jc9EhVO2F
XpVamfaIw89/OIoYxg8f7Icp2vqwaC6pisP4WPVjn7UOqdQG8EwPcmZsqUbquNkKmFs+oNUQS6VV
sNrMKXlWA3Fc2mYYV/UjPzsQ7F6ldMSDCwbVme7ZtXRLXHYFTWF4mafg8VbCXB1qlGglzeO1tsBE
XIR5Apmh4CjtTJ2s86ucX+yIFMH9XnSiWcZQ2aWiNQPm/Ald44y+JO//Wj05QYoK/yeGU0Vys1ih
2ESQAFCDZPq/qp0qa472KqPtF/z4A/XT038ST4XyT2/Lkoj/Bnlz6RjbiasO+RnxarkAuSDFSpNM
AID50J+3ITs6bcwUCNsONstOYlk9Iq/wyKzNlhiJ5xsTCVrxg/1Zr8A7WnWPbhhIGWzgZrKJlGGH
KRbHmjEa5h8xK58+YMlyC+ErYUcDqPRp9sUJ6sdnuK/FqO+wasKMTzCsKjwSde1sjAtIue1H5uKO
odZIZsGQR3UYjdw1t0iXcJ12iNh4+g47IXpB9RDzYtdvez8yPqOaADiIY+7PLGn4xneVhr9wYhsN
nskNRCbDxW0d2SDrSFnv2358lfS+taJoOLeZvx0G811i+PywxWbsEFpP3eBjo3iWLmNhF8u02Uoa
HYXybtESZTWWlrdDKq2PWuzQqEt5CsI9xyCX+eT69JuLCD+Nvl+ODuPUHVy936/UFIwaJpcSr660
G5IupRGqH/x4o+W9bTsYs6Z0tanNs3jF189pue8D1UWOJevdTLMHWrpNFC+XjnNKGhtXim7EnlYn
64xuSy48vGcZsiOy0xljUFofg486Go2u9rjN5j6S6gBs77erjyDknPV79NV/v6dE9pTmXroETvfp
T9kwRSK1s3rbDHHPmfIfjWeLecn1rShVRdw7qnXOiZXh0qljraqQyZmsSZVAVQIHgF101LtgcM1+
/8WVMnQtX6isJlE6WzZ3TU5FxfF1qOEsf+sb/NPYYaZC2HiVqoM90zM/BIf6PXT1Z2m0NqUsbr49
xYq/YCh198ZfGwtD/suJjO+xx5E+qa0dM1mYjF0d+QIfnOXXiZ3HmENtrzUgWla6Xo3oYO7ycg+Y
Yy6570AS5o4BccA844pTp3AizVOf0rGqcL9KWZ11yNQ67KFX+V98d2cTzkQdm7jFF0bFlUTqEWM3
sPeXbsvOWE2EwESvgbpZR8uJtJ0e8QVLcAp56VQ34ZmN5s6uykY9ViZDhyDD3doS3lHr+vcIC/na
FNTzSSlbIgQlMsP2dj2nT+Op8mDEa5oAj4BdEVd2Wom+W7/NWKNr5mdYZPI9c+ZU93nUm3VPe4c5
9BzrcyTV00I6aTjGhVb+P1884FY1zUQezR/RcAFyPvsoqZszE26xtLVpaSYRZpXtRgEwkZ503sRf
m+//WwB82M0snhkhNK2iXh5NUr07lcJiWUMPW0gjEIjCzMMlltNCRDu6rIPWQbAgO49uYVkJtWOv
+qzFLbEx41/W/sdb5o+y5dkkHniJDML1/VuUB7Z3KyReN2idIVG9TGZQmWXM/nGV0xHlLPI+8Xfd
CTdBVFAvcSLNtnWLIxu5WbiH8SrGa0KsZnxgrtvn6ide/jq3DM8Yct5WWOSMT3NMgBefEfeABdBU
oRivaT/9eMdHwYSMs0v7u+WP25FrYjVU7FEsFuKfQ0Qu7V7+DmMioGg3Ut7AAGhftCXS/XirmPdO
smauL86nrHtgeAmrd1HASSGZ33wuPJbEYfWojSyesTbSysk+KyqGIIB23f6ZIeGjHMlBaswM+E1o
7F0YG4C3efO2BzXHLKbxHc2sztEt9Yevj1U12Ee+AphegmrGoN+ZN6hfgwOaysMxD/X7uPvoGeBX
RMTCBcG4LPCWugy3/mxDwu+5m3mSSAKfCYvfX+e2jKK1AHrw9h5BZLhwB2q97pjG7wWTVu914kW+
tnHjXn8Hzc/fVnqnccHhA/2w8huzy1seEBJt/nws91ZLq346I/QK3UIUz8nacjjfVci7FduxQBGA
JdjHuWgP/00bRGwLCLBlD93xiTxOsC77FiWT+JWerTqZ4HRHGCYUT+ckTUuRp0L05V8yh0FDqDw8
phG7UyVzgbTvnCzikRKe9Quals6SItMBhutRqPW+jiHXOjzzU7N9qqeClKrC3XJ0YG0vgnSgo81G
zV3dVZ2qYvDENm5n/dT/QrZFXOcs1jUqZIkdmlp1eZEPJ3yclHikzkMkeDckZCulnmbLiAF+DdlE
NtGT3aw2h+mBAYQ+6E5Wwm6VPYl97uvypfLRGx5H4uZR+uhm5S4CXDXbQvKUSvIyA0h1eECGVvhB
1QFXyyVDfbl2k294pE1VueSpWR2l010akCDd1Y2FeJGi5KzoYS9wbaTuusncV/DjUcPN9//KJYVy
HvtyVQKUu2Vo7cVLIEjKTe0JbevI5dtXhxP4D3MqanV2dR5ayVHTs2vX/WLZphH593jhCe+N8dm1
Pkf+e5Ip94goV8tcnaEFBiJ90/cdwLnToCmKKqwB8oLX9JxR7IG+ajI4CbZtPxrL7YUTPEj38nAe
cysXZSULQeW55Axn12RiSNUv2YOvwoEwLPziXU5cMAFo1IQh5vHCB4o2eoiDH4Y0z2C8x0OTiiR9
jdaVDMGefPQrCb+4YsQ+2UT1ppqRJk6TcQrEuvX/BxyfsZjtdBIXzIQIkEE8MuzpyDGhht+2kXgu
j/0bSBou05mW7kZdDb05bH2p2txv4szXy+8bgZaLr47ku8hKDuemPXZN6ebkbJjIY3gbSRXIWA/e
Fw3SO9GWq2wpMlhT+jF5Ls9C24efTRoP/lH4dhxa6Yjo8dbpED2IfR9h/i0FPMaqTf+AJI5wvOGq
SIxm+AfUj0SE4hzhWMFn9V5jgC/GGzmv6E9+WxcvDNEKGpN2D75D69niLGQJAANwBnZEJP0oC66y
MfTfvCmTY2cl/CETcXO6ruayF0ELYG/80ZIzg3ZQFRXxvSZJ4HH0yWbxFwWP3Z7DxH4rLuncqZQ1
dcAhR78NErm/SDxczW/XbUzRxeg4h0KHQkCzubwanEoR9hA8Z7+Bjj1lfg59PxSKi/hTM617RFS9
bmLGriDxgjJ+ahDQATZc2Q87A9NEaIeAPnLbagdEKK78aHQxsCv7icIP1Mg+JKU6NG5tRNsw36qk
jibXGzEchQIWANCWAbYuz0hOsoBnR3qiVZPhrnSaeGRQuvPslxvq1H92Bls0WJteboOBqx6uXy0j
sghYsbnhJcTv7fTVNSNlmTqOcs7GFkl0WuXbHsVrXw33yeawwsd2uJU+6C7tSxhCiA4Q0amD0GIM
3dafEl0wev6Yzzl/ai6TYxTJQRucQGuMpsTxZp19INrYztZNAOordvguLr+xNMeZK8MobVFOQ7fd
k6xQrzy30MBkqg4Te3rNBpgUOMJFb8yZc2gnI8Rh398DA0W74zcGoNvgw2HhLd4gCAZdY8Hv8upS
HaI094RefzbGsukTSH3ULmG5UvWAeC2+d7AL/hZHeiFj3cAtm3Ggwr1ADUAXRZHJO9JkNm+ZCI/C
LfvRIhgMl6U3o3rV3dFzCEgaMsLXAHLgCIxdv1xqMNnukL1CFoMaPtdmtDvcYnCWWGaAtidObWe9
BAdHvor8quF+J+eZd9mKmF0D0WONop6eLxvzXmg3iTv6ZnZvvm6D2++zqWb5vB6yEyvxBwXe5KIm
6rME/XctSW/p8UV5oQBFOaB8E8I6cU0J91TN1viHr8v3XbwmqbQKUrMMJU4CHjAxWygKziBqqvc6
EyiuY1XB56SJ+SXAdviR8VX+Z1wL6bmD6BCnI8VREk4gw80xYwFZw8bYZqKNr1ayJbMnfZmyq6Ip
/uyyAQe9j6w5C80RwhYCsJl+OxuyBW1p9qSMW7TROpeToKh6riGY4q0u0IREOAla6YYWNVkGDi/8
E9K42A3gI0KcdxivJ35J8Qg+H5ZchTDepO4aIZWW0nw0y8egCgpzvp2ujjDCv1SlP2OfnV2heKUz
RoO5SYJqBL7Zl4Mq6N0kLCVVN/XflEG7yamLcqcw4bo9qCdWAQg8obIH/yBiCkDEEufgVMd0F+ky
4RyQwc6NoRpAMVkJCKkF7vdXihnE5RIojUQvEz1VMpSWoP3v/sqciOfJUTprxx5mF4OG1cgtCYbC
mqeZO1BpHxNQ2IVLj/vjoWuc4ECMTU5vswCe68kNt4bEA8UXSLH/XMDpgnl/rzZWbtiae4CVFbNW
wy/DnbuaSESFa4Zn9sCUazyST4DjC9BTAb2LH6R8/TWQawsubRB0ObIiNDz4YSJ+2XVI7K3pCqk3
/tmRTIgTfSRtzCT5srxx3zqQP0HapzLGWJZ6jBEIaN4BdND7C6gv/0HkiuEN2GNt9ihmsX4ecAgg
fqeSjG/mJ6n37by0yepgGkSOsjm+QnL3fORGC0ePj/YwYgYUL7/sUUFVqQHPtnrXEgAP7I35QcMh
yGh/xDheRzvM9joP6FAZDlbigJ6KmqIvvW+GunW2G1+9HltQigJJrswiHSQuniFPoypgxAc6s9AZ
Enf2L/o7W6gRBdcCfc4vknw+HcCI2X9lMe6btPdvxjS213KWg0RQeI2plXP4zFnNMltI8zET7KaW
wItcvznNyr4XHZFg0DtnFPHciMHeTDVMeiMZ5OnHKm9dHI+4xIEDXh0AGl46mvPMcUkRE15PiJJH
9oL3bq7Vn3NLL1Zai7qEinC8vvjagANzuJfDzCKaNg07M1ebQZVgBknqszRqFSJ19r37rKqniL+a
XUK4qDfNdx13VBdzDMRGk1P2IYQ2ihnpYiy9VTqX9NrbzTRz9EOgR3rRM7pvOHZV7Xgd5acG1cBZ
EYc9dSmQWg1mlF38agibmTzoMHTfyr4mkWeQjQIi5nzvT+A9Ih+KBKzIZnbuYweDIE3J9/egSkFL
2dOV2F7jqBDSimOHPW2Ncm8Ph2z/F7ml3ghQ6a3eA/ugVOQSnxBMaILwh3S1usmCXgrtxDmf3KZc
Z2farpWmzsoVEniQnzqe9R4WPoBZSPRrbn2YwruchW8wLEKYMrWiLWefUNQOuZyuvCZPd33NIqeS
+hfRmJ7zbZuwSI1beAWl9kPnrgEz4EMbGZlO4wBG6srv67UkVOS0A6M3XS0iaqgo0RJ8jiD38CPn
NuDA/dwMMSsB8N7LqbGEp9Xs7zD68L0e/ffskwgTPf3y/fw3rO+2KXkHgFoOFoOb7qJcxANgfA95
xVu5saIU3fTWV7bqRJNIVOBUxRzDFxGDrMXRbcCNCc/ngl/Qhl1fk4w1BFoyV9Oom9ilSxTprQDG
v91/wWUCG4ukxOgmtYDu3eKnMgJG2L+8NYeFOPMHUNzNXKXWY55bE7d9XIWe3yf0jXleuq1ETMCL
q/jehYWaEi3Va6GNbNhSsgBHtwoe9qRMN00MC8efuuJN2ziDJg8z6Umey8xVSLae04AzHBeXekbG
QDxLql7HWFZFSwGP06grGmaf3pfUNGszfWgz1OtPwSo81pous9SO96vL1VDL652EHhfc+E2UaIVS
lCxG3tg48cHgno8/bh2fMp3Os5nqCNV/IBTlM8yhx/kAuP7tBHelKwOSQItb6VAipQ71obbawheU
CReItm/WD4FXxI+2dJYZWnopmSFjzjugXaYEFuct7loK3nxSHw7NLWSTL1Jj37ufJ6w4OH11p+CB
QnAl/ySVsDIEcHxaHYGX3vRtqyIHNlfo3bMaslQlTFt06nZjj/IRi+ywbzXJ9TkijAt8YBmQ0rg8
oMvHXBMzqGVXdaCYnhblskk38XJkXO2gPaB0BsdXixMbfudDPMS/FoNyDYj/7CUZ3qeLzkduibLb
CTRs/CqN8J0ws+CQjyURZdMQqCbfQdHOnPtCnc9rDFMcbe+elSvcaJKAC7vuO+bW/spqsCTEhNLx
lOj8MFI0BdZdaTfyu9jLTX3di5JVrzEMqLEfQIL6S3rH804U5Bh2dkcpGols09qCJynW53tNaWl+
LJJueGCk7dtBRoQ3Y0kWwK6da6Iq5+c6AKWW/O3cFnfaxRZmts2Z1q9hHpEmKtVGVq1bu+o+AGrE
FhXBoZI0H9CVJMgwrbJHbZeVW1Ymoxu5ZeENbB1LxO35asEpGcx98U8A8YOJSkmqwkG5upWc4LZp
Cbcl+fFopedcdquNNIvtYNck8fIL23yYSTAwUd2fMxYYaIP1+f9QcPzbMImSh4Ze2E+6RNCBzRrD
QOKGZzSzgUr0NqBFXixmniS5sMauEYaiPviT1P/tWx3KCQCpY/lAiCTH2XM0Le0hHkoU6/CIlS1V
b1zS3riguI552NEeSbrwFQXyS1GFXOEVA76Z1xS74Fa++Mz/YhBNY8tEszIPFpUWwvW3ZgfmqCVy
lYJLDrCa0lX9EIu4XVq3e06Pw71E0cLRwC1d5pQ3f3qG6fMiO+cZhdSLMy4zIYZTWZ+jJ5QFYgsm
3a/QvGRuWn0ewE4tjwJ63vWm2kYaKP1NW11w5Vi7WQbS0UvFKvTwHX+7fMl0UcdxOtIKC+rj2n73
EbAA3SHGaCOu5JKc89CgI6MIvW8AT5YUGqvpsuoNJ6W1wTGML9uMXBTROea8b+BsSUiQUVboS1RX
YX/w3XSpNsMz9pFjeQEuNZhvHnS7+ct7NgKemg0IFPW/upbVM4DNI7cX/duqBapkg7ZGCsu0yBgC
r84lCMJU6jERyj5f4ILF1gCbsrHso8Cw1UIs2UAqkhNgBBMUEh+HtahupvvaZHqArH3RFXlsR5kw
GcfEjMNxBuUAFD27KCLAesIo5xb3eHQVjCFaeMCqVd1GEzHqkCiJHKbppQuo8ptVQ4yXCAN7HSp2
LUCof4dpNDki8j4/1l4g91J6ThkpA882kSPkBy+tcDK3U24jLBg1blUuQJRGIMdcMUupcdc694cl
UDhgRi52KXqceGt/G+Lo7Lc4J7Yw46luFR14wKxIvp/5qs4BtHmMtjAQe9alcy7b+Rrfnc2sqraJ
oBHOqHnCBcRC/13F7gtwZ3gu1PVb7/XPVCTpzkhVSt8NBtcaqww5rrNu1ACZqOCY0FyqmkQ/Xhaz
d7ticJ7gp7zgqpRLnUtgkpMbep5vv1/PphHnot4OOh7zgwEO2VtGMtJteBzVtgL/36By7YHtLZrP
pdrrcNgcGva6xZMiVpy5xzfkG2DTVHzRIl5N6fFTOp8Uij+BvvjmZkBBZgu3B3knYv2yAfziNOHM
fWdMIgGaK/kXSbUHQdiute8cNqPbOGOzWfcDMpiI5LOIhqKg6HHlWNYJ1SBLsABK6sbub6w5Ojvk
34d3IISNdGd+dp1thYYA03NhTX+FrMlBT19M3sbw/ALOaixCA0sIW2PTKEJ9n1f6097a67/l0xBt
HW4CanVvs66hysLsQ6mYa9B52ulTyaZYM6+c0kOJ+isljUh5iOXEQcDD4ERixjp2tsaVwapugtOV
X3xXVZlmD1oEuAQp8jQk6tkKQtOAW4DyyL20sY7NodDfZ0S/PnYcr4jpF2XuCY3xKnHtyGVp+PKj
rsjQCZA8glxYRHERPiGvg2R3k5QBPdy2/zQSRAuZfFzyr+hTOu6s1o/GnmOfOMj5XW0mIE3JmG7d
7cOTPmbe/o/B1smcs6gKXoXHRcujUieCrtzQFBdZJh+ZedgkCr93e+F9tHg7mLIbFdZWvoFKhOZY
y2BSgfJ14FUFDuVm0xr1+ZQXpVM8M3FOBU+EN2U1CKw3t0lPwddD9Q6o7ayKmvjEIe7IGleE7Air
/LgrLHHug/HPsIiqEVojzdj6y+FdNzLkmIMBPmlXkAvxxieKBbgmkL3uD7aLswVrl5tLqv4RA2HI
ZBamyJgx63PPQ4kqvV/J04DY0JV3g5cygOdwUGSCCn4KONXeSWPF0X61ewWs2ZCcISluDybmTJhk
cpvVWzw9J+Z2Koz4oe2tj8CGs8MlQWBgDlz0xl+K4kzDv6xzW28ZjIx2M+Ih4LLokiZfewOwhjcB
1EZwSFiIeB17XgixopvSyI/EYxbakrECNcS4Oj/SR11+8esVpq/E5lblv2pMOWSbct4gNjCpayIR
l8aBbtMP0wjwDyzDn08+NgQ9yZsWTxflTQrg0lyCYY+669gLq7gjSn3ECkDKJezYh8xtTZhuHpcP
EvIfDA9kXSKrAkkc5yaD6rJuawneRLpobaTEryE6aGoMrL5FhEo+U19ZqRhdwheK42rMOlvvbJmg
3sKxHck0eOWIvQwc9Wh1RWZ8S2VN2xDiNnGq6R4BtRDvMaw0eTC8N7sx4bIz6Ur1EcNXF4kjIKTq
rvdobukU09JLvrieMWCTQ+0RAq5YCT/RIr9vpif69bUuvUbA9VD4bCBtsqTmtZGWyotLZg7dTEAy
Y0kD4MrZ7tVkka4ufiWSrMhKDOvVc6XMLpqht7xaQOgvcwiyuga4HCxITxVju4HmmknzeylzsKg8
MGB/ayBqDXBk+aCbKsW5OlNjFclArWia1otoB8wTJpNmQAaSy/Uaw3gheOaQWxcRDTfvSCa3avgm
xjQ9sI2/aKPQ1tgVqFYsW3rrXVCUhbsnMe5JCu6TnYkjvSiO2WH8wySxwsk9OdGlgSEtQeo9hVMB
EIq3sYxANfgzetDzAHGG281RSFOonK6Lb3ZuNnZsdwRDh6WsaGDfGE1oCp8340TdG3BJWvMKvPuP
vKOtijuolpNcMqfJCRRnvzRMstEUVB0xpHv2IO52bwbJmZcw8sgEzs7GkOv+KKufOiRh2vNLzKHZ
HRbV2oQbsFlXizVKOXb3IN+tWK5lag2fcpKgt2Tz6i9tbHeYEEs/IkFUPw8K/SJnu9oZ8mYQ6MP7
7l49FleoxcT1L3xCfNCaHRjmL05LSbj6gkVa+eOz+aMiIxb+0cio0AgJSeEGE+2hy7GZcV0bPlFM
+v7Ys5+UQcSWQMyd0ujZ/FLX/mjnFGEw76fZiidUGxce7owNOND8Ze7WJ1VdGeM1GnkFNWBqrhpn
bYyUgPCU1hKq8R088s97y57V2fyKR3V5G1dx73u7kHcAG7ORqxRW7wkaatJfwdkqcnPSTUb10uLW
VG2ocwQpr9iuTLMp+zstJHusZszmugfnyku+sCRyAklqZ21A7kpFdcxMG2NdbnW4UTpjSMXut9Ny
jSuzAYh2dgxlSytY52NqQbxY3GlDLkhtf+p6O/Re7hUlZ7x96ThyMEd55U34VXvLXRrRH8IZOLcO
uFN+3pYYqt/VfltIUyUZIMXj40b0xhq6Cr9mG/+jGULdykG4M1htEXEMctBXar7s+jWj5EcjLB6h
iDxGIFQ+ZXuKjkFF7MfPwy7zT0DvO0MRY6jp+BCG8R04MhlciC37oMJuBiaQS+EbzevkLmBtmqFs
542HAT/PeFpgRUmCeJrjU6ynjkHQcY2PiHnf4sgHG9UtdQopdYUTL/bsiyutQ8o1hN1vwvrpd/+s
I9Ek2+ob1W5HEDaC7xFFvIq2/z7JB5iIh5TWl1+2vxCeuFUDx8FDQQb1EGfpISlinKizvSqfbZ2Z
Rxhf1TJu/fwFGzzmJEJ607JbCiOIoYaPDl08IQMlfWiakI5sdfMytzFO2Oxxo1/koT+14M4yvk9t
+LrW91TQ/KH9cINc/F3FV/k6PVXHDBFwre/mxgeWUwArsjKfPUQ6YsCv5gDAuY9yOWS20R2uvN4S
8LUO4A7JyVhOZsLv3u+vqL5XBth/3xwLNMCRJU0BLS+uVz16+B4CCThl2KcPHM9NA/UwXkb3wtiH
87/KWmQ9AL6PSYcRmFrtgvb7ljWaWtEUqu/JaRMQWppgibKxdwCIgwsusCeQouGbumTq2Bq1PGHW
HGvgCohEXhDS+KIgQz9BmKG0tSqQ8NU6AsO9o8+Vuvd+Sphaoj6Z0pIV5W7Gy6VH0IhR7/Ks++T7
c2M93d4uHOFRDmsYM3A8L+XInTQg5mhhk8XvBoClOI4B0DHKx6ucEw+j/+gAwOJw8E7bX7Gi/d5n
ximaGJJ/3vf9ggPIAzV32yvc0yD5YDX8nvK6wuRmIT7VT1/ck20bLSIuQCeIX/UecnG6SHupjIAC
kb0O5rlVnlDFSXUvX5lfWFRo5P32w5G5jrT7NrlhuIaThinFld8JW9evy0P4jMdFtGkD4RtOpZZc
fWVL1HB/ZqNOQEuPXekhNImN7nbcMBj5dNFvONBKMdbrO4BE3MuWu9vvViVjTwFv9oyvI+hYq+Km
NoXn6iVzl21f4MJWQfT7nrcVkd1uswoDljifDK5uKCqUE61ZwuaJJFci5Kq6o3KHu7IblPStLFUX
VUGMdbqSB2vURuiNjVVP+Gsh3A1hmS9ofwmLXWG1eTZ41j7pRXVeJNknCDX023zKBeccBvD2vcvh
BRRzCTRXODqClAyjZhfTe641p51z2Y6U8nb6gSDM/mYeLa5TGPBFcmZmjSHG/JK5H46BFCeV+uWm
3mlMy/ROF6C4bIYXhHi6gBN6siuGBQFa5E1NNnQtxw300c2RoQtUr502e50/DDW/3g66aa4wOEtI
rnaVCb1jDe5bXfujQX5EcgU4pPYyeckinj4Ocb+oBN49Kv0s+n/mS4ds78AGs6iySvnzQXoKWNNm
7+GMLkEtt2+d4uME5Viao53xImJGX8rnD7tgnVI6+cgOkw9CdVbYEBLFuwd1ypyu/8jBcaBgBLRg
tXPQqTrGopEzqBKIfQSNTAPVji+TJTByryY1cAEUKGiUwUk8m8hSMATIk1X7O6U/FCtQy8VlCCj9
4v6inHHG1k5B1jcwmMzvMheAcwKJH/wORTSNs3YvK8jVj9s8mgFTyd1OlJVf19fFtTLGtKb03yZv
AxXuuzbCi/W+BO/ZlUbWUaa3RbuTbwEr0LfcL98ofX5DHHJwbO2GJG74D9+mLJj0M52q2hbybSbJ
8w9LpAaI0kgvoiYrYCnvvWL5iEnBIW4U5VEEBjr8PhQd+ZltJPJnpscR71uLuoGET+pD36vgpaGW
UA89HZ34aCTZbPaZ4gUu1WhH8eaWilAYV2slWhGXjd8QIfLTx4NzLUnZUULtvvlGK2aANS51+SrI
y+Tz/VN6kseT1KR9F9f3gSeE4zyYxZ90ctjA8cqIoTQ1iTZJpTJhrkahy2Rp+cXyx6UbL4JdL7yZ
BLLBKN3r3gX2EXJfvFu1A7dzE1rwGpdep9lyqvsjwIS3pkkAW/59dbpETRa5XTELUO/Z3g/gpHeb
UsJFUHO5JWbfUSTUDJqScLvgmhjwLnxO+AAFs0TVBN1NqFLL2dfdEHr95UWVTF9/mF0TwXJRjnSz
UIc3W38LuLeD+/Y1IUicjVN6zvYzQTSkT3OkNpBzVRpVIR1SFS+infuI8s5AbIwuQ3QffBtRPqUr
jTsHyq7eGcLwmXmmG8o0ONUkvvLixq+U6MGx/J5+n9BOXJmtQVS4oJU00RlezmIqdWzrmIF2y4j5
dXPlJjEM/LJsy1Kn8qvHJEwA+0UIXDtrEqjJnEdR9BSJ2OZDWuVhwn3WwTtWdbCYzrK8+Uv8vDka
hC4i272K3zvHhaZ0UDMKqic1MwGdm4JVOONMwZj9VD0E/0hJQ4l7ZEh3s860BSjVrWoPTiSwbLGU
s48cm+uGt0iogGL4OFTbcYNnAAzF1ccs1Gk7UcIqwPkCOj3wIFZTwt5ee1BRT9LsSlFDCro8GFv7
Dg1RFfjgpPIKirB3/9Wi6wwsUhryuj8B3rWg5WD0rMxi2aWeN4iQDPlBRODYEERcc0TwnNlG9znO
CH3IydAeU2LWq3bavicpmaOcVbE09Qvlevj7BTY48z3pyOuY+FFBQU7H3eG0gmSPMu20Erfw/rYY
RB8IiK/eJYP3+J4+D638kneGJemZYPUmTp8L9ESoUG2ELQ0j8Qt73PxwgX8d6TsJhkfSgWdRAlj3
5Iku/0sMyZftXVBTnp9Yxq4v25NtBWtnZkAroRdqBfTTKJoKEEkipq3+tiOsLSJwwNCT6hEzqVZY
u2HOTrooMr3Y6ROz6Z/s9Tsa1sDxrbUis6h1J8KYw/yq1poh1AJA14LrImzzMYpNqdE3mmLhjtoF
EPvF0lbZH6p0x0e6OlojFVbhtpjepD5vG5JZhGZ/H7fUbASp0wPtztkcubFimCVfTGpIYQn6nA1B
5bduSSNp4gqVoL5PgRhmZ9J+ZF2/YAJm/XynDlErNrEVFLnU6Z6sUwSt3KzhHvTmnm22dPjmfox2
h49hFWftdFh7Dzi3fEGh/SUpz66Y+kvjm6kvsfVnhNht5N5mJazaiLx1ya89EuAjlxk/LLEZZWqk
gAXDNgE8/S2wJDydLjvoduB/EZMopc/nXP/Z0lB+5bI+3l8SeK9nRiVhr912V4UF3/BblmS25Pys
A0bmmYfi3fLwZSKRAOSkFt/viu9/66wlZaUWeQbb2MbYgA9DSNiu/tSmwKMiRX4u6BuXYkP/deKg
2kw7fGVd2WdNpK4R4MI/FXHEgalB/H0sOmOOqXns/FG1107X/woqubI06kEBR1fafxC3i4wrBwLe
zb06/nyVlsw5EOahbNpy7xhwIzarpVgcxgR9fHZ5EoYOfUCDy9W9ZyHKGGp/7NJqqO33SDTqz6D3
6M7xpzuBYAsAst2oLhlu9/83m0drREBLx6udCdCeqth51ldrKKW/lea22b7fumdFO2zIwzAmZzS/
rNwjnUnWm9H/2BSYviloIEBGsvVB68iSKxiqefBr+FKALH05jWDy19XLH/7YTiEB4Da0rY+BuXgX
/CX0z3F9FkH5qdPRReDMrWE114unQ5P25t8wEf8BDZFByvjeNz2I1tDTTUeyCXMpHG2hI46uxICm
qrV4HCFKD/KtVyYgwqJ7VsUgj8tLAPZbAAAKwCV1Ubooigwzm5JGcOFEVuSmQH2M0kKUlV1j8BD5
2N2V+saKYSfNUQpOQCHu9cZR8xOGhVC4DIgDuR1AqS6KEzl6ZWfscU4vFXG2Z3z6x6/HSizDehs9
PTRlucfJzGLYWgtPKVFqL4ATEcXXlUVICLHd9IjO4KhO8aRbdqEcQ2v3+hRrwIr34kBWI87I+GI+
hXma39xSPATv6NRyTcrt2IInuyheXSCw44O028gY5wvcJ8sU0oF3HuggutfA4Bz2f95Dxw1eFtHJ
U+zgsQKfZKlsyFoYq5IM0+GuONt/8U67LAQFBfcArQhRwlwTFc/+W7Ato8cgG0wg1caTIpHUBadA
HFh8LrRc4w09kvQkAhL26Wx5fFbtDHTv6YMM7p6SMarLt5z37shq1qBKq9LBR7/Wj4uFmgK7WmBX
Gy+WfQTWCdY7QkRSGCL53C0SML3mmIlc1zI4Ngmzjf1OEoJwIITtSYmSvDvEx9VDSJC6IAxLN38j
zLSuSGtEcgduap4mBy9yiX6UuKo53uE3vy1rqEfHbOxiGX7BM0oRbAR1xGPKddSEqVIVenHh2Ipn
8fK8+kifu8Sjsim04QXzzLNaEJ1hsBaMZKmW9Ytbb+8RTjDWWrW/LpmTqlFtAxzS/nx4z9GLUSMa
vAVLZpBqQd3Sab0Cq84ozpQyuQnf8jfmjP4505R/qXobskzBDSVh6lmQ6cNDWFHfEPWItMd0pnyP
DRIKmMJSRIdw5bJ21DIdUQecIcDjakymxLIoRUTPIlBE8YzFb8Y222SVVF1GB2IvT7AcYLQ0AYRv
lTo+sLmJYVsSmsMMucD41eAbmO/cgfsMjHRIyXf1jSP9lJqIk71Oxm4OCPXhdj8IqGSpUZ7uU/cZ
sU/UnJyKMI3WyzvO02908ISvdwDkwXG8WpNgKRtmjk6+sAr4sA3b+ka0/blrA/JLDK+4mMwdEh1S
UnNWRlK7gXXiKH4xjIAv9XkV9l+4WWot9vFlQNdFdQurGXwrTQfc5WbiUe/K0VPjw7Zoz/gpSueE
fOR9ncZyyqaNMxdEsmaquYETHORrhv0oWLYRy76zSINkpNEpTRnDu15N957vBsuTEKZbzWXit5Ey
QxgqIg6rgyVQiYT5CUSZG7viduak0mhOjV40tWdbnWOS3y5MgMpgm6fWIIU6xbq6irUkvVgosFK0
DE1iZkVi6NJ7u17lpxjz6CJ5GBzLHq0lpfKgqK3VQ45Ld2v0L0R/u//T7TiSVF6V4oFT5/+Mxmar
NLArfZUcIOBhBfjuB0ttViz+fAyghQOh2nyg5P414OwM6eQvFYH3jvdXeHbuIowSw2RQfh34s+0j
qUOBui2XPcjdmJTGJdpL7ojP1FA24pDCxlou3FBHW/NoVqqYNezdKc8EF6TM4FCZSXtlo9hvtAQA
88TdUZgWlCFUmBbh79TWtBQRBr+ksf+OuKl7FCfkVbdzss4s+h9w8EJX0RC8BqVSqORMaJ5izxAx
sQD70wUuHCK0P8qw8ppaDePpZvnA+Re1ytdeQbasyhYtaLx84ofUhF5mkPLEGUIINtyK1pQjcyxo
4rZ5iUPuOzUVUsq8InUuqxNo0xbvZuo/812zbwX1s70Rg4jREZyCKhgPMnJgB63x8RdRUj3Sm1yY
I1qn5aYsAbjtEzbqyTgd0aZEEzjgqEC12jK7nRU0/2r3Sh8Wq9ajAjC1gvpireEsDuAXzPu5nAPK
s99eZ3ugK1ohNICZe0LyyDklA3Qbv/BlyArLbIbwxgCBooqaUYBTQLGjsw2bBD0XIral2NG0VpKv
mkE2I1XOsqvP/aMZFE+gNUNC+/AZW7AalShfm+gaIipdlhw/udldHhaFf6fWZBqSXXAZk4hRrmYa
hy2uRMeDolBi/ba1urYtPCv2mMWtQoAIeKXM4+4QlHwUwAQflN4eAm1xEIJ+0oP1fDfAhl+1r88F
y4lFzPkE0YvePMqZ5LJmC+nf5V/oZDSZS0cL6nyYfzE/4O2NPDDrRh5Jm5loG9eWgDU/v4hKCSut
H0dQOEYWasCoaS8g3I98NYJ3/PpUmSVffARrNxRIuALrp7a3sJVbgizjUMkj6X6Ti2tKJFIOnGqR
ALQs6lhi1W0ol5Xw/FbJ90bcRQo6eIvUhWnQwNw41aJZRxNmhgpcnOHbHkJdAOd5sx8uovsLmDzP
1Ee7TPHAdZevvaP1Ea0La63vglCyo8bpw7qclMmh3AQYnI0+v6tGWB56DBTUTa5qCoYyTPNSFlXv
hb6rRCtGH2XggVniCWVyqleHFxbX2iKK8hj/Er7wzUIy7Hn/TAwNnSWatG1/GnCyP9wjjIlQukZm
KSbluzaEPog7E8hqtI0x4CBvXlOciv564Gl+lNUUDiWss2vuD6RXTiZnwwSeQv37sl9GuokSMW7j
PKFTOuuVPee3RF4AFD8w6vmXdTA1vy4625JXvL0NswGlfw6qqqkc6VqVJ62ZhpO0KASULX3YJvF4
yBCd+OLzwr9h+sLezHSgZc7fXOBJ7TJgEZyGmGLcMur3QzO/nIWcwmvbJ80gVSROF/ZU3s9obU4A
Kiggdg27MyuQZklm1s0ObRqObDF0DlcM33qX7jcH7h7HeLidZaDJf201ms6nYDViTxYMJO3pkU11
A4AX4w+l2SikC1SzIDgfYFR0c+RpmiS/eEJuoiaVm+6xIhKAIOgvryYAXzmWWS5QNPX51kQ6uX1Q
IZeHmdyVCzHcZjgq8xM7vnanPznb87Wv9nA7HI4HbDF4aEnoz2Tga8pVMddRVIEF69B8d3JWL++m
9e0UUSrfisZ60A7VnMrFZvQbQUhydna/Lki7p2UFFmjotcpFztHWVHtxygKha00GYPTxWo0SWaBb
9hm0MHAIYF5ghalBKqGkTa3PQP5U7sZtbk2ZHi3I//kYagrOMEIIs8IBlbGD1QIWii/sKhbkl9lt
jcSb7FbkRyRZd1ETea4kdSnJWL626XFv4HDha28FDn1XqvbDoux5xIBtmUwW/0o7GS3oBDUDQV+D
3PKehYYJWIEj6um9XY40rD9RKI2VM3m34HL0Dl0GFOhWl1UjaWBvOZEboY2a7PG4Y8TGM6hRCOWV
q8WX2zE4zx95vOqRcaTiPb11Q2MSr8dbOf4dpo/mniWMBrFfBe+BHA7s4XRhQ7w/2a3l9aNprebh
ir3afVmvbFolkptonxWCf5zWH/W0fKZZaetvrgbuO6TcNZkBBSlFD5tkVaG9LfH4wNEVaeF+q6k/
h0V+gLYvpFpdlGv/BLP/sEaOZWvSPnREEwuYP+2X5EvFJPvuPZ8adV1w7xWnBEu+bkeRznl1qPaS
sfpTqMTDRO38ry4/vs5/YZ0dvthCxBt2T6W1ggaRToZj9r1zXi8Sd40F2PI97CYdVydADOqOFl3k
Lpy2Rzd1pyieREX7Sm/x6JyBMkBNHkVOl1T0Zqj1ItL/6Z87QcJ70hX4HdzeIieYXaDKNvJIjca+
3t52/ISVwfU+HWHBRkpku468ZSQKVzuw6YBldSqUV0YO/rEeHVrAjOb3aT/PUGybrnIaprKMe4EV
qCtSiEpSWqw/pG/VzYPbS4TmrOiYWL9vB/Iz4ts9WmimHj3yViS3pb6rUjcVIlbXKJgSdF4hqvP5
66EPbwABu9oLkTVkGIGPFHKchZrs0THBqS2FrqNDDplqReeH7LReLaKfabQNG2hhmNTfIFagtnl0
ARcdXSCWjUAHsvnim+N918frQvGs/4GWWLL+NIfoecSJDGeUPHgqUSTdkLQhuxhoWE8uL6B7oXGv
cg4hL409RW6peJxQA75wpmmw0gDs/01XmfF+3mvxAMGpjurKgyX+QQ5tzAKPi2AaGeCGccpF4vvw
E0Elip5HxWr65GwxD2zX/f84KffbEvu76MyswUapNF/EpGG+tNuG3b0/SA17oyH86v0XwE38konR
45majbzKt/Kvlq3S90riXRCkEgsalHvlD32vhP3wRXgVPa6um/lVm8PYvSC38gxRNryHec29bvPy
3lE5fRxihLalcm1hVBQaJktUaaaaTCTgctAGDg73uV33GKAb9qFzz0YerqvohcU3/NyKBsBwM7XP
NZEz6fFLxurI2KrU6/UiaNjo2TXdnXAEbuPWfGU/2CXaugya5f0L7TLQLSz+NhDDtQOTK3JEKud+
malCd4nKruChL3FQJD0nrBY6DC7qJWZMvPk6DiX9TtmnWYSoNE3uiaJhKyPqdKfKdVOEkvNPvpa6
oLxLmBB4WmdBFp4YoCyZgF27w6tW+Bzjt0FQ7OoH/NrdMFPlfE2gBdP3NuujbxpPqEuvgo95+Fgt
/Eu6Qv+B3d6/pytmC1xS8KkaYSHp8rzAbjO+7az/3jtyoYSvMNoB/RjcP3COVv3O5f2mAwdPlFuD
2k5g64bsfTlluGVY8l7tKy6r+PVenHNlusjVF1xH3GbDTwVOLHDowB0cYtk2T447STbC5USNbCZL
SRFIsXP/cFZXyKTfRQSoYW4HwVX45r7D5K5LM1Je5dOunCpdEjVFwm4eLdWhxhKpREgaNjD7wnYy
wueTZJpoyp4aA0L0kzKItYnypAesZ6eOu0lqm3VWQB27I0z7nkf0lw95Mr+bXosKuqBmjsCadps8
R0WyOJTj3IT1QZ1YoBsg2fkWEu+voSWycRxXBoHei6Hc7dZDem2Lew9nV+8pYMtKRRO1IsSHkV0K
nmlrDq7Bkn3yG7jPlLvxGu0KWadq6GyoHcTkElOJYdNnGAFCWwv+bd3rHYssIYA3TVoq5ojuCMpd
doPGKaxcTVDgZYDEfLSSoFBnMa/tmpLEpjOqIRveZhTFhzQ6ZpknERgm73jrp1LVJVlKLxFbCgSc
xoTLGUiEFd2ltvhXWmJGaFliWh31/y9JoBIxr72B6HJuyi2bYxop5aXHGOO0Uk6h7wyumZfSEyvm
2SMqYpU9RK7Lq4YjbB6D3EQloMRUKCBI7W5/R4wukuw6xBAXdW+Hgut8beQp9857XKusGtVENVAe
vXpK9YQaMI1MKL4/kLmzYtoh7xRhxu1wFrqGQOlqM2UvlEFMYPkVKVWFT1sE4sHbgr0dZ8Zo1IIf
V+FSeI4g58jIgBTK8pzzBS3So47IEAwwIy1vv0rWK9/irDKZLu4bN+BZZPWZ0rGBLbVa5pk+acXx
E8E9Bfwwp8NmiUuNc+noCto9ethOK8H3SrfVTIteSjXVoM1kyhUcbM2cfJHe/KYbCxFD8HZGKOVE
IhufSF4iBv2P/lBkGqvkBhLMFEBaVxUjYwCqnVqvoMMcuvdyI+Hk5w8wxBiQbteaPPP2lcxTPgp7
7bVWReYRX8PhpWIJXLgfgMX5ZOnnB8OKvrk+LCL/JvQVwACO0pctQ60Jd8aWLEmQhfpfPq7Rhs84
NBOn4/vRb/NwMGUqhPlvtmMRAJ+wtucA0ZLAArNrnlw9lNmqojfMmStisIgz/PIDIqwBncfXOYVI
+szgHsY30XODChg+k4TymLq3u9VDyh9eHUQE7ngnONpZNr41hnNOcIzMqytCFkNQn0REvl1Wr36r
RIM2l5vfeYmh0n2Y6ntU3kox5nrOeoTeCnmzk2+Nv4vUGkANKTExIPr6gHTUuDUHe4BtYxpAJlY1
dwlXkaXXp+hM+/1NzgtUJW+BkIgIEWiQLGvrXVHKzRuhHFRquIAxB5yKohh0fhNqEmnSU66msQg6
gShUl9O4L+1d83pLsdfCRcBw2lB9tAUjw4+gGU/jLpa+xUsmjHH8vr0l85owUCjKA+z0xu6Y39TV
50ra18H2PYbOGqVna87EwWB9KQokv/ihJQ1xtDGVQER8DcxcWwlmvR3anHpXG+z7RS6FN8dk8ES5
q0i1/wef5wtq6NiytWtf80BoirU4hgSwwlrWQ64SdWGOpTIkA8c5cgzdgJwVYTfrH0/1D2WUXtnP
aUlCHl+e+yZ7y+BDLHHvw2CZs6nc3VTrcAun55pU7R/aAYqWNG1Qsg63jrZyVaGAsl2QMYxQcHR/
7ABR8T7ZTIGj5yY8iaw8FkxZB2xkOsj+uxg/zz4Fb+mMQJtmdYv3fV21qmI61juYW9XF8/Y62tng
EcJG1amesAsSUwGYgA9q33CzIr08zzMzFxSIYLGZcFNN072g0SdFcOTnwcAxz4ufXYBzBJ99MpAg
uKmNpo+g1xEoiSnpTPXJVOKbwZIpEBWwh/m+4kmviQPGKZsqry6E87ZKmgdUoVG9aDwjtPx68Fua
y2YpsIZ84Lrd8v7G8klX66Z0r0PFzXNf8eEEGm1nYhCxe6STmvAvLYE0UcB8LTmA1D7YNCpPy+U/
7OqNCjOZ1GtZWlPwBGdbSuxtFe5zftO9HpgCR4OBm0PhTcGFwZsXXEP0vJ1EWWsseE+yg1Sn6zpG
wkf/j7HKQBd/kA3fNEVro0mBW5H+Ak0/9yXSqNPvkCOFY8329cI4qjgdyCsoLLXK95GwfOIWrL4Y
l8g18DHPEjRxT1gx3hrtA/KUFjnFK/ByflLgDIRwZnYluCcy9o/0dBfVmDcJ+TX/FC6Dd62WO0wu
q7gIPMtvYgj/peXccHYgA6Rgb9ZDJOkO2S/TeBlxH0JIimv1b6zSfTsTULh5KEO2GnaWCVDRe8jc
d5OJ/DBhyaQQZuAML8XAWwdUu/flbkkDXxZK5zsow9d7WPjKxoDwbEikAFH+1dQ3pBGez4+M9ONN
uYNBsVJ37bb9UYjZX9f/Yexrh4wF/PQL7Y51gplQnyshB58NMl5bArjPxG8wXn98u+jwoaUPemxS
4wvnMtjBA2er2MdqUCMwR14/p1LQumKM4o/tFnBkt52crtW6Mga0wDYIPDrZfUJcp922Vf9XjyCl
HNsXiVpbiIdpcQKJhkHk79P/To3TNqPvQ9IVjlWwRmGUBcg460maWDNihoiQCWfkAj9mjDry9t2s
bhWDIQb4AE1IkKh/JXfijRbWizw2bGDTN9mNtT+4XFmlinDMUVVLPyfbMQnZXg2L4vFUXFAXavYB
Kla9Vl+wNnPVKNUYrpZnRAIgAzCfV3aK+H1bPT5LW9S217uuqPJ0zF17XIjzyTXFUvSv6dJVAE/o
TSTk7ZGt+6QDK2N5aBDnB9rsRj3JFrIs+fTMr0IvpT8k6wocVmP7EvDqN9Z2yUeQ1Skji4ZXLTMK
cyvwrpojn669uBBldSK/OB25aGJiAgrQZQmdjpPICpRuyniBeqJZ03bgRTPYVNXEnUDSRcxGn+4J
9rmr+0bD4qb8hVmZ4DHw47ZNmepG2ZSZvL51lRdoudr7c5CFWt7r0xwDSHHFutMH7pzqBatSnVxS
d4mJwgUUq5/jEbAGgwjLN0sPczdMa/e9GR9jJ76QHwv6qdmYj4WRLH6bvtjVoD5L8hbWhDWIT75R
9qhkYdlMEHabsvuudkgQv2b5sPRh18cz7K3KrLdbxbmX78FK6gaYxE3krR7kb6aEyF/jyZAMN0+9
I/QSLgMwR8sC/9FzXl2MHsEZK1FwoYbzjMNwonQyOXTauKt6NgFjVdWendrLj38gaiq7v5szNgx6
CZx2KMNj1v11atwxOXKtTpnodvN1KKVDTrjlpJSMZ1B4BplKYJUSBI4tgpE6uP+Ut0S/cL9ZljKj
4I3lz4cRPF/d6HnY7O57KiIiAnYA41Pilk7ItWAQ6762gC4foyfZT7gWVk4a0r7V7qDmFFJfsCoo
2UFo7pDGC/OGjeMjj9iyd57lLarX5pyI8oaMWOG5hbA+qPNO0xqWDutUCwa9M43y1WzqAGfsohPD
ssnZc9UpbciwrfpMRGElGcnNkCW9U06dUD5Jd6V1EkuK3ULrMfjeD80zi/2Cm60EPs2YNX1tHSeQ
T91AGmAKIkBRAXSKpFrNP0viqB0e/rLe/YnwtmhBj9mK+0kn4CiZvEHsVhhfYo2XFO5o2R7Tl3Gr
+0IV54Tr32WOmB0iOnaGxfossbyyIddoCM6yERJIRZ3UwvRDHLEMCgZ4DZn5LXBJ07jNc9vbtUTO
ZWK/dLn1dEC242EcCQbuuMcdWt3nJqhZMPneses1fRQEUZf7LRYNpqa5uALEdpV1V4sjDWputh40
iFbBEgyUPeNXUGNSn5ES54t7NM21Gsa7Qi2m6wImHAlddgOvneBh08QfoIIe7Kl0GgPybQ5lE4er
9aTuw2BmkOPrc7Ul/Cq6u+0qf/ZQmpurw30e0eNI7Jll5Dt9Lv1j5zxX3iAWitR9vLDa1QT1qb8t
/RNsSOW2rjBjKCl6rvx7ib5trmcADzlY/D0MNLN1eMKaLvpAZAlAYZdXkrL4P5V3/zUteuzmKhqM
1BZidUdbqXhyveJ4dmY2CR/6M/yf8cOEiBNxfEX+UoZgAAH7R8rWVVgHSsT8sgmB2R+jXj28002V
7XDh+EAD6jQADRW4aIdk9zVvRgUcu6Bapirpnq2P3z+zO9tt30ocnK/WQthHsFGwGs0CvM03oM5g
vU5NBkv3YHLxl2Dchmj7cOAi3hJtqN8Q7pW/jTVznNDguSu5bJPJkDn2hSh2x5vkjMYSNqAupx4Q
4zwgrLWV3LissdUaa3b8i2HkiEVPjo/liByXGu2oECFzkgS7Vl4UlYnipf6JlMsJ0xtI3hUKMwdZ
mqvoMpWY9g48KUEM5oveRLWC2vzItbCklWPSvsSVAa3Inbgw5SEBHeIQlu67lSbOOhv7ruYIB32m
oEP8Nyh1zmUJq+hZELdoQDZxM4VtkgF0kwLb9mSQbfr8XsljTbwyuR8EOy5Y1m1hOoXyqVqt+Yb6
krPRytqZo9zPSm3KIuNcJbRW5+/2TtEt/CFEDCI9m//1HxN3yZLZJ7gtGR6QZMjsMREbcPYXU7E4
ZMVxAwsys0IyMIqeIzrRzhoGJh62RItRxMpP+E16lCcduTUI1W/0k8/rE+L8RCOx5OsXqhbeJcfq
MFzobCBwjC+H0VUE3lcSvOrrVO3Mmz9pvrlYYj/TbOAEWJwZsdU8ESJg2g8RSfu4GmAN7x3YaOMK
BUHdII62iKGjR+Ya3bbWVxxzePDM/BfjhGUuqqPE94TmCgNnKEO1fsRLq+IWl6RTQBy9YBo8Mu7Z
5js7lCMYHTGcwhs56I+pczNJd5ATB5x4165fyX9AfFk3OKezH0L1o24zK2vcRN3QYDYvOnS3dMSB
tWgfawjZ8JXvS78s93vk6dSaLjr7uB4cVS9F2X0343uo5+tSvFV2yYDAUWqrfVhTurfCabihbBfj
ttmsssKOglsWAmIZ2nOfYSj5+1h1mOcd6S9obMb8TwMihLrg0NYy2imupYYkGv5IgUOIr6i0kivw
87RkcRRgBxvpdS+okWtQqqFg051Ljq06YdI+F9UhxnK1g0ZnrjPXboOSVoRfIt6H1wtpmApuD9lb
JX+mhjsbV5g4AgT8t6Qw95887bQ5l4BAQ24ok+xks6dbPO6RmYLDx90NX+/MD/TKZqp74ib8yKU8
6eYYCQJAZAkF5O1bvcqC0UTcbjaVdREi+5V2uKbddYY611FXjAUs4moERkVnafJ3w7wSXLrb1NOA
4JfRGp6cAYO2sWuTW135ray5Zg9Rtb3zUHEMwBcC24n3suIijlxoN7KBSYtjiUWQq8st5y8l1ip4
fHTB8IRgmNMD2Wb+Ouaod5qfETcU7mhdmRRpTi09CkvAdZLgOxPkWRPOTUaT7dtxQRhavvX1gDJR
I3loJZTToKwbkeeld/t2P4KfUyB5SSdzjGdwT2LIDHCC6JC1nf8rQ+QOs0pP9HB7sq4otb3MXwCp
jTzTFxtlSqyzO6MLVpCxAJQcQX8eUrpREsd43iP7auMY2LnpYfYrIHSN3jrMvnmwlSRvRP9NpPvG
GwfKXIBV7gKB+MbmbpCEuXZIKAQ+aUGR51EUCDHbjjCqB7ZIPYjSa0SbXj7abGUg4MfPxE9omN54
Ipubxxm4XdRCxMDSAgLGjSjy3wK/T/KOKQF8tnDM9E6qbn4P/3zmiZxzPg3Zy/GtAXXRC59hAZc7
gdC/glr/z9fB5TF7ULMo5EeyNkRhr91HZg5iNadNnKgpN2u+ZHRKk0kIhJ9zu5ANigcVXX30v/T1
3gYTIwdVMKFv7Wn2n9aK1oaAtmWpWsN2C9fGgKUyJyo8mQbOdcGzuFYsvD8hRLCV/jFZ6D5x9Ho0
yBEVGvPFoZC6C+Tz4DdFAwDFHTbcnlkvJG0fdwoo2sV1QKNzGFOqqeZxcqb0Z618cH5oD1SCs4lc
ig9mawRpSU6dYj0ZXtRWOdlsagpUmb4pCCcPp8cCnnXBIYn9NQNCUx/bV3oOwCFE6bkstlrKUv42
hOw43n5xeR6FUg94u8BXctXuNTao9TCXUnXbM2W3Fu3/Ncq70NTEC3/w9gKXx6JDFbQNb0VOllrJ
Fgxvpn8LKaBns45rHIFovuMWwX0YXiY4+UE3WUkECgBCdBmw3wYGhw2vbHpjN/uwkGhNLk2TyyOT
MClw4YCWWdWdCe5HBJZI3L0Kx3BXVsEm3GlyCdgJlATLb4MfijlJNrgaN11aC/IRk4pmvEcDI3nA
dhHqiK74qpKRgsAzl2xnjf0NrbCmLBCkKrZy8oyuJ36de5qYaR8knAeqetEupFLCxnm3LTLOVMor
O2Fq8RSSidgrDj70BIc4VgACMaI2ZIQKp7ZHOk3/k66DLgkQVQh6sRtnngz4CXK0khaZw/4KwucP
LvMb7UOWopx7xdo5isfClxNIZhz3+LYP046XNMm6cF5x8XDlj9MqaeZutCi6mERq9wuZD/p1178g
Sofk5RB+lfNtY1Zob3oqE/LWokRJid/+Q3wgV5B/tfx8b1eSiSQXcKs3QdpJ4cfgUCrTedt/q6sN
EMfqJAYPtYMq5td+msWOps1BkqaY0gtmWTXWZ4aZ9d1mqn3NMVIP5i7oJ9AKZaGapkD7b6ZSM1MT
58pgXhhNJq06ehKJ6b1++L3S7yaoACTE3uuY1xLOCBZ/v1wcBom4aNRgH/eR5pk2u3ZwXLR3Ztrt
H6GMQ1oZBvDbfoBu/KD4+yjJtyZOBG7UcuQErEJ5SHJwHG87MFAVHBRAjCE6DgrBfTItqu5qi60N
bRGRZGnqgZNuXbPeKD7eccmFMrGQvHoc3JFmCo7Y4cptz/yfRI8rXBWM0f47jm1+1gtbhOU0az5R
yQKZsRGXKfpNXhXiyBlm8mH0DZ73QQmiX/Agi+PxopsNhAK/FFiVmdYfHESRyEBBVwk/JcLXcaiH
fFW6/9RdKMzaXeyYc547AUE8FAZawQZVVw4kUYnFvJqGZzdnCWp4KfhdyUxePGa/g7bzgD/z6N3G
ZSmEtpMbm0yt6DPWRhDD7iEimvmDFuSJHIj+Z6ISvImXyCJG1+Xr75Bbs2RxUxo5IEXizQv3/Cji
pY3shY9ObS537aSliasG3WOQ324Ocdn83fVq2QoJvF+Me+LKfx1ju+VGzKhZWIDQKUI7eak7WQa2
BfG59BizexXln3gwO8gRzhoZbIkml95NDOAl1yF8gmbuedtr3NtfShLwsakE3ZQF6xkTRzMcoXt2
8YO0V8TxeYVeJD85OubcYvbWIndfVaYnRuh1baqUn+H4B2Wk69TJ8DRlBtsHUb7WVYoqeO4p+vL2
xCsT/2ZEXr9MfjbI/FxpzT851JZkaTC7t5K5ZtCTfT1o+9KEd/QkhoDlGJjMsqWFxPwfl5fOaZFx
xiMENzuz2vN53j//U9tIlelNyG5tpR0eHwbd8lsDItUl2aT3pk1a4QX7lPZGF/OQmUE0SoNGvPjY
nVR9LJyyWJXdxmUSqroF1rtFdHAGNMXrEq5Rnl9DLsQWFKmeMhOqzZ9hcbSakpusneKiM11gl0Yi
Qunqer3Ih9+s4JKxR9FARPhgXRZ/r3LflbWvFzKOKSROBdshL/IlFKNCKa3O8eGh+dBuDfxs35ZB
7BcZKjXthJHDBmW0Z+tvYcmtk/5yFfhel7IKNZl4Wjo/uTV6wrJSpX8MwdkChElGcGOnlCq7MhpE
5nqCW5FU7gQ4L69APG5iuBG+DbZ7NAjMN0WkuqeDJnR2xw7xSPw+LNP7OSCG67V1yJJo3hhEBxWl
jEL2iDqi9Gnhs3fy9XOod4MeEr3LWdv0dpiSUOPDaqaLsXgCD4R5TPcXZmWylF4w8DvPPW6OHpoc
H75ILUhYfW7MiNc5mQZ2zHfWzKQ1kdulujTwX67D8rg66Fx1oxcVQBdqyPvOqtqalNKs4+fRczsr
rLPAWgSZY0+HJ2FTH8jxNbTA/pfsFOCH7KATelNTCo7sib/+E4lgV2Sn/5Qn2GZQL0BRH5k3StM0
L/9vOR2N+WqoaCsrsMAorsA8yx2uuvGIfcVEuFvkgGRH9446xKNqJnZqqJE9PHqkaheUtuCTtiKV
RC14EDdxyRK/Bd2xSOOQL8hB5Uq1HAC9FRVWaOGnzYDSeVoH8yRgVImQ0wbTbeHPP8P7iD+beUE9
osYJajLgK4otJEUgR0ZBSJhL7NEOe4DtrW54Q2BDjGoIDIYgk8fFgbRjejU9sg2R4sHtP1+ykg7c
j7K0k4m3EVB5YWJpMCrfEka8KZXsGc5s1UGrREaAF5ckKvBMW0Vl+HyrSq12KEZHmhc3TVg0EDPF
tVUkdceE2nbkO/X3867NKzaB6OYXBMizjdpQZ+RkwhO/rVKoE2Jqv9Gk6UrIAK3fItyif1HBSL9D
GYQkHrQFPW0EKZ2WXeB9mUM/YZ/lgbnwf8an6juT9hXi/CG1vtK6RRMq6zo9yoWrBiV9/708qPC6
AzZXZwFM5K2YexazMYSJIhR2WylqWTRM+B2MRhS2BnC+gbYvKM3xjjBwYEArC230zVYdpxZM+p/v
pckMimdG5WfDihVMH+ohxJKm8bFgi4eHZGHMvoBHfYUfwgcv/9QSnk9iPJTrE+O/rr1CjOiT56Py
jJh+e8ELNCv+pwkS17dv6kSvgf4hW5HNf/rDrYwyAiTbXnYQN04DEqPSn+y7lJEAoxF0bxNnKA4E
YzIYFQb9/MMsgknmxpyV4ndr57bK21Czd5389/oC5IjgeuE4GrEW8oci71DpGkRAjXQiIlBJgdzT
fjAiHNZY3bx0zIz1cBQRhtUOklAi5l9TleNds5oWojjE2AMXRbxIkwIs6nce1kbHALvVT6HsX5LC
wmDLUvjisUmp+ivSmAcCIxHgSJaF5FkkN4v2LVcqSlWHLSUwSN0URH6PicWvWeNgie5L22i+DNV0
gd0KmMbZxUfVlj3Chq9zqBoD0RXly6sbVmijpnLg2f3x4WOgcukPWZ9O7bdztQZRIV4sMw2/1saq
IZvJmVZLh1UX2Pd6y2JjxF2UxcVM/QSVuazToLwk5tf1nbBwyAf8GU8Vwrc8vOYs0dW23JJLVrBw
EsD3KCnmH9MYYxemz5KL+qNqgs7pZtkV1wE8oIUUkSbuG+0QmVRRp2PWVmX0Nwj+ZSD6hzvlYGGI
RkkhZTFpf4smbfRJjMA3dOy+tqSU3GutGw/u1dPKd4R3IjujsgsTRrnvJjO+efvP19+Icu3Fo1pR
GZOA6C2Lxjhcx5sXhFR8PGZXJScjy3fDKNe+ihS1pFssc7/V9O3RKJ/bU4mv3kelYexs/UTfA784
yXpjEC56+3l5pjg2Ib/9hYzKQhlG405emYqgn2xFy5g4fV0DadCwN/afVfz3DMjfzWu3mmsgjB2s
zD7eYFgK9kIz11NB2KI/0bXgv6vtmDlbnGA5r1AL0yiYqccLYz287Fqy9FNrKPUENygomUGNpLaR
ATttdGka7RlJAxZ8VpxPnrNXzydUMaJsHWP/u9YK3d8bs8dwdnp4oc5wCaOAxjpm0nn9FlP/fGSj
Q3jFq+LIwXZ32hGoEr/BY9aSnLyTx+7tD/kmBd4hiCImiEElXoJbDMRpZlL6T0QFprfv6u1K2p6X
Aw3K/+6MF9O+ex1j5gSWbtqG1LG9HHc6t3rzctJLDnyRL2LA0Oxet7FKRwb11PDUBoh+9GdnttnU
TJB5aix2HtGFzlQsy8gCABTifrciR5ZotE9dMpUB02Qy2eWLRMX2Ol1GD5/8SxSdLbSOEy4CPkhF
ufMIRuLkpGVi7xf1OzCcttODCtf1cgkNd7WupYGVz6j5Tcp+K0DnbLhBKCGtIVBnTNbv16X3gOkx
TA7VnPvEES2lOKvrI4NewsiIbEFsc7nRzXyrc01FvvC9Xpbuf5qv5fyPn9kqteCKtlLFx3YWYQz6
aYPaRZsbDUq1EReLhgd2ulKIlDYGyN0WMYDaNAZHtHtmCuWcIcTDWnSlIOc7IuTJVUetmNaIW5RB
8g2MeO22WNVsA3Wp4ixSJ2xGS9IxvnbbCCSgTSZgo5CN//z692Zq147SEDXuGj6hWZo0NvivLt8X
u3yIvsuGgKxrw+V5H4bkHNJe+z9bT+ROiK5i0hB60mbYWVQxk0kCpRKs5j47tB9Q8kz2UQn6iRCl
h6MP4vKZ6riz3vkJ7lVd5fO+WdZxHfkENK26mLa93QWhgF+3dhYYs7d5aDIogOF+zeL4SSh3kuM+
DY44PpNGvzV9Gg7y/V0tINlC68/t5kE8Nt3OLq8ln1/MKiAipc6glsXpW3DOo/1dqaaMSAdN+XjB
+U5Z1UGbkDHkXj7B8GxKknYYKnm2wcN7xl8Lqs2S8SxMEefOG/SCfmGjx8Lx5f6WGjomIBNBklnl
hTNTaTWxPJ5UrqDL2Fvq0GDcIdoMgZNzvAqIwuxSRIfLbGdgJnkMHgf9rXJ+hyMBXxSATiompQB5
d5qjnXoQ/Ci5qIVDPRWeknV/+Wqb+gebDFyZ1+C4iy6IT2167k3Z/VMSGZs+FTKt/146xweMtWxh
Ux6JsE654wWyGebSC3cQm6ceAeplHCRt3dwRw7iHdZYzIxIbtMOLD3CDGSk46ajpyZYyTi7vPzb0
CRQ4WTLWHg20yifCC9h07brAXE2KyqM+wiuhF4Gq0wKyfbBHEHf30wxlYbkWaTFYMhYnJUnrzMuC
n6Wh6KUgUxUWh4c5rYFBPC+7a6qXtaZC2K7f1QR3fFi692OhFCP8oS/eRAOlhTT+sf6ge8mFGjL2
wEJaIqA21eLSgiVmVBk+fqv5alk7DD6Ztv4nVrWsuO65QJHWxGXkWn4Omkhi+hoO4Blk98+lNqwH
TF85XgtPoy0v1DnTCNG8uqIJzsXzBa76GYCt5/74syurlkiXQz8I/qEf6gZ1r8KOVbXG+PybjEE+
eeAmbzxV+GkFfqACv2cvKU2oyFzwgcSUmg+Ld0J42ZcbxHugKkp/kxpf51x6riCHbGLYm74zIAIR
OqTJbOiv80YsTxTTQhVJGwV5kIAW+P40ALRUj8R5c6+Fn81RzxHKE6r17XE8NQRPA1/dwnukDdLg
u8V5VRxcmIuhMdv7BVY32yesmHByjpqpqJ2IrlAlaAYd4327HOklpgQrL01LTVc2EFhFqV7Jg44s
XixQ6b5lzaAMZAsb06tlPPqwhzuWy6oFyT4gIN/EO1Vmasz2drvaJkHstnTd0ILJNMlR0uGzgTHa
DwwzUq9kXYmOlG0pXHb8RQpo+c2N7Wq2ezdi6k0cbYDOla1U9KuUp0YF9k+u/T/CzqvwsJOKZ5kt
f3aT58zzV8aWE5g0UsXIM+H15XVn887XzxWRFy5OgVYqOsL5+hRFQLJRkj+7mdItL1O8P9kzxNIg
Pe+E5E9ePhCWCKptlQGx6PYqF/lvpKd6ER7ddHj6YNbcAW6VWrFevfJdBBF19qXGEkvC0ZnSYQb8
oQhJkEiu/zXMuKgqwk6yG52XraisaTVWhNj2h6OWDgpVYrQHKeJ3DRxQuBZjb2MEhbsH5adx0Til
PFYxPDJPSo+7jKXX6eM3Zlfr/9r8GTCSKzT7r2F6ZvX5MUFVTHp+td3Yk8poHm3iQF239/3y9ZrJ
6hGrdpAeeQ20v+LiEVhUsaXptfaxcX4ctKU7uNVhuBM6PIE1dfWE2W4nWveUQGmohnelv6ZbKWL1
oPO8WXJbER9+euJ5GS0o+QYSg0Yv3MMA/dd3zl/WQ8RLw4Ld13Us2DZ+NSlFtUoqe7SldJcsbhY0
nvBQ6NJJxeA67mYGtvr4SkQj1l0/NRoMcxmZq2ggwRCzzxpmwmZAhKQiY2OvW4AQCQ/kVLki9vgf
ffIm6vLt3X10nypZ/G/A/2P1epM3emRYt0oA6TutnZX18FUUnK86SQkQ2EtupcH5x9lJPdG1ZACI
3mqYKWwMOHZoEM4B8c5ZyCFEhITJebcyaY71xSczM0VTqnn2cdLIbVFNVNerIPB3lKVip8mT3phu
qv5fjkf4EV+76XeaLggTaFvkbRqyKiNGPVIksU7V8mlM2hdMsxjb/bTxvqwNTGbTPOTs2Brg2J7B
xMeel5OZeJrJqe5OE0+jGVxYMiZR5xa9HWVtyq5ju1LcJ+ob0ahce738xYRatLLVkDbU8CPLpOpM
6O67iZu4aXnXHJs3BCc9X65qZ8RoHQeXacU0CdhEB7wDA8lMTiMFNzToTJyrZ2HtWcC+LZOQCTaZ
TwuLZuOkBiiv5A7jCmoBPrWHfHBFAypvlzTjDgecqPn6XIL1vGeTZ3tdPv/YjBXzro6iknYxyS6N
J5Sii6iaiQmL30nefmYHN2G2xAtWNJt7CV992Jv87WhUfJSeBdEtETr8JKVk2KaED/rw7YEOngF2
EKAIQjF6KLfAB3kbGqrWb6Sg35N8wBwCRJe23JqDHWj8E2T9vLm5k/BY44scsZMTFrrbIt/oY/cr
CGu4c0mg2VxyFgaxAn99P1y/hcKJsHpY4sU2DXoT3ddYyfgLpxHJ4wBTE+MpoCDKZySux4HZjfn9
rDpT8bdOa++2LWP0RsLqs8mZP7j5LPvDMmCfNIEI2jF7l0modh82f5pM0s5jdfg19hDGGs/ljOFH
fm0tcg0SkCvsvtzaFW4kHn0IKHbDVnTUDLaMzUA+kFoliDR3SR22CSFW5yEtQ36Lk/32yxKni9Sb
RrivWb49RQlMqGn4tpV99k0bcNgweeSeSJl77E8+PtFEuBSxmUgHZFPjmEUZiPnlOvlEt+oGH4uL
uCzL/2Dlvylj/YfIC0Ms0BeXJrra46cTTDFYNODqZeTPDXJaLdVI7TxqLbS+mxfglc1X3mnd7js4
M4dFg/wPUkp3z/BTUb82lmcuyo5H4FGJk523Z73yE0M/dtr8/JPOnNynktmEsX6yUlpfWyfPUgwc
5atr4lU+GVgy8RtuccBXp+pkRHln2gWM8gl9f4p9liJVuI3c9r1gECOv2RE2f+knNtwIlaWHreOx
xA2JLVYoFVw74yF9O9HSGTLhO58gCb/+qIl9GCSgi+g992kcXpVR5Qfl6HpHCzJltqsbTqXn2A4F
kr573k6iC40bBZVmGbJfBvTtyKowLIj+rxrKhtYubbdU+U9K0T0SSiyI+J/8hlQUTJsMHJwM0Hfp
YKuFJz6xP6nbne2+jVphAJakOwVIQNQLGApTDNoB5sRsMoZNx/fpMin+x1Fr8ZkT9/UoXvSP6MQw
GDhUWXkkDBGfN9TYjaALNeFDECPa2+k+ZPA0i1J3n35e8iwW4FyqsC4rrZls90Q4+Pkg6Ax3EQKx
1YWHfdSY5/UTVzq6Qn6mj2y4/ofcjg3Kn7QGp5CY/Z/vGvnDxA5QVtYpd51e+7Vc9VvtoQAPsj/0
5tIL3J+y+8MN8Ck2Ar3QCvBxXd6u+qnfhqVKsEJpEfZHRZRAlmOoufdZbmy5BKEixmclOQO6hbZI
QwIehRKknON8VU5CTCXjtVAsof8H+HFnVsR5OasaLS8oUw2dFNdwfrwiuEK6snpZDORMGzpTJWX1
Ebi6vAUCzn8FACJgqYVrwctKxvdBy9buAG9qKFQHZSFaUZmQ92Bd3e6aCYzeJ7GE9uMLe+gCyFhD
gs+oKKUu9n9EmKgZT79OIp1dvBF9NZsJQB/7AcolJcGNeg8LMQhy4hDywzZrzn2fnmarOMP0g0sI
thQN+Mp2kxkZrWiM5EFswae11e9KUf0I6l8ilYz7e76j6OnQePEx9IIT7026IVvEt9qNm9StMR/h
1ttcrqz1ESFMFzF+kT/OCekHIfbueEwLwmECfgOxIDcSP/foJpfJlviUN0isejxr4L4qKt4ewq62
Vcbg35LX9+jZLns5/Bysd9JBN7OZozTgLlR836i7AsXVT9T9Sg5H0iiR0w2XQtBx7TlNvJz0ZXkI
rHcTq8DDyYjJUquT83DZS0QlFd5xcvH3/rkWrgrOvnMP9aDTF4paGqnceoUhSDuvKf9shsVeo/VV
KXo8ae0+898uuR1/iRcAYJGyK3aGiHDJrELuK8jMFDhOQTD+7B6audoOoJhGiTVSu52q+uegiD9U
N2gX/FDtVLt6cSUwyJ5A2hYLGdZVCYp0PAK0sGoJAMQdkmccJLPYql6ZHtNiIXJhRYMX1OJXd3a8
Z2fwVlRhqIMPRtCFB7DAE4UQMgi5DQNSHozTjZ0E0J2eOdnrRIMKGw9Q0HtGnWgeljbUDVg8zVU6
pWrEkYgz7UBPkRMU55SYqzpViOynbmMB3wYSN2PlU32jkvlCWZeyoy7Ayt4hiin1gsrjeW+iVulZ
MzpP5nGuFb7SHeOgf0wTp3lyP02R9hPtuW+0/OCvUTfFgcq6aa6zHipzcFwA2rVYcHM7zcYqJjUO
673ydzeBTDAZPkdlfvGxy5P9BC0LSNAQKma8gloYFZR/76eu7nvzYi9ApnqnenP6qv4XgJR6MjYV
f75S2JjOxzO/j3a0StayRYRM+aozUebdJidkbKu3w/pVBkKqDyDRo1LxNDUrqTYW3dS/jWKZgyE1
EKqz1Sj1r2iSwpctYQkdLNi+Zqe7uQAqevXF61lfYSWZ/ANgZ/6RR/6jI+kqJt5RXBDnXgYkDHYb
IXpYnp+hnkl4lnsmH/dr9GVaQoxfXIoD9o/KVWrewOuBu+m9zoKIpwsK6VlFQTpB21eQdOGIB3ZV
yYWeLMsLZD6nDKpAg5fZdY0Cye5ciQZdf5hL5ozqTT+v4rhYgOHWEAClsIPVDSQGI0ds2GozYH7+
Byzsq+aVJ0llkYPHHs7sbPJ5FtNEhHTlQJ6t6CJA3npBDHJKOTqW+4XYQ4cylduw488pNcetQ1sf
fCHiwGY/CHlfHys5irgY1z0zq7+bKr6HYXZPPLlNutD6I8jEbjiZyeM0Ct+1W8wRQXYhyRrznGeR
uLjhDG5wdFUKxLmSrRGiwYvm4BtHWe9e/CekF1/Ncj/yGFJjO2lW1CYwMKJkQtr6CobYudSwmTdh
olLL8lf8NI7BCUogymbuiCJtGO1Is9oufVUXB4LdBbqpOgXE6jUXto6fu4b1QyZtPO7nJOC1b354
+g1owLPof0oMxBNc+TeDqEe+IInQGSkDXfMgod5HsDiXQTz/yoZELI+og9jWokOgcpnRFrNXjcxr
GX/ly6N2YT+q0S1poxxp5L3GYJA2gtYG95uTXmS5d/zUELdjomLCYKRf7QivlgiJIc3C4UHANPZr
KUfdt+6fWCukW4fjuG+uSyAZoqA0XoCX4a2vkxCaTO1fmXGuvlV1kdwVLX9sk0g/LgGgPhx/bvxu
1ZNBvsQ4B3CRb1YtzsZ/egckFEAgdnNDfbePHP/+Ab5CR1Elkja0eKiGWCX6Bl/+C73V56+APYGE
gqBvyPj+xmjbGGkFz6yq/ytl0dfBThJ3RrvrDzIM5muNyHfSGV2g2z3WiCUWh5aVgccgj25Da/OJ
REweIjYvMziHrSQpnP5LHBSidf4GH3zirO0m53C2/qHC4Jr74bboa055PG+/Cw07mEuQ6bk/t5Pm
SkQutyX2OAy0BS9GdTCoONu0UjaiCyImuNheOlJmh/F7NlzpVIb3TaE32sGfyaZXDQVmLKgca3VS
jbDBaq2irfu0t8wXkod8qSVEwtAnANHC1ZyC8b8qu2XkOoIRDjHf3k3e9Q0kJRgIre1C57U+tEuC
W5Y3+YiCm+Dj0LL3wHx+i1BLIGhB2Uyr/AwD4trwsFC5VBoC9JuBCb7XpJM0HxkoGU8sKWMoiF/C
Nk5cwmendF5422OADR9WHKoe0BLkf7Y7bT8YbXg4qxxL3a4/O9o4oC+9M8LbQdbSJM8G0SDi9ogg
aUYs7epZgfYb/fzO4/vNh3dGExIbWlflN3shF9+LKQaU89OpGU5dybvQN4cAR5BQiI3cZ80nO7Wf
zInT69Z8II4twLdv43NM7E7jvZbronqY1GoPs46FQZX7i4QhtU+VMrVI7LotBS8wB8SHOU0brt6e
CyUz7c9+RWimPCBUX/HSGuLXJE/9H1DVNU6d3bATuWw3Or+uIQBrPHPqbs+n1veyH5wB4LCKu9PT
cYmHWHX2ca2ha4stQGFB4haNFqZDxruOVrO37+sW7QnRbSmOMYyXkaXf3bd9JuF1da5pZ/aacErm
i4m22XglLWU34788OFwY1+MQ2ZEV8/qOnSh7l7gm5aRtaON+6sC4FEXe5wxgkAhLLxvGukz/7IJo
8HeEPc09pQIN3RYxhELXObjniuFLqSswNcvJpHWxO6tpgeMqf/xDqP8NOrk9DJ8ZcldpRsjbDx0B
ajBaEFe9E8r7jlvx7ZPdPXmzCmsQaaIXnSWGcE4QhcrrNho/lEQ1daaOD8mMnWywOjtSt5D9HNrB
aNHrY5K6pN13gAyZzJjsIahz6djBQ4G8qiCP3UVAuPO1ZLpBN2D/g2WyGNOKaT9xOzxPSBwx6bay
BTgNjduJRmz5tTdVu57rDRhzsnzkwBX2BXCN2BQPjy5WblfGXzGEge/T6B4l6RL+P+JxEZ8QXhRp
zYeSyabgQIMP26zdLfZaaWzAC3nj2s438R2nDnDcGQPnh1j4G2Eyl5FZMthi02zIOHr84FvZps0x
X+JY5o1tTYOHjMEZx4kq4GZMM+fJqWTTHobdm68rqkUEf8lbz/oYSa5zHHqSVNAwpiHF+bkYT0az
JLr2HZtsP0QWT2Myr7XQviB+hzaesjI1KSzvXNBb2qKOyA5JkRyNqpWw+DmSyEfbqpURIc8BZLp0
nTUOVdw/Vv6cxgCQ+A4SuO/96PhjfQQ1ClBMJWeBxeJdh/P3blBxt/OZNhL456z1WAx4v8cKMJxf
RIfug10vK0B0IBH12vDbAw4xyaN6bPhRsfZUIGzLoXxkeHrrDcoQ7f0qio+0lAgfQGVo7BGp9q+j
dnDdC6Vt68BWUv4/WHBaH6b4k78QDdh1MQnxEozfBLvb+kPonXx5oLQt4ngD0m6o82d2BpMJHDne
VVIpT8mVrX5vdcyMG/O4SK0ccvQF6+5HndFPA/3wImluQJSDK9cqku0I8PiH9Rn14LhnvKKx7MA0
EUlydh9frsVXeTXQAn74aZVgZ+DzSXsGdEopkErA+8rPVmrD85pE+HgE4hczdL1aEABxGNq802IE
H0j1EIDoYm8T4opa5Vxk/KGsV3PYEZyGWmaulGxiOWICf3shWbcae6D/BnVPhSacQtrcqlzVBlZd
XnWN8n+D9zN42vtpxOU9nikgeQ1jNNEECBL53fPWReWun3Rbn7kFFfy2ZRGLy4biYy7r7AI95I0V
Hz0VJy1j8z6rgSdFKx+GhI6B1cunJJIWN4ArC46EJY82G10fJhKD/TWUIhXwG+ACgNjfTkGANxYt
Mir95oDbXpC9qw9MEQXwqj25diTSPD/nrqVnYRg7yIS7axZkd6kJl2R1zImmmoK3Xj0cGKG4wXlF
E98jYQW+sv11r5s6eeuqrJWnk7hAAgjcKmVhUt8r6zG+ekEAkbnMwd+ucOj4xDzm5u6BV2CUd8vy
25QvZ6aFyitqNDQtYfMX7FABeVg7BkmD7JG5ZsEkhJd6pDkD22h4VAA21Z3Uwfs4JVcQku2Dkf3n
8M6MALVp56qPoMgAztfqnRPZ2uAlxFUvGGreRe9jw2i0GkIGm3kPOZRZTRiTT2Jpt1ZibYQHgCXz
nXu/zhIYgvocQnE1wBCgWsJAX2Ad7IDW9jU9WF0sWZvxFbQn3auGjWpwXgoWK6n5pr7647l+nfKx
50NOrZ3jcvpw7uqRRIwg/LTZ/+gKX5J/e9ABiwlKCiRFsK/MdD24PNgDftkP9+YPVkSTMUdWO8Oz
gTcUMiHVglUxEetwkcRpgmnkR9eoJDseNSjpxpJT6rKCIHQIFTED0rK4z5rz6Rnf9zQjGS6SdCGl
3PHZwaIZNrTMRdVg+FNCpg7uwIIWugyPOcG6R4ElsX9qiMeGBUr/jL3eL5uhOmT8pWCB+DTT+Xap
Stka/i35RSlKPQcjlmKVddu9aZ5j3dT3t5uZxdhR8t3d0eMQ+ho9OTWJ58FzVXGOGu1WJUdbN+xJ
6v+W+3v87RmtrdnVEHlL32ipQmiVZpQmKrD4E+ULAdU8CFjkx2C/ZlwGm7vufT7t5sJSHSlZJ+Hy
QpQniOV5skxk0/LGAIyaRM+GnA/5JjAmWJQ30z0F1SRuV8m/As98gHAA1xqRBiLIlq85vxzEqhQd
pf7D2jLikt0RY8Xw+kNiheozS/P7PvY4dtAn3UkcK81Jt8dEp2iNaYjMWKnhZfbLkQOYK+xWaq6q
4A2fX2C8FBpqWTOvFWOo38RC/+aDZzAQKS5iQaD6CnIaKa6pkEAsqc3zevslRBgbGJHmy0CZ0dAn
hY0jmxkYjt1KlUB04uU6lbAfUIa7VGBd8pp5FWUGNuE0lJMVFabv2EQWh2bs2s14Dt/SI4tWM/iT
sclWzx2qnqRFwJDCIS+S/chnXW1OdaCJ0lHpeVSy0C7XnQZhpA2AXeadT09L7BiYxJsC6/5CSX4z
qGpwIc+Rq6/XTVF+Yn52ltbqTzVMuCnBti2THS1adG5QhOyOSG7yVRuooQSK3Fyx4cDkRYJZciyA
OpS9nTQI1LEDLNC2MNkC8wAJkGSREFW72s0RaAXck8iNs9Ka96Ujm6OgFtfdfUZHKIfTBMcUeEVt
XdsoNY2sWUhFlc0rH3DPyKOh7gpZk9Kh/kgmC7t3G5U5TMZOIGNon1e2j1HchSGFOoxGvWAsBCT5
TwTgnpc8TVX0HRZxgujspWD2HsddgjnSjxxOxZ/UIKnHtbTX8GCllhXFhXcUTcOoXcuYSJGbs8lI
f2L3V8xadDtJ3OCqZqUDJ7KKBhJADPbeNwP8CnOKi4jJArffIb/l6p59HCQW233N/OJoLb0rv9k+
AkdDXOdJN4apQML+STsstYyalICCYWbdGJN7zmCHwTmU/NMm93VLUNGBplN02A8K/ghja9nkjZKj
7KbcjLVVp3pJAPm1o4ny6yQ8a/CXnnPWR7BxI/zIw+AkZ5ZyNBmX2PQX7QN7k/i38SfVC9/xQQWK
f2ii/T/JGO7bZDEIKUlqZTZoix8Ecd6bHpeApcplIKsk78SfVqGl5LIyYtqR5qYkRudWO/uBgT5G
GbNRYvzpjT9/ZWfxarJvcLeaEgd2BvTavLeVDCFJcMJ2ycGcsmRhNz+0n7F/oEIQPobKoZaW9U4u
wxm+EFscnDXCV2JTobidmur5qiIKL1yiTK+s1FenwR/pQNFx7GjNXSU0egl/TMNon5asxJFqZXrZ
46tZtGz6FJRpZploruvl7CgIXAdvUP0IdpSH+PpeOsha6mgDCBYAWVlCXEM3z20b7dzl6zcV2CyT
jC5mJRWupbr3zF72CHn9jlK/SnEieE5MEXPFgOfb3zca4mbTMWoFA1IOBDfv4fPx2a33Wp4TX19X
GWxKdsLrlIf1EulIxXAvwy4XRG87T5f6lw7ousRL0mRyvJz9gXIRfGVmoZy53AHM43vHZ8ud3guG
3w+jvEeomfD2zcgSnatIVq6WrCpQIZGKS4jDohf5ORI09FBe8yrkmQS7YN3czSH3F8Jg5hDvnEqV
10LpYtAzigqgSDoYaiqKjAVgxfSJcr8Y4A/7ZxT6kbRwkFi/RJvCLBjGvvEYiJ/1gwm6A+ZIaBia
ybuH9pVZIvzCuhTWkJQHT4uZt7ZdGW/G4wcHElr3ESZ9fJjfrOBzPnbqUPNXzM87TybtzNBXGBlU
56c4L/8aSbC7bxyAa114voKtsOYd/q1mPEbwh/2A4Q5CWKg10Nib74D/Ce7OLZepg4XGIJBHOGJJ
Hw86qOZaeLdtQx7njr9D6CvPZZ1Y5aaSnAV1E0YCGXVaskvGWqoszn81GlfkGZkj8zoK4Ezymux4
iMj6aLUSu/1vAvMfth9Bc0DiiuliURRTF8s7M0CqNBrk8VF9cB4wk1dVDXb5zVctyFVm1IDhAzF6
xN/ay15m5rL3vFW12Gpz5q8ooL6bS9gZBCqankBQLnr95u+rRcMglaxAWwCZR7n9a2a+2d91k/eD
iEJAsNeOVh0dj/vQmBibWd4Lwf8ma6iYrznjmijDbXHfjc4HdwILJkoi3DDTBOEELL2pzNhiain+
htF9/LUqz5r+5MH4KEQ/yrPdGQDyG/VwNs3HOBYUJFUdFXRwAzEBgerEAMTib3oThPojjqvb5S53
nugfWcuk0/uiLrFaDbno+S8yYPgfzGELQek8lHgceKGKISzlABAmrpCVYTRa2K/dbErY42PQO1+Y
0DEKMbLXmEwIp7u3BNQo94MuPE+Hf/d+ne70cUJ51c9HfJcmjFXmbZQH09SJGXnEdPSKzluzuxJ7
UqiaqGHvZ+BW7dnA1sWEfv5dyytKsSumV9C738hkUei4ZWojWMb1gIGxgMMrHlGBvwYojkZtCRej
3U+WeRThzKHqzALe8Pppbd77glRSr9q0ZCuS7jjTrl/Imx9Luncfh/gckNnUgaXKuumbmU/WK+t4
q2g4xCwDYJ4zCWF10/5+r/0WJSLafVbfGM23BuVK1MIgnIfMvR5IIbECyrzHv54UqcH3YZbQoH8L
j3lWZJWju29xeAByB3WPvi9XtwJ6gIsoWeeU38WO090P/r52XjKIlHY4UyiwjulGliauGyIKrbgN
Jp8WQIr0YDDFhG5rAerz1G1X9iQJlmGyHNdMAfzr+lT6sVtwNmDAeqpmQSO2l3uAazFbrg3aA0Bc
KgPv8Vsqx/AbBDXt4MLwF7CAGp+QLy7tBYYX6UYe0gXkBZ6e4WxPpF6v9u4b9XmiwafAfKrFYEBy
xxtv0dD5DAuEcwuIMq1pdtPBZgLV3C6q8fIgHTPLqY95c2rPWIhKDusHzW3py1axKJSPM+rDb1PD
rOZ6+TiJBtg+ZczN3Uj585Pxt7JStfXTQb2WmBiBYPklNsyMiAR7UyGPzGuboVlrlCK/rRNV1w39
+8eFoMZ7wZ0+GTb/r7WW3ek4AXS3rtasUSEx5RqyiObxkI/OdYjYOQ9Epewmm3ABYvzMwVQBObhz
Ng80BvP211MkNG7HGTRVzBwIfJSSVhr+MbGIO4OA51ISUQpzjAb+iQbgUSa8RJs2/Mj9pDs4eyj4
0mk571e7EokqeH3IFMzXqJwmFVHagQyOgIPKBX7G7ypmsAVqDsRy0cgm4fdBWgY/LVv85GXfV2+V
Ch48BfMuqnPDj7R+m4c4j+3lIlVsqpdXqlLrSqMwcuXRLtEpwpa2A5rS2YLwwnP+GhDlZutisQI1
+V6CIVSBMuk2zFfQ/F1k2KGuJXlPoqOIpd11t9z7kzwsVj3pLeNaCXDLZDuPgckymVByGH+6/Lhm
gwlAR/Rs+tGSQ6KBtrOMiXpTskuWBLVsLTt0F7HJdnAlBBKPtKuCvF2nyCylr61FpzDtjhYbJmRx
L9pIcLYTMD9U3ybop/ZVjSA5+jsWBO1JtmSAtKvKVHAMIXoDMRzFwJRTCRZn/EQfmiX/7fcBy0Vq
i1yVOIPtDsdyAQv/r2f50iLF5CzoNK2sYT92Vd1EPBa3z+ewClEM+5vuQAue3zcT3uygoVDeKrsI
x4BMYgUC2dmb3gH6ctgYh9U6WGhgaKfMYbHcgwotzJomjoQ85hp4IMVJRLt03UMZM2QjrfEfzeHM
Zg6E/ZSuimq/7cQfhmQ471q4vYweJpuvrV2rAZDrte43rW3KLuoQn3Iir46yjL091745h0ofj7Ne
wTCW33dWbb2Xl5A1VBMfsxG9jGRrJX8wcDtsJFuFcxQqBKldfOE4V7wQijtsI4LdWkvhKObdwIqn
eUbOfhsECxgsM+nmyC9Xi+OGKQMj+y6qr4M1eXny+PGZ9W8YKfUqNWKeN/Cedgn9gi0VoZQ4wgmn
5U7jynllL2FxWvfmh/qyxa21J+AgmFyD+asEICqHUp6lV23fl4c8ZwzTIlcnSalc+I7EFzS2/M5N
sRkGo8c4dXNhcwxtREGGhrEEdcR9NkE2nk8ULm8kb5B8IY52UmDs87ib770XwX9gDkmIkiUFGIcs
9Bg7OJQ3B+cGDOkvIURepr91eNfd5O1k2ptRvoZ/NNvdHUyQ32F83v8rYgFbXHG/LwXvE4nkL+2c
LNWRdaJ/A1mjhYf+HMdC0tF/QlEFb4kuq1Ni2/66GPyxeQ7E/qmbIgbdjf/9pWjX3NtnEZA4T/yj
lMTjyOgLWsrEOOM47ikBgsBFmS+/xNPj0q+TQreUsr+5FYLds1t22lyTqbV1/xl4z+hS5KDx7pdp
LbtPy5douB6VrT1ivqpp1G5GQQw60pWeYnyLJzguyyNDRr516LVb2tLp8vfaoWNFU1jNOImnuFJk
PLGCr5k0wRCqUuKkhBOiWjK7jrbC1oB9Fj7Bv/86X0Lph0Q25+OUVDdSZR7T4AlmLrnirYMFprXL
wLTDW/pUPUzla11DDc2LYI/rhARMYANFH+lakjT+bN7nYZ7Ua7OGUH3DerE409MqoFZ83UYXGKTX
bnYAKWCNFyl8p2yRbJwTQDM90kIo3DoFgHy+Ha7vP00fMegXivPOQWPHf+iLAahKi+f8/tjdS8No
QUxIpk54Ub15Qh1FECV/f6YP2FeGc1BWwRQQOjhYWrs/foJYl8fx35l9SKabHXxHhmhnqk+UV1V6
shcifng9yhgVSeJZuCbDpxtu8WndGF8EscWuAt1K43DNotSMPnmJNL9Jf/fmGizW98Ei+XBarR0Y
eGahS0/UqPOFsm7hliSJhxhCgkh8J5U8MYXboatHJlTGa6YxujAQdWJrnaTpDeHcIMn2GazhXmw3
QJVi1qAWMVDd6eZ+ukWxy38yrvdbctSy6jm4nSdhiy3eM8wqNRr4eoo2R3roBsTyqOCqB67cnQCI
v+qEQzArNYGnynQK/Nij1bLnRPuq+/2biVwZv8cJKmQhSVvuq+wH1MHuNQlfYrEegLiR5/C2Znxw
+xquMyNdwEHY4pPx1+cfVhflz70429MxeO7v4R+haoHRRQIew8O54THwrZ/LaChq/AJMO5XM9c8r
VyF2Oeul/Xksbxr28ar2vbWD+6OCm7DhF+KyDo8N3/5tzN3jJj/GyBhuPfojjlDw3RRWrNTESFox
ididSt50CLnorJOpDtQArLrP/zYi9FBFjNviyrEbdx7bXHVSqWeP+An2zcNC0isHWbK+zraybuH/
hrC5GyGP7EPibiP6Wh4wQp+fu4ZNsRYopceOM+hBB712fYPxWKoRhb+3wfifzcCElyof0DO7IsYp
FKjQPHEFtuwL5m3czs274JQlWiayl/KtC1TXtXRlfTk6mIzCCYSSAPOwBIIApdJEr10SXPfSHUm8
YseUEWIvcjBPqw1a4ZJIhQuF2Py25XQxeLSVefcGSvGintVLj86ob25jDjeC3x5f/GeJicsJEweI
yiqwJ9QI6+7iD4UcGXLLQXLWoSX46KxuRTDbH8I4a8eURGF02JI2cnW5/OT2bWrO7ykl3xV62tUt
ZZmiQ0w3fT/oRu6Z8u5WYqE7QV/cNkqCf3aKyHlr5YG1ODd2HgYqLpYbudkP/7cN+3K/u6+bhHw4
CJcSGSvxH6CceV5vSGUXwFr3keYweH303x3Z7Kt6kYfaPNAHrzH1y0cAb3bZGRGuLBTLzyA70c4l
OJ8Ma3CNhdRWAEMjPbgOtEEadkUrKVu9tm56Uiiaow8XxyQOcMchAkhg+QGbAxjBTljpGNmt+91i
IbiftB139+2hNFI/TdNZfIFN48QeqvX7WCvjSfLew1gPtwB+uOyEWBE2hvtAnq7Obw2Z4MumqSIo
YX96LodWA5452I2oRXF+lG3F+dEu5xtbTTpwfu/1+pY4pWzZQGYVPTtNFHZkKHmcLZhhRGjSYgfP
TVeW9FnxIq5BFADGMEEJwPrbQ2Gbhv35gfBAPDgHHMaevA+8mUQyyV0sscM9NpOP+d7kgyRsfO4H
p8iLD/YeVvdwmLLDuPKCXLLTnqGV8cA9buuMOpbhaWzcNEPvmKOeoLxBBRZ7ZD+UdG7gTa0Z5C/s
BM+RSgklF0nrnl7TGkDTp3ulh9mTfSq0NUBEyIH8nDRvRmjBpxCglcJe/ednoGvJkTnTcilwVv88
8yeWmUs5Wv6Q+CGA7PQW9QnfXJNUCUNGpB0J/iSFzCab8CZCsiTtWHAZMrNI8f7gzcC45JZktbNJ
gQgPyxQ5swYTwX5/alWBaN3a8tzSpbxmZyNb1kPzo+Ihub4no3Xuv7H9ksTHu5tss9ttVVctVrMI
DAvAwotZKcFwJvep6nqlaULtI9mZmyUHwjdlgsdti0gvFZHuAEce1fbc+oC8me4YG7t4M0CTYGUp
rguROOI9Ut5VaWQoz/0jMiunxUXNHmZooyXnsjH2hmoD6nzAlSSZ/sJsSjnXiFBd7a1TD4zjiIHk
md7yEZpYfIMky8YQhrl3vgl/F+CSbNzkRRVUSy3NkK5SdvzO6x5BWWKXdrcBPMsoYJvRgZwDTgiP
CunHZFSUIBGLtmsmhF1KoKja+vabjz4Wa17EY0a0sA2iQLo+iGEMShvegHD7J6XyLxogkVFbiqip
fE2V0YdyMT/Wpb3gjwcMa8Ap1VLwkURvWmIllF2xhyWMBPWtnldtGiYHdRoGWTHiP3RrlFi5xlHd
/LpFazdSi9fuZ0qQ2gRnNxSbHbW4DOPoVn/WWVXXaLXwyRc+5RREF/SZx42PQipPVBipLCrf1ySl
j26h00GIDUsjUzYZFH5EhQLgYPmHyhtpCYvVLpVgi5kE3//V0hYzMju4/VR9MQdnCoaNVTuBpOug
j6YLg88bjIVP6PZxc1yAFMY10s1Rkjh2eKLT5Y8vEy/yJDDuubfPovShbU/Gi4uGixThgjKRhRX5
5rAXiezQQOliEGeLaiNhuB71O/ljsY0Wt1o0NAYTFmMnrnvzyuVKoHrKNNKZxjjVoJEUgCRw7uO1
kPmcYfGfT/Lo/7Q/pvF+th/t08u4RltDj/AGeIbwr1h3ubePzRsbXe+wL1T31LjvkaXFsq+hkscF
1Cc6KAcv81slLdx9zd2+i+Qj/jpTTQzDQZb3oNpabZQk404WdAOhgQzqpzEY/a2NM9cIR5ogMJYt
L5BpbmlfFUQqtJfRCE/htg+uuK1HlPuZ+8XcDi+YolhUYWqRV507cgLuMqzaPFIyVlOHlQ17Spdo
4d4sQmQSsj/nuG0IwRPMY8msF1laQDVXi9y3kPghHNQARyU6AGFSxJb1EnZnVP9PH1fNF9+g4L42
DPk1H9W26JTzojAvrNv7E+28iakQtvf43rBJT83OJxIR4Ela/2TyLD+lNo04WVyMulYgJ86Fktt3
AexVSCK5eAY3ZEQV+TyxAeYf93LV5mv8wB9pJEoWBIY8fTURhVZ+O2N5ChdIOBEtmlsDg6hsnt/g
doYvak9B0WVXXojnpI2ElzEYWTamAP3qTNyCrpYoyS4zDekvjR9XfBHwSZ12GSBZL24NwbtjzWHo
h4d3SMf6+6FG4FmSwu2VsJjSAoGiDZ4+I0tCMnPPXTG4n64UsQ5VCTcTgzzCIzlRxKqfJPivW1ex
hzjdjDPJia+KZA6wEYhPcymNNS7JodRSIgOhEWZcvsIrO+ynrtSxCJcq3QjMQgsyP7h5EfBdicFT
4yKb3G4oqJOjpAjy9BTVyX7fyDsgpd92PqZ9CFh9twLz4P7fpy4V9SrKFCrXCbIcCmKHckdryGny
9clN4CUIbfQ+1jPKLRscEJTxZX+fw50mao/qwpF3XtyLVAE6z5kQwk2G8dRupSRFumXgEhLGeGhg
5Wrjkez0hkRt6YvOjTs0qtozsEJgh6x/RulheOxXR9CejiN5mBfi4qFZW1MO4SufoCixd3zvzc/d
r5MrGx8aI3ZLZOj1RTPPtalTtIL3CVtN/7w+Ic8QinH3xMPyqmWfJvpeUnU+oTemgHxwgCvwHVFv
jhV3vVfFPctB8LTdymoz+ZLFxNVW9RY802iFJnLdZyEazxa1YW29rGv/nTK4qGlQeMiKJ7hBRGlL
QqvuxPRmDhUztgJiPRpQNDLMKuAGNl37qOfV5HWMNskKv+NG+29SMwo6152CWX/yz8fbMJfOAzYO
flmGwaxTyKoZHOjb7pa3SRbwOyvL6iONwYxSzp1yB4EFrEEIQwl59MiTArWQmQHNuNL6T45mkxtO
aznAMM1NOnv97MpLs3CQJ8URjdqp8xyykWUDY/drzcDyQKVRd6wsjAOX0vSCg5dg5kpLlCrxoHCm
xXsmN1JoyNT5QM7sUHVn7ppaMPg42ih0bwoiGZYOBUWEfKiIGr52h0RT78Yw+09rJuKDWrt4F+j0
ouJF7AwGHwj9XIMpXxGprcx5pGF3sATNhF5a+eoMqa18vhdol/GJLvyZBnCurvTw2reSCTfHdoAi
7AqHJggsiSPLKl0qi9hLR5sxx+wIuVDCTrkvlhZJxPtnH9pvOhDKTf1x6mDRON61RJDS+PAD08hL
nMYZrOsXgVs7GWRAjm8RbHAlMpqgjgM2QIEvIE6Syapz7Co5DyKPrUIp6pTpCVNiv6NeOtGeqQxT
EP4z5/Qr5ddondZCrhYUckbcaRivMfNixF5vYFhXo7/yU/En0Ioph/ApE7vu7XqW0NFE3vQYFNIe
G7vmJ6evS0wX56dAU5r8NqzQI0QgsR5mrniPFoCUnmMi+lELtbG6kgw2utaIem5eQVpOWeRK1sJG
Km22HIx5OnW5EcugfOorS2BAFME5WdevlJRT9T0D6rMbOiWxpdFCrN1Phlx6vgFH5iy25FTCRJdJ
oiP6tqc2lLmtJTBgA33R+6yYlP3Jj1xmPV+izqrRNEZm1blAcD6PwhiZuR4FMigHOD0s/pHOsqDY
k3+m9YyZVKeizOC9uy9D6XLf79eVBFIsSF7awStgyadQnSRJJhLMQb0bhwv8FxVrQtEWFnXm2qJb
KQ2OMo/D9r6bbHS3cqmasgMKl63EKMFrBz4mpnlJNLypThZN81gdhZRj8P0QzlcRVjR5PK6r+OxB
+vKGFP/24+Zs2aauTtF5F68nwMJkDro+gue2U/m6raBHrskPotX4OfDtT6RDksqarkVmZ/P40AN/
LKok/ghxOUoCkY8jsWj+/YLNPaSxQ6YlVQYjTbEIbd6ygY27TLVXXrWjS0rsBrrycLYNbBuv5BNT
kZYWM2YPiAiydgVgyg6kF6hdxABv3SlZKUGTAKSAp3gxicutnD7IGBJFmu7oAfKQJQZSXxJ6SLgJ
WKXUjn0pNdsRtLJDccmz2qF85FqlsKyw8pINq9OSm6RjsbBM63c3PcSej6hvZM2tuDQ1thP2XOnV
6XBzdkMVRsEHodPPrRUiYZ5MfS6zncQUwaRHqM56NCiFvvOYnJWPVGML28KE1o0hBWyxW0SyQuWF
Acqa7OSBfCGrgj21mXd5/IAF5XXt84xU6YWagIum56A+58Ro/1DX9l8ZjeoE2tJuBl69kjA4f190
Z2TqeOTsEcnTUxt6OtEydk4ycicSFkQpLgwZ/r1LczDNh86d1Vq7P2GB7wnJWEzdX4j2TwP3ms1Z
3twclyJytfbJjtHfSWy/pC/GlhZ2fMmMv5HHmKXXWPbXB82q9OJFdqIMmTZEmnrEOkKfTzmq49BZ
IpB2jeTHX4gs4AJyiQMdVkUE3N+vrj7TZ5ZN847y6yIIJY09hkHyn10RnbDcQUXhl3Hsqw6u++4k
V/UyV5t6JRAU4RqoAbUlI1tephmrBW/BhmofU+40X5nMO+oPXJHfSqY2bNwuxnvln7z1pgStjCtN
/U0p+cpwZelqA80+g7VRVEGliwoA0AYdTr3tVjT0PQt+7z5VSnCiHMHmRXRTNi4jAhvknStjfXTy
3nJOFpk4aqT+kbG6sOpQFAk1i7f9c6leXtzH9JJT3kSFxMXeHAcVH29cu59TkqZCCWeIiYA330RL
nXL8NXUrhYeS5WStITggwCdV+q6tEU4yYdfKTiN0BcDQ/oF6/9DtFqEctZwf9WkaIwsIpQB/xLmc
vk6EPSstaU7y3Zd+trhKW2IP0krOQm0W468m8vFKHq2WKfqj/xjYXgxN9A+hWGiNwdbbWaSGX4YG
lpwWh2QwV/YlFzQmT6eK/q27uAqIoY6mdfJhzbnHHS0/Jeaok/EEP1AWvyAlcrP/tpHNZ/JYrmub
rT0Kgr7a05kcOyx8p4H7JO+jqQTgriE8beKzF9H9Oez+zsGRb5LU18DmPeFquIikTxV3r+oX+8rl
uqQ3jYWGAXhNU1P7/Rm+LzMK08R8NNyDvtdEbySgsTqrEeHykJKx33IiAyCRd/agh0LS6SuaEcgl
HetFPZ4Z4erdg2Uc3mAyyQG7BHcZ/GyzdXjVbtQwD40+t2b0se3U+TFoqawwS+zS7yqkQ2FMX8ru
Oy4VSJhiUhTMw+34tzkYZh72LgHcXS/Ha+ACBkb1bw2U6mXIZb5amMZluBgU2485AmtrHqwRyGhh
uFOKCHl8gTEESbc9XOlzzt03aF+zwzt5+Bbsg9vZg+C4qBC4aokihKHeDF0qeGMtMBQgv61gWkbY
rMd9PqFe9apbYl7lMYoCevADAFmtEas5SsmzkHCFsKsRMZarMrQjHbWHmVKqpzg6tFoDnu/vH757
N84uJ6weR+kiYR254NJ2xzHNPxPzSC9oqTkpheW4jfjeX+d7hQaXtPw81E0TRLMUaVxeB0bZsKZs
haQ/a/WgNyx7rjhjwpNi8zkSjLOyDKzq+9Wmq3tfiHFL0XwzqmjdA4aU30c+RIUre/IZiDOlTdqS
q2PwC6+wO54Q8mt5lMvg+wFErDSSg37YK8fp3zgtbPLNOybc9wAyQ2kJBmxnigC7G+7g4jWwsXev
60PXM2iaLct2DBzBGVdIEMTGswC/Kdip1NUv3Jg897zRZTy3mndNP5RL979EOCIRrXJtywDOPiTy
FcK9i5FJ2X00J/4V8aP43tAqFWnqmsNemLn131yQki/+gnkPJpfYLZGzZZqV2hNh+CnSA7eSpEcH
2uch2OiVW3wI+qaL9s//REC/KI8G3Qw1q087yXQm7p5c4MXTBk6MLhSBWle6YeFjPV+vmUwN0HTK
XTtLPIPSMZIS5xprLE2MrCEfH2QfdCfRob4v7M99eRpMuXFEcJdWAk7YAccBei2/tfOVI5janC7U
O0NMVQvL2rmd24O4lpsrIO7DML9UVezSDCh0r4Mv+hR0we7QQp19wRbI8IEvE6fDNuQqhK8/lPhy
s8MIQtRJ9BduDwrPw4gRaz0tCI7S60vfM+w9z2VXs1Zu2j/fyZmjzJj+6ccEYs+8zDiv+O1luxig
MDoM2huMxtEYNhhqBPwkYaz+az1alWwFbiSl4xHJl+u2o/hzweiiofM0BW391QM+Z3oqwUrz7Wfu
hY24Th1wPxPQ9V9HcjAkzJGYpKSmRJZ8FMKcNeeNW6TyngBJWktKKsbUiKOtrzjlmd93q1Hr6KFm
Ju9wT9h2xot5SLZMxdq0oEiJ5UWYEDio2Akzl6SBh6rOPLAGjZo/cAac/lrhyHS7UABWBQzXNpPo
3zvSAd+9Fjyc/H+dqE2mywDqqLACKuSn3QaLmXDnwlw9cOhwqWneFeOXLVjeTZS4K5Mk4I4+KW54
WxmJe7amqiP5AYipbHmigHQ4OpAer5+N9GT1U6fOnuzhfNIN3K7MX0oFinlvlGVy/Ial0HUwz6Pj
L/zl0+xzE2M7leurxa5z8uhp0Ns1XzERjDV+g05EAJQHhs4hsjwcC5j9+7eMVPx/05NHIJh/9fkw
K8HvbOVBEKdKAlzHZoNHlwLHDlBg99BL643kKRciVMo+nilMuUzg5Bm8zYmj0MV/tByg7wJJ3cAz
a21wJIr5RVx3QkgvCoAtK5wn7BwdSBNKp6LlpY0+mL0qdwMDq0/LvaL3J+8gPJtgOwZxNlW61gvK
lVJsbt2geq8nU/lKA954vJnaTg41SYfp9rM8gj3WXt9tiLPHjbTjr0Y+BnVA0BVWBStiRkTLDRoz
5YXnxdkhBxmbrqx7O3nuUWpRuLpEJ0SrJDTa/hqWzEzKVux0GuX4ko84CuMlfUAjrhhTpDZN8tT8
JdYhb1D9auk4D9AqXQZzR0+Qnod2NbOggUFM/cp/LHR0aIBB49fIb+Xj9OKa5UgZXpuUndBoYAC9
2lBFockYAue6MJ9Sy822tChr1/Qxm6qheeNnbEkO5gHZNYxC6Hn9Yz5MP55NSlqyfdoRH7KCrRG2
yfZYFYTA3AEaJEydgOlV4GeETIWaHXiRgv9HLfpXBXb/658xb+rplPOMtvTn+4xcBILUX/SJ/lz0
/pEHvqdEh0TGLVFI8N8ReOI2r+M7/Rr8+RLHgXljTSqSVBMgyJ9wxZ7WOB2KnXG8Wm0Luj5pwwYu
pxPmQ2zE068UD7/R3gvcvxtttO1IH0ioHxZwZpHTfkkWY1wgaeNSGHn6IF43oSDWVoxfNjJ7OwAA
VNdbpuJCnigNqZ3SZQXPZ8U7ftZ5nXnqhPkziNNII82DsW8b4qybuXzQyEykEMa6sfh37Z9ST+HG
INzUsmQhIk7/usLOmBgIfmQRHcy4GVnivtpENrY5BptWftvX1h9rwMGpeDYJbDzJrPad8dL4Zw6t
iePpDu/mqFeZtdghUhfeQK0BQzSepmsqTxuTNuL+di1kXm55nVfM27ljsaJj9rqzfW9MNHl2ASRJ
VA5K7joyotVhi07LxVg70ac8+ow9m1h15Pfg9LbYrRpKhcuC6TdFtgCe3NJCfC83dEObuYtjbrx8
8NkDarHoKg5h1qksZFohV7qjYEYrxZh4RPduaua6ph3zO6Xe2CqEcsf61Rxgg+OY9pb4cT0JLtMo
65k3LktC/Axd6MaG+UI6d0u85K9adbClcQVgz8boYvHL4CngICfAFEPhkMc2tYYn2As7YdCxfNeB
ujtiX2nq9JEts/k8kBaXmS2BTxV9AnnK0sWNEduMdKbpiZIiuUghov9dYNPnx60V96NqpdnRvJ7s
+N+UCbKIin6h+5IT4/POxSP3lOcnTKo3+xl1Yizc4oF5jRQEjt5SVyGwMCJTDHFxpLY0yXZfhSDN
/UOwGQlNvseko0Z8PXxnlG+O3IkwesSAPgGyAHgtaGipj/DF4R83GoXmTmN3E7w9GlKByoXlhWS1
MxhrcV+hIv3tPvXnoLKK7YIht9BbdKufcZGa7w7WdR8W/W1UIzFtelglxNIqdupzXmUhpF64808V
WVSMIBrfUwEfW+i72r1qBr0qQMIWD9YbSL4tKXkdDlgSOy5GStnNXfpZr26uS0GoyZCzTWZLmVLX
oDzwwXQupa+t5Rwubs688XSIq3VaPgK7pt1SR8F44OWb27BX0tk1nPzaEP8xw3qiGJ9flgFWETqm
5x8LTcxufKEe2keOpSgwnqHlPpNfQ7cRzVq3kp0QgvzyIuFl+bp2kaNXG1/aadJ/PzpOVaFLuRvN
lcbQMJiCdA0XtjijbJXoRup4DrIb+Xzo+MBFT/0kDNYBnP0+3TA2ZJTgWyiMk2TNX8QG/35ADcqW
IZgvjZRbWo3it7+TzOpgWu9FWsfxBdEtBoJvs/wuEY+h9sXgUr4DR4h/C6FXmqVgDaVLVfYkf9cd
OUH1M0qJlIXaZ4DJpDlndOX39o+75FCESsUxyfPGxSCG1ymSOjOaf/ug/aVJXXHI6pb/iGiSQdWh
7b6QKbvrJIUUJG/+/mtDNi3oSYmeeMS11W3pVAipI9QkcGiMPowaQ6SPdu2hd4AZMPqoBbmTr8gr
sk/dMUWzkukdBo3pIz6f4Kb5Vy9qCeNCoBggX6+1dDJa6t7Nfg5+InsXkrTBaLf0bHpWwL0PptEa
/HvZ6oLJBYTKlJ7w4Mn73Gx0DpU7Xw/phiMdK5NuoGyYiHqG2uP0KQ5gcCb4IO1qTEZC1HjJGMu1
lnNRCiX9SAYDndq8UGjMzOzIpjgKgR8uoj/EOO1S8L54TQDYc+/KraA3Z+Gqo3+wMU9X2mJRp4zm
qBuOLs6/8yW/jdUq/XreVaCrqJe+wn1wj1XwPkdrLshu75CKgKzbCKrTf+0Kk9qNG20daAyq+N38
1Q+338c1vkhZFio1NDNQjEfZtvt115h0VCxXcn+KF3wyZYYpdYsxW7KHQm92eoPruAfGUCpdixan
ZXemVWrrwtyzwnVcTPy8HbsWA3cZ3MFlbchb99MvLxUp2GUnHJom7B//xaQ+i/YRfkJoYgzlc7YQ
eK5jKp2tXFm5szdQok1dQLQ4LIeaBid83apa4RxeTwoHeL+LFAlaxoKXZMUSFHbixnqL36QZ1H5j
Gs6DTcBDHWcc/PtelXYxk0rbLReC/HW+FwqZ8HiEuhStV65shYKjvnAu17/Vw8Hbv+jwU2ZGzGp8
UTEZ8r1T33lvxVfzIX7b4s++biGMmEsm3lf3pemylxvZ25He+AYelO+IEZZ4Us9Qhm0fAorOlZ1J
AFq69ogq5K9e6ZJxQswESKHNI82HE+2N+QM7dl6iCBpEvNgdo7dXlo+tu4aIcWxYdQDtZ3IOiva+
LZ2dI17Jle0IYNEEhEhLoXpF/YwlDdHjpq2lc7/dnUy5Pk0a9vWF5vHm1e49qMYcfXxo0mdZjzf2
/+hjWSBi/3V04OOtcP32+Jiz360attBcNCPveQ2UgghZulSg6XQLdifjlUlnU/0eUg8GhPn+xs96
N3oYT1Cnl767dLrwKrs6oN1Z5AhhnK4+WdpqlgwCsQjeGXRgnQQTBUHg2HBeeOK12RpK80WPUY1g
tGDCEx2IZbBU9E/gLqOGXdr6KdNvrmrbNNr62QpBGXM/ixW55lbYBL43IK3En6op0HQqvkG+2A7I
uwW7awFVgvHhXwy1A8Ub9pgIMJ00vuboNiaxpWp4nCbl3kFWBmtKmxjODrNdL2O19LCOqgI8yhWZ
Wq4+e8ObXPLTFGoLHfWOmUE2Rt1PcP/dcY4zyTudID/udCFqTpWAmybaOcRf8+RkWg9zS8SjbQjZ
QhedJfzVwExbhHQgJuR8QHVvv44mpbVl8WzTw1kOKAm4sZXgYDtzwDVQfx4eo9D7NIK911IG7GGF
M1nVeffcjJKJvuVHZZ9KBmSWb1TwiOmp3w22AwwiR09f2vLM7t3YOxhxPB+7CHWk5cCQt3RhYcEv
PMP+n6eYqi5ypRN5/veGvLfzZIO/DuLa1diPbukaS6MB6P+w+LOwz9t0LffYqewRa8gMvvLaikng
JEjpb8YPIDhfOrHlBIZUp5CVtYrQJdD5m0rOWm8dT2rK39d4a2FWe/f5JvrVVew1Rrx2nwEs3tLN
QfISJBaNJKC+WDinNPEFj9epgQAv7lK7wiwzBjg1DtJ5ssSYt0HR10TezDme1eT9V5l5zbFNcyn/
brq2HLoHWqJduJakD3jv674QwxVjeUybX0VQcKqsr0BQv3yb1upNcZo1fZm8fPuUGpJ8q7feeoxF
kGgcpMN7KoZFwPBnkJ/R7URgvmgCnOmxZe2VprClNaYpnu1WLYNyttJCe0CTHeDS6M1Q7aQB+jTe
Ol7DW3T1iSp6eDaY5/ppIUxuuslLfV8BKOBHlGNU0WEgbR9a1oWAkZ9uNvSIJzxJo9tWw4tKxKMD
Tt8FTTLklfCJgASmWC8HAzTY0YtfDJ5sR5azziNzXgT/tWOe/sRP8zoGRgUmH9lHlY2PnfaaZg1r
vTG/S0lvT3VujQnUxyCHW+i8bVoQBA6B2zGOvvZk5BClo/sv46JMMXYpaQu5aRQUP3LYETacgNBl
YKaBsyrnTNFXrL5h80qvkn+JWTrYSJMFThzGYaHAvSroGcZuPhjds1LWB1oNtHlCFVtnupWUMtZI
yrTlekG0Z0vDGU9+Xu4BtjstPIJvvDR4J4oDv6K1RqNxmPViVJgv7Xy689HyVhev8kKr0YQK2qAU
yEMgo0zl+Dcvcwy1i+ujKfA5mX/khOQnOrzzyKrIwwIWqbnSRcGRbsolUYYGByK4V6B7OHrPgaB1
MAUTO9qYHKBgUlrEbpOe/BEt2rejij2NnQnaN0uy8b/qqtoarBK34O/nCRXBPSjOubykdOh9rygM
bw2sbhH2qabmGcBZGNWTy0iv5p1oMnNQHLJldWaHKJJznK59RARjZV4kQnFVuREQpAFsM0neycEM
r2R6I6OSCIbczUIkULTeh0zCzMvKzkjjFEzSL5Z+4sbHjUiEVwhrWV9Njjq1yu4rbF30L+KM50nc
oyTSJZD871TZOiEnC13OYzYWHovOpVeUuB2Skincra7VnYNH03q/jOgrCh4GtCo5fsJGSY45OavL
mhw4soIYH+eEghyKDmIIMegtfpZxLSS8Rx/mxNGlEy3mjkR+c56/zHHBpESrs7UX1pEYaNs1tt4u
m3nvj42BtuZV/ZYCI91n7dqbl5YO/dEwg4PGwQs85IfWog8eIxsNFRqy/qT6GzA1etYrr6A21HlE
zxeJbhCyoq2Qh/teL19npiWF1bz+8dve/R1C3MGybngy+09gHAQjPR1HjxHmvuKMrN78ypdglOtC
L0N0T1tW202b7/AA0nsnJ4SQBygNDy/XvA9kYCixUvZ8SiajumTtpRTzmkexBlBwzQtbJTfMYI2S
CTuxz+26kvijANpeeKr4bpNGfcRXtpqZ1aC8ra/sb5s3yfZfuco1C6OJgPM8mhvWUQyQ+Zl1mqIw
dD+894XX7yPShoA+9PRoEulGTTN8Exf5KTuvSsu2/jmHeHbHJxsUNngwIcKi6eDWCtmD+k5C1Gbo
bCURdoqFV+kjIzORFgj5niPm9S/FeZCEqSF0pMn+ficZx8QBqu+JJABrmX9ygla5eN3VrHTAUwdg
nW4YYsKWJ6HaCYjnnbEtHnapmjpkdoiRqOqZNpvwUXs52MiWLmNF+wg7O7XIqheUawj5xng+itSP
UtTIN+qz9er1G4zDxcB+tYJ98CgHrgfqN0F2vOuku28h2e3iyJLrHCmUX8H8ckvmxkZbILa0z1sx
p0II8RKmqQJIX++bDBHY6vkZMFZNpx0e73rXuDcqfXibyg2XvZoyc9OFSEMmnbwZr3RcxWzULeSi
RMGbM4Ia+CTjpD+VLSiEQJmEPyPBrQxhSgDY76d1hou+PaWUr1Vo5+y4+j5OwYatWcnjeQrFxD7u
ROchrvy2VAVlUlFLmORn1kBbVBJ0CrHGA43BB0RqnKHJPaAYJiz3IhHLMNVsC2blDDLJcsAoFRpF
Euysb46DGYTpLt5wVSCAjlwD54ozdvjBXFwb9+sHnNPD/dKi4vn6lzspEh3yrELDDu7WEMhUn6NA
8n/MxlY43U60uifxVSdgKNOYpNuN+hYtGOtDrAt+Y8e7wjvfcPOVf51FHZ6lnMOzk4JO8Simb7ts
rQ4ya5rAQwEIWrqSiEOkXFhGsBgtDqsVWdG1qw0Q8UlWWBkMcZwvQdcdAqXQzMChYIpC3PQ5a6c/
IVVzOFylepW+jG79vVfaUH1YJh8i6rV5/9sj4Hs+IlTeIinX8zaLmNgq4Xi/SsZxnvqpbZP6mRYD
oQE3Y1YDX0w56q633LyMBEHKfkvDZfoKJNJ6YJV/VYELAJ7goCc15Vld4uVDVkls7uV6VbbRcQtZ
39DfnOmSL9UOVlxOoy3LfWJfQoPOmcDv7Mdw53Kh2edIK0L0lp2ZnjsNCkhNjhfmXvX47F26B5Rp
+F7pPqFsVGNNtdXHdYAVabcR3IWm/DiYJGg/TmNDp/Fs4RyqZFY7k7b3Cf/Bd+cZkE4FggoC3GAF
hBLzW7ZmifNCmk1v/PUNjwrg4q1UKBIwAjbun2auNF8MinxGZnVHYHefO3vN5GNseUyBScZ2SXT2
6ptg75SmpQL+sc4WmakBYaHoRUz9WUMiQe+H9AolL5wh86D5yaw8oTNN/N/XMDs46uQOXYrM8Jnd
WMAcPjscSr6Q2LngeGs4nyEB07/j1rM1tTs/Y0yKbrcuAOScF8D3RIL/Iz/+qw+3L+/JQlZl7ScZ
MjXh4ykRLW5GkrFYLhLjM0cJbyTSTNgmU/q45hPPo8ABRdIZrATcdO1M8KQKcxh0NQ4t7wPBSf9t
+DelljaZVV75UmFWQAMsDZHHsv9JNT23uNTGh8hR1LGZbEmKPC1HngDZYd0EEl2Stx7U0cn9hLBY
PFg23wK5GdQWW85zj2zTktkowb/g22HC/mnu17cctN8qEFaw6xiD6OeUe7Fvp7MQEW6VSHvPLY5+
9HrJ0VYIm6c+wOUfLWTyFY46iZCBSIujPxi3fIoQCkXAx5QUQFfywujRDiH4zk+KM7kI2MbZycLk
gH24ar1JD3jAn4/fShLTaeDBLYRWxDfwVEFBnVhQXBe4EP+tchBLmbsiyIKmNgP8WvNOiWxFWufv
uPTQh7QKcr7ebG9F2SdFDuoORw+9981uKqa+hCJgc15y/8tuM+yHhfbQBCzlaV1H9QVbML3lTPbo
0Jl8ZxwV9OxCtdHToKXP8h58pOIplrMOjGDJBdglFm0pKFmo1DIBhTuPyTlgAB5ph+Hl1bJrGQR9
0JN7e51hym6FBRp+9PcLn1USO3E6D2ZNfeQMG1n2cVQkstx3faoF5QStx0HeUBxYQfnbYpGgNo43
YRayx5us18Ry6Tc+viYwa5OqjXd0dJ3IKG7+BSocuEE6h+9PrcYEPhZiBTfbIm7sH0ugvhtGIwCr
UPbUzLW8RTYizEmGcVeWU9blU63D3P+vAC1C24UHE+KdwkoaZTI2hhPnF0XKOlUrrWqcGlzzwPL5
tS/5Nc6IanXQMEEJVda1GNqdhS+6ZuUTPVzWfEtFb7JOmoWshulnaopD6X6k4XfrIqEYHRqgv3Ce
GHXv8NjaWd/wQM5byiExF2n81uNslD/O1KItoFbreCWMPjVrVB7fecVWTyshHwUztJ9aMZ1Tq3G9
/2W14DeCAOM6ouOegklh7j+cixj3Xki1cChdV6Vm5Yl4odlpPxF5Up6NqQFdhdJ0KpHHGtDiPrEy
Vnq35B0XqF4egSQtaDvs9s5I6R5Df1OaXCrclXehVQdO4KHbg/DaJNi7k9xQs+qretXrraa67DTm
FLKxt3TGEsfxpcLLHe/+xhdwilfT7C4ahYLFgZhi+xfsqFp4c6qOZS3n6YEBMD9OxrfwbTt937Nq
9IxVRoyoaM7Sk5EtLdbWh/q2KqEZ1kqO9jbM/i2VtNiJSl5OLVRkFSmioZIifPpD+yjeDNXne9km
OnWXiQw+XTN+FzxQxEW5WOzdyNVPUjeZ5YeP+uBl/keNviYwq6HKVI8osevL4Q4IP6yB65WKNNn0
keI2GgtySgsv+7+J+uB4Lf4OO5IEpGNwYJPWqG0Fu/7ZN7SA/H5IROKGN2Yi7DUtQt/exo5bvglT
KAPjPeURw5irI6xcH3LL3rrfzIwyXZPFvKCSe5jRPexLL3qCBaLzcb+aThmZRHBHqqZyWQYPzwPT
vy1OawBkBhz5diLpjXnQUbHsghcNXiI7ep68EY3mt0WSDXMyuUqEURr3fGqTmu5iZNZAc6qy6C5f
06vyA0IkvCqY2ohhYde9K6qMaAM97U7vlhowcmAxnHkpKGh8GfMPN5PfVEB4fwLIge471HQJlSqI
jXBU27eUkhg6gVfCK46nBHQI6wQpGrb4SSiStOpANdbXoM/Mm3rWIEpwf0R5Dpxk0llSSDJu9vu8
ABdSxHzIc3Ck3pylAq2wbG8t0mJQKaW9gQeATC10DgZ3CCHDSHKMrM1o56g4uAFPC9/XpAo77ez6
WNUGFbHaV3ZesRQjuBtifG4T5sr5tm8jvXAhU8Z3q/TSmaJVJTXVoJfKIeejCdZ/4vv/+f3W3VyR
qk16iMvjCpDIh7PQ6y7rtjOmPZtmSe5sKC42AFip9gcKuW5/Svco6tKjcDR8C+9lOsORS5D0/BlT
sMEeGEdaba7EO7Xl86mPXQ62rm25kOdDip6XMlALOIdnEOjXpXjo3HFDCypxmNjiDyN46T/QDSDY
xyuEaYMuq1XZpnmE2eMW4Tdi0pKv0dOdSzH25DG3HGJleOHenS2kR7Pw1gNkxkhIFnfg7YDZ2vpS
cECfa1cxm1cx5cKJuzkaffys/cEZXAlA6SlHuVTFMhBWl2nqxjuct9KJWz5bdaXtCVJMbhMZwZLa
E2nhrNRBY0l949KVbcpdnAfhg6ScFdnDwVcRdi4abpc3HCSCj+9wK6sonKrE9OLcdMNI5E0BbLN/
JyoYJY8wdegqEuZfG8hS5GBDCn1iv5vzCp52cnS5DRSDrc7FGc0tbZLze/wdT3SCaHlwioIHoQp0
OCNLok9nL7HXvMyaGKQQY6UOOUiAZN0iad203NVAruOlmik31hGwLgCsEB0Yq16S7zdmeXwzYp1M
a7mhOaPFhWK8AmCRxnP3Bct+gDrVDwIxYn18qGrtwZLkZcz/sufDEwkygGkkC+mIg0Jy1laeZKbT
njWjp5DEKhjq7pbeTqS6H5SBjNTG29/3HkhYKISWb7abOFm6X+4p9cd+b9yvOx2ux9KUcIBmYWpR
48a2N+pFU27/myKFq+ememIzLMmnjREoFLhD68lQpe2xvIqHnOCmqDtESzafuv3DFsUSu2Ve1m08
Yq85yuiKO/9Wtk08+2SimpfgqorIpsCV+70Zl5mjPo+oA6MVB3pCqCErO0+n9VHvsfw4yO5IJk6D
cakJaQI7vSRbBQIU6SaQ4Qo9lh3e5xl/1XpqiAacVnEi0htOpHsk/e0AFE8pw/OH9mKZ28vG8am5
8wECBwfBuzKWo7EyyJ2oRnIQzL3hT/Ju29aBGylvadi46Lo2WxDVAB9mjHAWWwE+KoTC0uc012Fv
eB2KHuzXf7ZSxI63/MZ4LVMYcQVBuuVbBfFvSIdiBM24adgilW25BEjtzGpvekBRUJccA1Ao2p9X
hn3ckJEbALmJsxfKUJK0M8I7udOpQ/KcpCo9jrEFuc329YfrlhlR+cHyGJP458PPucL+kaOWQCCo
0QnAA1UUu19YsQgwgoDnuhahTc2/DJnY2Rg2U74s2seJm1bnbycA4y4sWWWlPXWNunVWRc3GLkr8
IC3E1q8CQrEw8Rfvmlmz0MU20q0I48KOO3NCYdGTUW6r3lgWAT0+PunIyqmNTewy5/w+5KAuY03s
7uETSsRwwq0zPV3fNljTh9Az2QSumfZuTvq6UyBqwarJ1/xMD+psOviCM2vHPEDpxyBTSRhZ9DTj
8qu8DbUxY79QKGeRnJj/XSX+DMAYKzhRONPEFg6RuQYU88ozI35DEUsffcJXZm/e68cde1VQNDsu
Kr/SaIaqv2altOW/ijkNyb8uU2yu0LE0knsp7Wq+IxE2uErfhIeye7Z5gqgWF+LC7BZeFY5zggYh
g7ST3oMt1hRHTtLtowjXLnQ2PsTFuBn6jBEoRXVtLG3pPg/prGF1cYLtb12r/ok2D8mUw8kXyAqo
lCg5FDI0xBIKHBcrAkQrag0N41dy7YeOsY2TtzvfwqzYBzPOuGrfCRNjHmXHVtBBskhTGhhFcNKU
Ia4rIB2PYtZJ4meVhxsdTzSa1VBOs1oduMTy8FYn9ZOIPeUpAGvnv6l6OOtJzNnLWdT//ypOuybb
1rQMIkjLCNlUGMosyvpqEpmkvCIsQiIxjsaXWZkPzwmW8i4OWHcUuVvnKBEnV5/nyCTX9gCVrr22
JTiPnvKlmpOpMekvmvfK9k9kTwoy2107+YpVHKyUKakMQqrK3xvzakENgwENWgVnmVbjafV+qYbh
BzVtAP4CQN3bdsF6BrLbVW0hNa70aTtjjvYzENBJHqWOURF2kmbDp6f3ukPH5/10jlT4WSVptekf
P2ZDhMVKvzICJ+d4X3HipVkTn+PpLilZKR/8e2RLIVlDpvnKzBgvakO/Ns6405CYooFRko3xWhzk
Nbw3U5Gvft1NUMUPLms3hZ4azjrXeiw+cj3eKpmhOZeZIRCEeOFPJ5DTxeRW59GYFd3o2lpcvvwS
ujU9fcHrILkQtjXiBpAvHvUUkq8WvR/UVvi8Rl0RblL2JF3by8YMij8XN7w+3Mv0ZUEzylQZ/Hf0
XJdz/KFHmTroKxQwiUew0HMYm70pfPPTPqz7XUsncz2+n2p1T2DFXptAxen75zKa6+aKP0keH2Y0
OhiIfRgA5ojo/2hlLJgKnC2ZodTc29zRX8YsXY5XF8zwfw+UihxdSHygyjTtENtIUzS8wWfbM3vL
cYPT9F48mwvfp6blr2RLxL0zxLcdri6SrtVVexdLBtXPJ0wtsP3i0R+sVUKGBqZvz80HRVHN8IB0
SilXX07JcfCs+QFqfJVzcodZiAEgQuQHIveSGYue3kpr/MIvwf3ISmFUFkvExIEH2P1t3pcJy+0b
huOPM4IzYmaPk5nTi/GLM60bhHRyi7C7djzx6lJucnK72K6gpk4O5fhfzrTr1AO6YDotVJfa2BpO
VcztIZaqenQDHsXgOg9P6QJ7bWFBi6IFl7H6fWsgLljji2hMgM8XBaPPV/r9ZE7d3RsZZwmixOQf
qNlAqGc+zT+q4TS9OQDw+1AqMRCsTBCpYwOl9HxWWe6U6zWHQG92Oo+WXJ5+L+95FNhUwxL8kGf/
MTtvvPA4sDzVxqP7IFth38fw6b5ADQxjclye7XTCfPapA5Y0LmMn+WiktMLsvw8z2Pcwir5q6hwO
mnWx4dMVRk3XRHD+n3sWRJRhigSTdCDGAuTDNK59qPMzhKnXgBxOmtGKXDlhl+lJxLyyEoXFC8zP
4J2jXQLrpQwcO6gR+ISdv5NH5MFautgLga/fjWZFhtBJ6rrAUBRrQHesuUPC89Ibyhl1m0oulthN
Z49OiOprqa6oHaaX6ZnEsfMoS7RV5+ZRkpEZRSGNs7c1QO6c6VW2C+5pwh2puGmiH+FZzLxoUY0c
YNzMVwka7RFqokUf/2Z3ozb0xixA3nzWV6quXFzu/ocdUHoFPym5Bsb1A7mCz/xDl5izIQGmWNxm
oRgOkfAcwcJ7R40A/5+FzbqfGdBOxk+gZHnSAlXJQNT6BkZJ8Gsgu7YFm4jOD0wOUj/kz1I4s+ij
nCnHUyby8bDdbk4FjRa42X0y7RMOA3QoK68CEY2S3uu8wymRb+dBhYvaGPwvO3Pek/OxagfHEuvq
Bopx2H7D+hT2Zs+p9El7yVxyGJ90P2SIU9/ah1A77vvGpOJj3NEUL9BVbA/5bbRJykkIF9ZMCOtn
RBleOgqsdZJsauLedfdZUU0+4GV1l5dPbDaEk+ra+9f6c91/GOWt2VkfMujG3Fd4qym2NgLnZGxe
LMijxz7Oy12Zi5n2zH6FWh0WA4L8gdJLkQ74VrXud1bchm2mkPWBY38yQFvychBWrscDzZlRkDoe
fpAN9me7kvqudP1bYcUDSs+bW++XsNmh3FNl80Vr6MPhTtxaWQSVZvE8KcvpMQPHbUm81RRjmSOB
5RxiaLTlWZQWYWCeIrhZa/yPjh8J9OgJUAGnmleQXge/XR06DTg0QMXShwXcCocCrQvAPUsrl0t+
eil301ImQoYWLuKRdrNo7KvHlDe1VO27w0LId7hmwdm+77vsjgWM06FWlT30L74oUVW8/E9IWKdP
PNZ1sFmYrHl90RwM3D4Vuoq5sAmEcboqSBpaVRVFJdON1D4ouRWSu0dXzuDz5JknSIiMzSl8qQG4
rhHmWUHmmZDuR8FD0yOtK766bEWKD+5IsFWhjfrPIUZBF14K6HRiaZYJacYNwRZS/lvonTN1axkn
na+aCulOwvr9/j7zLTG1k6d6iCPi87cjkrv2jtZ42UaGuvnW0BEPGvyHIXRKWMPmu7vD6zrDq8bJ
hBxFA75euKSkKv5jE6T4MM+9ehCvWfoxqZoWXDXXm1Qqe0iafx8XImPFf7LcAPOu/9RW7FCR8MjE
j78pBGQj6cgSbm/QiWoCo4HBPzJsJQEwMlTkCQNdsJBxKsqhcokmcbsvIWH0kxOgF21k7SwNC90J
79WDSoBoYxveIKrpID//qttlhOiSR77PpqYVBdOBigGzj7L6WQfkBX1b0vb7ZW1mSSmspc5zODax
/alx/Kxs+TKxtimCtPNWDFd5bjIdMQ0cqg9amPCcCoiESMRsqzxA6iwg9a4Ba1fLuFogUMmxz8l3
W3pxK6q8WsS+TaxnPZTaqOCHuAXE8PxhPBFdMFNz0sZQf9HQGKgHS+qpHIgbBcfUneQisWPSarYa
aYrXUm1s3oYneRy1R+RD/MwYhN0AuRUFNWQ7jb2FzQL/JirGGOmA0t+MDs7tLM5O/N9QOSq2fkwV
Xe48WKQuACAd3y/dNcgPMe8GtQu2Iaeg6Es0l8Rs+58fONtRA/Po2SZ64hqNcEQ9Qxybhwppg76Z
zCZhHSgFLgsTFM97ckyD+yoKOaPB29CeumyOG8oJKtXTlCs2BzDdlpb2XWHTtuqnon6lHUYUndg/
Qet184r95K5+yhwTUreEQ1ElBgWMDYdnp2CL3JxyAqEmyfUC1SOyPdyl9N6iSVzoSu6os3QrLlQ3
xoFbyJdSXd4Q/54Z+7+95tltcO5+dbfi/AfbVD+5YrsDvoGacOu7mPvTmjMeUWoVZ/wHSCU2oLCX
FBCoiHviaRyMal80okcOxlwL1pLHg7jNquRGN5O267TMrTu2hYYvUVe7rXx9GyxYYWoF+7mdCEOS
tXdUzCA92l76EynUEZ++93vjlN8vfUkWNvW+heR7VhjrmORyUlbsrJkOYuNyI+gFDoBKK1WWKnBb
D1brHsBARYaXlUKfrsEabWPcr/RuA8X1DtCQo94c8121eKXqFJBmwlWQTZASEYTGW6W3GmPQmHk/
Tk6Q3Md+zIpzjjI9dlXfy3mkNmyvU//Nx4su417Pkz2slZoC5W/1e1JypGgnkVfRemxAxyjkg4+H
JyfxkcRgTNKocXeVoVRpit65E7JtnQfyBjfXCp8d9MDeTHalh9sYs014su+W1ATO8Yt5N0dNFMUD
5JbZVTO1/ZB/nXJ5Cr2j399FAMF377rPzS3OeFOS+MBY7Nah9yEyTaQm9NdUVBGg32wzVCnvFLLg
rhiDeC8EZwcen1Y1XPMxfZEJ0c4l7lXPTH1RRVc7POWh3VhkS4mXs7gCSjc3Pq7uwrj5GvTkz0vY
65xBZPQmjjgmSq9a13BTluKq/SKkZ9Q/hIn0LViXfyeQVgTFw0+ngjHJcO2T9bpECAg6XNw2sC8d
kVj8Ri9RC72ISzwYIgVdq2dpJk8QFKrJo8fBGp8USzVZwOgLOsqJ0Ek2jmeWRocmsyqsngAM7oCU
fZT5amuCZLCS0IdDYdUeopw1HJl0EDY6WCP+1kU5PtQkQLKqWeE5ufX5CQ0wcyKVuHMa6c4MlExu
eKcN+osjlIqIiKvevBRAMoPmBemqZW9oWOZAFVa0P/1w4viPlxVlGpNFK/UDRaBr+iCJ2Yxjmc4i
yz4OjwMvFY0MK2HzovXGVzWtIR9Fm3ZhROB9IExzogyIzHPoG7hr5UzobsjucU1ZkTKmX7J+yTq9
Gz3yarkAutOWR0jkcm4ThtthTKeP5n4QVsvSSH+c1DweK1actdV3NLubOiARaoRnbIvjS14+aeTP
hlov6UOoDmQuEUQ2brGEMThsuJUVo24NLdHjU125h55M9nULClqPyuVKW86vBmjPYqqLiB5DmiWs
wYAPCqG37ScmJQfMt5cndd/ZV82IrdUWaTBXjDyb1YYcOup+Z5KJ9DHSpmdqh1owcmE/idpxsdTf
flbx6UFROR/j5tDfSf65tuCvtKDF/p0uXlI089sKDciAh9MDoaZOz/syEqAe3NUhvUT4bRGtuAZb
N2OnpIQr8FHlIOotqBncbm4oalMte/dEuP41M5XlymnzMHkWFepDmuAWf0GQSzzGf8K1NUPRwxLJ
J+oNZFkColM/jDJ7jQqef47jXA6p5PMM1qjhGkNRoyA4QqrI9DugyBR03meJomn1dGLbMFCXBsFO
Z0c1XtQGCDLEOFwl6IYHqyDCGZL9R+XjMuGIjIjwlDSAA8gGaaezQu+oBi4ukKSDLt2xrISWv0js
tX+rNiWi0WLaHpPgRlxtV2aimBLjjjbnmJCZ+XWrK0JF0QVgAubUEWk25RkU640Art/3QAtIEfzw
ctK1zKRh/xn4rs25YIZ3PJ9EegIb5wPcGEKM01PEz0foHPvE1usN7eRfwqZOfH0UhNRIUHj4CSRz
4cBBnalV9265t/uJB606tKZDhdmqU0QfhG+v207gz6eC96xRJmx06WGYdqH/LKXBV13tOhqMJMYp
A+15z3heaZX/wzaoKHCOyvkxgO6yZHdflBK2AqxLxiEOn94YMIfRbdHtdYTHUJMk1hgDxAxmP33t
peruaVNyJ1mKI7Vvo8cqb45oe5fnRrdahVpXqbmpEuWalGSrDAjxcV0SIg8Dxp+dZGOK1fPs0L3s
a0wAJ3pERPIX+N3E0Z/PK9zRJ6peHN293FtxJ4vfyCwWLTW2TQQnVUNneZ9uv2vxkKoYKJgAc0OU
Z6GDf07cg6ey8varvUiZXG8F6NcO5AP+3FCb1gy/FtSNFz9womoIO6xsU/xB1f4zVKwCT4IzHosO
P0yRlksnYs1quUj8yWALRqlSvc4ZgHBwRV2iE+ZBxlzzyndr6inWcndo8j+Y5PS+3cYvH1YV9XdN
oMZPsC+AXwT7X78iYo3OQusbCXPaI05BNrZnqfm7kYmjieJ8k2QymDY68Fn16RSj/esfzqjsq518
06v2tIM/uxZ0BH6oPfTCBaPvJRgkmrGbXhIdUfoCMRxmyz3mxCKcfo/KyrZ4ywAtudI+5hcawGew
9e26WURVV4HzVlZb7Xep77j5kCAwP3hCO/97hSMQiLQ6o/dHmabdMyFTYwhYS8v0JopjghVLrJlk
PKPtrq28HTb4Y2xYQo+fAaMlBbP4+EJ3f2yn6hqLB2ZsfxtOPyjfx4c+Dta9go7g9gpYbNwTELw8
pDSPuCSMgM3OfdpRrJ4/hIunCaWXwJ2iHGsSBOsu4v0LZKoxp3IFz1Fq/6XbkrqqShxJyrT+mDzt
jvSJeRhXz15sO+fKlHDXwoYHwMSqTzjSFbrxlgLfDCZbo8J2S72Ok3TSeVBcn6Z5XLdOAo3w2dn3
gpCfjH4AGsAslWSF4OFGjbr/Q2oS/uHAzEfkC2uCvsyEg98/5K4CsMFwBWFEoj0LygSe+SMHHaPh
KdCQNBaXZ8isDS5M3nZeQyy9wtucBIKZp59v6ZAJ8b3T6g5FCYmSiyJWIBo3t5hlWuZSdIxiAvLC
kbdSFv6afLlvJW76Ig4s3yNExU1rJt6ESdkZFqDbWoCsb8aS85/XmNcBVr9R6IOh68CYAwG7Zttm
WxpdnDKtTivh+nvOmEpoTC1tqFfJx3cEvR61nqjrE+AfmNV68/8zXngNf0rtx4gpCgmQforuT8xh
J0zv3DoS3NBlLPOpZ75b0saSoVlUXupGGNejA85tkLrvaBGuAVrwGgDg8TvmzJYH4mnK1ZrKxVzV
8CC/9GVDtKtcU6PVNIa8hXl+jD0sLd2djjCzRrz09Hy2oKhYMM5H/by1hZtLj5J1fyJDFFJJjsOZ
IjEKbTDB2jWDByQd2CLq9eYrmleTOvYYVsQu1uiA2uq4+jxM0K5KkYqBApXWqDSrIPjoj+HnY7xt
YLNmOfaKdRWkfK9dtPifpY0NE7Wwv5rbgqSBwGCxsjLU5QetBGwQvV0S9+aCvk2HwGo1AiZSxnS3
NKHjCp6/f8kt4sF3JIBexuHOP5bN+3/0XxLFh+y3ShPOOiRwaKOZ5poXw61nOmgOdti0/hQ1nCTW
NFzTfVnwohvucOKPG00QMuU9SYt3Ni9uPaJSVeAKR6to7U/I1pxHK6bNsaLl6ffdzKrlSBsqkNO0
eyDAVW0NTedXRR7MZMVJxcbvPkCMIxqGMogVXjw1MU1fdM4GsJNXsaGe4tpf2YLUNvz60mTTuZec
POxCgVgItgHJ03qTkKxw6jOd6fdUd93wCyrJqOXgMFynFJL80JQkLwc7dQyTmb3awlgPo48fYgib
COmYcEr/kI1yVW2jMEF+W9LtEytoAWUbkQXo2Z8DTTXHmYiavYdReYJRGYsZAGg+6YLY7ZqD9vYW
vZmOWvi3SiJZ6CpAzxLHPiIh4Fg/kYBf6/JyxO4VJgwck1rAMCnRzrOlJazM2zeC6c48zz2AttaF
tyhAr7rhsSTar77k5stJ2ktyTh2TWCPNXN9KwagEny98nLKjnIUc0OpGP7Webx4NqkVRFBket0J9
VngS/JjIKoHFWUaF5sCO11enfGU6x85yaIAvnbRseaS+ouoZqBVk8c2rTpS1ZMcgXlMF1SpH5X+S
xRajRKq7LsigrGhhMOOQuApq8wM7NolwiyTPn4kJF9qukiCWmK8gnPX6cMSTB1c4l+qmfmMkhC9C
RTxx4wKLkEhSN+/rkYwjjAkCPtRV+67swbus3NVDN2NpIV0t6S/EzoJWleJ09IjEszrVQf2QO7Bz
3o2xkg4JgkA7KD9LYHAMvtZ3ZhzbKawUyMFLD/eL3tYvQspIx4N7hb++VQnGtQRV5bAfjOZKkNni
3+WGcCqg4H2C9x5eJY7dp3NvHVacletFBcNYnPKX7msAmcwH14S4d1E2Xb++pMfhaAFK2Ru/E1r5
Z49PWqy/dCw5AD6b3WmQJQJKZTbJZOvL15gk0G+3nMs6+zGQNRtqp7XqDDkUYsLyJPkzzT5UK4HN
Y/XyyvyQHm20PyM9hMy3OLuPo88D2tfFmociSJZ1zcx7/zKjE6cA4KDtK8shgPirWRK2Udc5deWa
srkst0vsVoIaiu2NnTmS80nlZkLD/wyAqp8XS5JeLa0/+Ag/FpOc9jkF7xt2VuD+a/DWw3wkE0R4
C7fmm1k1kHRQ0IMhufmgwLIkK9xjdU8NH4sSKCFMwf5B+NCVT6xYf2ZPSXhSlEtRzfMdQN2zE30S
SxOPnsfhodI+os4nKhopQdxWpEHZ0vu+73WcK0baTiuEsgLpyOl8jsnUHvAAr+esES0yHOKU4cHz
3gIPmjIJyhyWwApJLY4ldcFTp6zlP3VgGx71hjovTWq/IcyojGpwqY6GVv25H8aTIh6dbNyxff6m
TDmdqTmpIn4RahFiY7bKp1VWeq1KtGethQuQKMX7PcfanyrmxPCgttvy7O7ZlWwmx6CY65KWE5jh
ukDDKMSDrR52NoRr0KGILY+AIRF//R4vxDaB2qMT/Bh3FnMAEkrIqyNKKUVEJo6UNL3bTwj5jOi/
5KqU84glucyUQGphcMCCcLFA66oeDm/LX1x1iruzbfUaJOyx9pv+pNR+VHQp/LO6/9/ssONYrd+7
gWN3VHCQfbjBqSE9j+PET4ebtwyR5g1ubmNACzddXnYbu8TdfXHa3YVsYd6lpteTO6txNB9P7PCT
3wCe2qgfG0zzbv09ID4WmKZz9HjuXgOp67ZK8G3uL5+O9itZTykCYv1C7A7BLpX4x0Gy3aYYRM2G
AFQnEUxvarL1SSDitzD3EObC/c3jAokTLPdyahZpAJBzKOfOqo5HzhF0rOcBHqvDYaj9yyZjhFPH
2yG6JJxJNdRAH2FSld2dKMlQsSgu7G5tOkAJqwUcNTdXgZ7XpcPzcQ7anCZiV3HxMpzDQjyAHjuh
8rZp8Q5RZxdbXUe36+RMRCib47L/xbp/DXkAlz9jybKlzEBxsPdJ02Rs2SEgOlZhwLg/XtHoWwVK
J9VmOLgN17Ozl8iklGuxcEULoF9buwQeJPv+Zh2RqGv7GXoGEaA5kJQR8tanO6SiTqaBlXnOxmBu
KPdSnV4BRHBVVqincFYq8D1Q28bXG9Kjk6A0Dm6p7XlacfLhqAfnaUaUW9lWA4YA3ef62cPnYZmR
GWWOp+qVhOplgqlmbj/1lL+opw7FVuBbtBpPoiYtEBbNY21jW+cVsANxSYejRSz+EQ1GrB8DiKdf
aejPNPgXqCcijDEkxTpoOlC1XHS0r+Vg2EaABJO4F/h8iqt5aOMm5/LF/uMNdP6u92WVNMhSkiL0
t/08xh3LN+5rgaDG5OTs+05QLmWSqTQc5vbTW25xbZLeU4od+3hIcVay9/YovHwi+1Mn/TEeWlOP
A52QYBGxt8TITXZoXB1HDKKpkTqQc0jH2nHrUjcFw+KV8QLqXYA/z2SGh6yyd9DEPAoSXEoKPweM
JA23KN1VZpaHrZMW3tASMP9njUrh3OlAW+mqkUhy42nBEaYmnDy7WzrI9ysOp0o/1u9F7P/R8aJT
EMOjb5/7B4+C5yve6FY0N7ttjpSoqj+5ISk8NX/Ppu6YibZrQvqmU7DHMisVJ4JZz3z4rwyZpwSV
tcRnKRAYp6eJyIBbeYPS3EfEXYmsMVbo+FQBSstyQp6Gi0dbROclFkbt/CQelCV7lMIbOPnkw78X
+8+EqD/54H1cL+Rihod1uAYByrFxcMTPvG+chWIOPilzAgdSm54QTsrWC9BcCf6yaWiNKDjVHYc4
+obK5iwwCyRK1EGKvPf45lYKU9dtmdPKxJsqmkWTB2UIgZv7gxyZTpIocE2Ssfxh4hdOT3QZjQR1
jZUzR2iWtCZ37X8ITyxwyCl8CBMQdi4HT3E7AvTMPlyxF5Q6nHvoctTIDR8du5fuD/cZYuL/HKnU
O2s+q7cvy1kFJMT9NwQC12WyPYY/BOPLe+haGjlcvItiq1rlS0DbOZJBJyyJ7050XZAUi4fVSfg4
KxjSh0w3ynhQ1mNRtgUXtvTfv74JXt+mWC4eNGYuh7NvrQTpQFDQp989ZIXW4eVNwsOOVBd7SX0s
mfLZJ8GqRdx4/eUMTxtqnq3OHnIt4lb88t33xdESgwoNmlb2Csk0e5Whdu7gNq43IwzyX5XkErME
pdSw8hj5KsAlZ1qgBMWy54OqjRKOi/Er2pRoZVcvhYbDmCKN13QbZadFyL7s7OFz+NIA8gCbg/0L
uDyFS6TFghoq0/kdQbFHtfGgjzjiz7rcKu3+SdtKlo1TNb7w3cAKJIjqzNt3iT7ga8CTJWdzseAq
sFzml543GwbNHrNUVDDsJ773luzWBtrTTBvOODsjYsPHUAr89ucRbZHo09yzRNsMoqLo1Vu7Om/H
RLygfCgP0xOYDNphhcsQVYT4piDdtEJQ2axgR0eZervVR7teglHJm+ax19OFqDXoSU5XqrBqarmu
0hI+scIjJBssmy41SRmU7l2S8ELSM9NKujrElpSEDIwSkeW65QDc02PrXByieXRyrI3KOL+CTnqI
qdi5fFcwgPZwUw/gwsN0JHpOBf3pu7hEzEU6Fkrhgt0jxEfLYAPWGJ3Anlmqb+fAEXLXFuna6NL7
y7FhLFjxFPud+QViXBOezbc260scAb0oxZhpmTHZO1wbMDlkDLIsqh6eU0lmoPtZAAwh1tE7CW2n
mxs3S3VKEo+qcTbRtwh3RrRZxvnZRmd2cRpzk5aE/8JoPESB5XYFV1CKbQ+xTz5X+E3Qbao1tuic
tC09dXEt3Q7sxAtOr9pP1dORhOewhUIZrWkN7XciKY6PwDnpDtfcWn29F9/B4l0qO7iRApcsBrkM
uj+1Rh3ScfC3VGNDZa/umpU/qRqnQGKoNw2WssSzQsps4mpwz2uGWan5qyopeALgF3x15bNDyj3G
w2kLF5XTrnD/gzJs1HVq2MBP0k0VU3qW5yqDW1lvIa6vLtRdHmlMTJzSIOMXcJD3SBU1eGZzI5QI
ro2jzlqIIIPl+38u46qcaFh1wVCig93RNyQIFKVaJYA1adPSuY9DCmXv8qBH77gCCiQEuaReQdsw
2WieV9JZWXXGiuPWoj+6w4TflTUGjtdFVrn9jy1t7GD9OhGfcARRwSHD7aV7uqpGlbaUO21ZzEyk
9AgcdMrELRcrOmoZcfGKUoNtPXx2UyEIfc2AaoSv2uojplAqtj0sKOwQv0KepMNKRGydgQWn49K4
80OJPn6dbz5CJP3+Vwcppc8s9Mzy/Q6zfnvBDfUzYiRCH2XgpnhhP8k8aOWk8dC/HWwSLzi6k4hc
GzcmgLIMVWXxqDiI5PWGuYxcWqR+gyxYDFYNxA+afb0yudDR7mwJPhNcMhlUYUr9ewWMQ1da10cE
gnKzqGDlT/003w4EmdWuKqkSiAMIexVLYyAtYlHdh60FU0IqF4IHNvffgkLGjJX+ltMRi9zaKej8
azzCiQJOjAxFHLAWYOK/oVxj6pIuNoNXo7ijWatADqCaZydJB0s4zyigtvcO8smXSYK7rJbMY+K0
SI9VTu/QenVhKIjc/C++yvdWv5YbtAPJo5lqf7kYLDeB3lonmCC1vhxR+6Z4u1X/ldedoRYes3DQ
mXGhiRPR4PbpV/SiJvgiDC6SQ3v6/fEQkuiB85R6xY/H75/pMqhlzoo3vH7qYpC2njqEhIINAJ0f
HGE+0eOCTt+hHFI6sra5ZCtgJkBXWW/aKbImVmXaLH6c7olIkFVPGth2W2ITGy0KXgteWnDzIe7t
LxBJSsglzrLsY8YxOrQiwJRIPmeJIfRWq9rxQyO1i08qgyEe6aTRcCXd7O5SbxS3HjXJIUNzCbRc
J0VZRrbk+qJGb7A/0F/1Iq7wl4Gkh3DiScmpLQ8e/9Dvk4yXWweBIXYr+RipfiXvRTC9j77F04BU
6OkUzaDFMBBrNWwfWv9giBl5GZVqpkffRXpHcJkocDdaDYy8GR60zL/odxRRnUfRMgg86OyL1KGq
EryCCS4aHY/fUoHuxJ0ylJ9rv6O8ewynrizq48h7gUCmFxsnXaYPFe1SjdjC8/VtyunQEhJ+OEi7
khEIKwydEUnsnPJ0C6DEYro/uLKpi8NNOYM4JfMuOrhUuE33zwbAYJ6yMIgsy1A5W7nJoyyBb2EO
Qm2lxdS4hEk376gsgStZ6/GE9Yu3tz0+VGS+WcyNDN/9q1N/h2o9A/CzcYw8e68OXv2qIjIaQgUe
VVeI5LXfNMP3+IZFcgKZa2jBGZ7Qs8z7RvPEpKL/FzxPF8uSe4aCMHhnWN5rqmazTjTgkPJhtAFk
G0lbLEDOyBwaLRBlUdKwEMHcvedmRBBPXqh4lYwoYf8daw9HAE7E2c1zrSDZvF/GjS1DLWxFNCJX
v1GLWXtgkJ/kFYqf01fFYPDR/wCI/xWjryX6tKl0xNbFYBkDULnMukBt+5QpAFYndKxkHirmgqqc
msnGynvlNIz9Fv/d8XGuuyzyAZ/Jqai9vIrS5B+XXf55boJLYFNdsIOkthlY+3H5ibBjdokpSGu1
Ng1J48/jc/aAmsNTcqd1+WDcUK3nG4ZBBmonoJJBgWD1Okuk1JXtfCcZJAybzif/QbZOw48TUw+6
f311OLpnEbMQN5I6/VJgHT9lvDsvRosVTp4sL+L1f0PhknfcWOiLe4QRZ5joWIxr0Fl4p+jcw0gz
+t7Nvs8Jy4qez9dO0hYYhf6Kzvmw/Rh/uU9pNG8Zy6/G0IDhiblkil1RwZ0pIHQjZanK/KDIBpnL
tkgMesaRzX3FIkr7TQzZ0Df1foZU7L4GT8RTKuzM8EfE+Tien2+BS7o07qhG5ThixJvTa2hU7bQm
Vi2a9vtb4VXv2wkKJepbrswFMPm+ZpvhIdaC6IT2XQpbfPLDkqnoIA3lv9+vTHLxiCCKLv5Diiq/
zLjAIrUenq8PZ4kVMzSUnynNYSdpUdxLfRpI70gJ0XZ1A68DDTwFcuQXIrmkvM33gVQGaQThb7Xw
G+s3kmwoWOiYwXbqbkqjcSWHNje5qASYPPQR22lU/jTG1Jj2CDWTYYcKRU1JyGss0FJ8komtTx4D
85d4s/5iQ6HZbX3qhMQTwQTNPvZGpR4F0zMPA49O1FD4CdxRNe+qa6n9ETp0uHQC9zMzVPdxvp73
jpkQitiI+79Qa6E11moHWzg9TL8Z+in3Cl7ruRHZ2B1H/7GPQZjRNz0tb98/WIwSx+PKRCNazotL
Fde79awYfuhjKFM7wZb5E0dK7t1jSPwf7i3C2B78KUiJR6v0Fwuzj+d5G7zqH0IDnPoKXd0R+CsQ
6Ppw1hyORPiGJOH1eEvIlDDTj1EtY7aDlQ16zVHwKdyD5AOSiYLlfa7fhKKd6LZsm4aMP8J5fGM7
bZ55fm9Glr+yDUVRN2sKVcFSss3I1AZwhUC12HqOEqx5Kg5PKdi+xIdS/kQmU4QER1Ogtfh05Vl5
bK4MG6YJFWDVXCuJ3AQ0KMHGv6rCtMExO/HdrgE38GSuhrj9oHZTC/r9lnq73CLK0fEce1tXtUQK
OzWL8Q3hmCo+UOSUx2lAMiJVtKATyWP3/rIy+PzLsskXyIjN8pijI3Ki9TqP5iFAqCRfiJbm0J22
EFeKdMe7Gno7eWv9Pt7Heq1ZASfSLJ5Z1q7TRp8ANYxrd26pRsoyNgt4SI/oAmZTz02ufmzfA/px
twJTnfQgh+CO6Agq7NeSWezVFGJ8V+4Duf6ua4EE+SL1KBsxuUgrU2N28BqE4mVgYzgO+MdrIh8u
F+1UOlW6hz91X1ycEoTwcbfrGIXogE+7vFIWjHCacViC195g96R+hiLEIk3G8A5V7Bp3jp/teLRq
TzUka7spR7fnqvCB52VIzQ4pZzxOJEQ04FBy27Ki3x6pFUkm62gLpwPCxMKpo+k3Ac1rA5SGFA7U
g/Zfe9q2k1wmtbR0NB2/Kf6ArcleP0hzs1Vn1GDmnzRhkkziB6N5S0TzJ5Xf2Fir/VlnW8DhRdi5
Es0hLC3ImNIQRPlh5DdAUl9PyTsT11f+M7UPeSBKn7nsh4h8eZllVcQT4moHcMZ4S5z2tzBKZObA
DC3+oIY/uVmoZnpk6hEEXPPt5Pt9bbliKNqlpwsIJ1mnCnI1wVQlkf1v9oynkZHgyrkdYCPHCyH7
+NALBiSCd5I/M1o7mkmnFcQoFAeKBG+5tM6DkU4WvaGKZtA4d7Ab0j1be8vZzEVoKMHQ9iByAjpZ
QrLHjt+kuApgD9mx0TeMmulnXwtJKq94cYnWB5abN8LH8khrtxvTmFLfVyvT1HprwhfGKH9LTqGq
oBLgBTCxgH55rvALszJDQUI4IQVZmIpmguL5B0M9CgKjOA7oZosOYJe0Te2d0T30yhg0OaLAemlO
HlIBU9vHTRY7KRmyzN8vIkLvayYuHVDuNELR/LzHlFuKo+L2C5dfLL8qs9LKOxn9vcJALhjmuCzc
enqmEXcr854M/Qq6cIB1gOJUoaO3GGU6rgWokJ/1QcRbZ+HaLe0ODgrsL6x2acXpNvwyLYzPUKIo
leglATyDDt2xAri9Y6/K+7Ykg0VwJMjpyk7nGQ+60PrXAJjSy+PE/3Yj6Pk+NgtgHhw4t8cLpBLv
0HmhVHu1Nl6rcgK2bT4yWwZ9lYiPaCnDUyKqEbz5VGoAJzcnK3fW/jqIUh3SJNrVxkv0xkAJmf0+
up6VAoxNoSOOPWrgp06piR2auln4kO1wxvKfSL2n2LNzc0OHuGSemf7LdXAriaX+P4R0D7aUZb7y
IMD3BNKc95COqiSQdL8TeYj1Knuf9O+3G70ijHODqOhwAmI5cPyBgSEti4EQRv6ZtQa6SZj2RIqQ
VPisXG5NLLcvLgTmf176NbdsIfzw6wrnaj5Rz3UoXsTrIB7NdPxYMCIWyYKuAejXp5h5ltCfBWty
JxuhJd47lLLigS71E+mUJ1OXCpjmAlpbHFbuIClkTrLZ9Yrf0G4rgJ+WcqC25i1ce4ShnrxM7RJN
KDtUfloqORcdujp1wgWJ4Nu2QKT/toy1BUhpqcyBZaSPhdGTD8gIJDrGufoqKyexOk67efNn6kMd
AxUzpe3M+RGS2XS10fV3FTC4ItGMIu1sHgClvEpJDOweM7MbW46fypbkfSXK5EgKBpH2wwSTODP7
TxNoLNBAPSUg/1lFnBm3ydRrpkrBIKxQGxtUdsAZAPwhkh5zc2o+ehfvFEYkRtma71hnIVNtshdy
rSXNnPvQIZJQlJ3dh7jscR6XEk5omXD6ItY9SZ7h1oP09kkgAzrJn2A29RNNJhcyx7ZcX1vlFSSb
D1IF9S8XbiQnyA6xGaWK1L+2jVr7thHl/G5V9uCkUWgwV9oUFLaS/rNDboUJyQZwLL989Q3GpdUn
Et1rkuDVGatZvNXcl9kieJqRxT3+Hdozwe0N2EQjNb8J0UXFzSziEikekhFX0L34nEQpC8MAy3ib
K9HfqRL0HqUSRRtyqKsO6jYQIb+TsZ+cgHGVVMwZsNt/A7OFeW2Cl42BkUR71BllDQX86csPtlC9
ZwiXB314ZvulZFMX3brhjWyiSuB0cg3jLLqKBL92dOl5FSXQizzc7fbbsyPSpPEierffSNtw8+Yw
BQZwdfcUjg+tGbg96yz3allTjEto230a9v/Q+ju0HI55Xr+K1AoSa6FeIhpUFELDsg7SR3qcIHYw
ljf/MfAbubobovi1L1A5Z4nIj9IMhvBraR5rucbeRdmY+E235wRA8ys1gHMUdS71s1JXx+qA1EQD
dC/4+p+ztXi0HJaB4EJ8IUSn5qTop05LnFR5GEE+OcYgndv8mlVj05TaG1XBtoTpATCjCyafmhgK
ZajvOfNccSj4kSefv0V3/dCB6P853vZL6vmbpcRzKwBPVJNScDQ4IXATNgeO6tYRzu7VmrltEMCw
8PU5AmabEdnlNrXsPQnNeHP8s3Wwe1+f3yajAcEc3gloY15jwpXg0kSd9zQIE7FbVtWptrbjGgsE
PXXz1YJ863sLqONLOgcnwi2LjR0Se5lzYLg8eYFIgs194wBUQlEXM6EAv55RWaxHGhtrl1ovXTZf
/vyT/aNmW4cwBElKvWpW7X80NMs5YRyK2YQAb6BDmb5iUVGh4CQSWo4wLsgIA2wYDOqMlHq0YjpQ
x1Yg98TyUn5Df3Xs7lgKipMJG6FaKdje5rJwW6euoY+76tJZKdPJkNzhGL2z6VR34ZzcZZpjYAdI
CfnksqTJkBJZCi9TsSJzMb1omfuWUBb10jfYBM8+zTtbKuvwv0uAONhNZnOeBPDdpkUwLrbRDgxs
EQBnQvOPKTO8d8rfwPNLMbYg2GLNPdBx37NqyLErldKd0gm3Zu9qWd+zBYd61quiBnoUCnV6NiOz
PzmBnDM7nGrYszXjdH8VLz72nk/S7irzE++sRhwinIeW5HMB81btp6MvB/fu+difykL3HsJKOUR3
f+XEgPSh6S+TwVb3Fgr2pf1LGDTGbSRQoZE9nJxMWbDMIOkcNZ8ucxFP6aebn/2lRGRxqGrOv2sG
pbgqTaQLSPT3lwQfj2EfpcfioKxDUH4I1o1Vek5HWgKL+itQkZwkz4LS86EDacN8+rLDSoWlw3Ul
GKUnTdRfThe6/bNO6xCLMFEdy1f9nGH8u9AaCOo2OJ7wIVGXWJOVmg4/EKmaDDLmwtG3cma4GLKZ
tqJCiCH+PDj+N8/R/J29QoKC+ZEIK7h2FreX1jliYC1e6JWDT7KbW6w8WSdjHy10ONHCCiDNfb8B
wgd3RKS/BG5SaPQmcw5/VO1Ctpy/VrLNb4fyEES/CZARhsNLX6esuLoadyTWte+LdbKjsaR7cYGf
r+QDKv2s1fp2UZyUC/nW0s3+um8Baeffojxzw0p7zMHpBX1f3IMvXyMGGhEVFAs7NN/hb/hogwQ8
rBMKIsaWyrXySNeTMdnhIUaAAu5b7lageYJZswW28E9eEqq5VBZkQkF3/v+oiLOKkvIgykR1P3QH
2wLKxrVtad8VszMHbZWclBPaczS9ctoToEhK9e4Q6vf1JSwO2nEhNxSK0BntRkwH8bmKSpUjIvEB
rYqk2iV4Kk0eCxSBbdjBdjfCwB421quHOeMiwIjD9ATSiTwPzRfk6Hv2PW6ZYN9YVUe5JcAk5rvx
1hjmK+MHGXkzycvx0jScYnYMmd2AgThIah91ISeE/qVEu6X9BJk5iXkriZlTANW3qvytsXSnp7nv
Fi/MHTOxHwU6cfvzNNEmjd4ahkqmkokLi5cx5jQDuVKeP0PK+pRnQoCKj038hWfFvt42mOMtT1S4
ygR/GthTGygvu+hisHMASQGeV41OFXEriEJ1e6yRtnd1zoL4S6QHYtFuocVjKsDMeOp2837Cyx+8
8pNHrYSKQlsA/W6Ch+HvrWbFlwFCUtBMSsCST1ntbxWokO3ese8ACymF9gepVO62nKLHKXF8ZmYU
CNoEolIsqEZkn/43YWE0mvC3w8SsioxtwrPq3DnxPIM0UqUZO3BSniXB8qqbPB3rKqhsYH4AKZHQ
Lja+tINGGx7KtXQtuXnvtZEA47VVINakjYdAD5bKvlQUaQuv3M4Ui1gOrJsCpkWzOohLUC6TemRe
xIHh+MTOi7CLm8PcBGDahzYmpLrMRvgrz+elgoJjtsdYzARNFM6ZAne0VPDjiJuIQg/mbpE6OQdS
HNXfJMtpG2IL4d6qnPOrftEWeZF4p8MYLzIYmybJL3vYAOIhwoI7gzTKWqdAU7JadCbP6yDHuCNO
tz3qX6vtJpAJwkk4RVkgU94NaF8MODjf0F2HS4ms606J681hvG2fMUFvwZ3CtS/QNL+UH4Mf1G4d
TFTim3GMAjEfxaVsTSVAA0BKhkE+mfDQojDTCa7zfy0NhtpfBjh89fZIf9GaEhxA51J9QONVSDPj
K9ef8xi79er1MkcL/4OE3Fu86cgK1qORMVjcF7OpynNkpZPH51Q2z2q6wKfNlo22fZVLEALTHqxX
fqrBgibMwl1keiV/ljQ/xOELyvE9F0RpnEY7LNen5o7RAgjaigbpFnTe+G3tNEF1A4ENkLOllSNR
JK4y/cUlhmzeYizLAfreDVv+D1EM/VTwQ/yYO5Dc8wK95aBTSnoXxWPAiu9vJ5FEelfuraA6Tnzf
iFjaZZERrd0bfBpLEtZPGptMR+O4AoOECw+AJQLOmPwApMKz4O1TwJgtgQELzfuMfM9T/kKojowy
6E0LgtIsdh/Y+HnMP8yMR0hSRFm37Ed2I1e/CGdJWnAazUD+Nwl49pyVJh2/qukqIDBLzWH0PtHH
rlgoAWuYHDFcpZrjyMud3iAk/edE+EZA97dQZRJSSaZp/lA7LYH70YPFXjiYYK5Tii3DKxm0R90D
B05ZQP37QEkZWEBcBWaeCc9px6RmPTjdRF5jOpBs8qQFyQxhD+1voDZqjy5PRbB0dwFBq28rvmoc
ergYTcWxdSZNmit6TzIJOj/oZEKMSBmvhGMQiGxN5KDE4v0NlbrhjdQad5gfgXInYij5uklml5Tr
da8TnT0WWjSZF8cab69r3UH8AGFhp1cDIpphLCF1MNbbP13SRXhGmNLNCm/iodz5uVak3slOETti
J4wWUK4Uyr0B3DIW/P03RohvgnL33imjppMBS/PO+uoHhcFBXM0oxbHMJ/M8QqwZjH/46fN4uWnp
SN6qb6OSxizXOGDY7srnL94ojFjvVag6jJB/NV7H9c49p38d5Ik9ruZWwpYQi4AO5XUcczgiArF3
ExnUAlPNxxAZNDJYLNBaUne3FUzGxO/JAEVDoCM20pebO1p/yoRXOqHBby9k2zFbYF5hMkhrCoqO
9gLWGwez0UQ0/zU/STSJ3u3uf89wCDO1onhkebOUTN8G9tL73irModAA9opzuppSKYE59Tv1r0r7
jMQ9KAXsqhAl7lv8EJ7ABR5kU6YFIpGD2kM6J/I8e41GR8Y31aTydGIn3KONYaJ9UmYcxzb1XCA7
B3DZPW2OnmQu6jqIPFP67pA0tPCtGoHBsned2My7JJUVB1vWl8/VjmR75PSrwIW6jAZOjttJCLfp
3BWPhhuPZ7dT2+lQZ5Cwc4xA9iwq5qVgQr3v6f9Wb8fvR/bzeYLQcTIeq+MwjzOWhUueHUq+UrPo
BEqPdVal6uo3AzTp7ZeLnSXfkzSh19e4mMb2Y1+ChFu7XaPv+oAVITYL4DXR4ZVyj+faxvZxqQwQ
r4EK26nipnNJ2TP2LJowuod6ebO7hdnVuCKkdkJfFjAINsGapSgjOicK+iCEri7rN9YwXQuO6vBF
H3X2wpqZOgy5ZRdrNLo9xj0PwjPhmA5ccGg8v00OdmeJVCU2R9qvn7HSBSth+R/f276+1j1fTR+A
6DwNXlKNFRl4L4J57GTkOQ0Km9LZdIogdL3wBX1t/cL/H+o3MOtfaS0CUZcEYzFIvbbowN1SzPur
feOmJETvq4lqztCBVLEu72febFG8MpMhukvElypx4n5xAxyFF65xypfBDKl/7WrpekEB5UnAcXE0
24kAsl1e1F1EEsKqmDKpdXg/p9BxTg1hMG7wW3fZ9/CWhCehMV8hF9NZpOpFRKea2wvyUXIeFYf9
FTpLtmsTgwBXYwYrenKLAUYQV29wMXonSavb9+x15wjmJCee2ggIoXfbBJgp3dq3wyhziDdtwuIS
+LWbAWGZM3j5n/DANV5YRFTxWKwx1Gqy1aVY/yUj7CTV/fbEf7bCLeUUW8dGQM1k3mYQ8N8csov3
2+VlwA79Y19DaUwD8j1+v30mb4xLsP3xh24N2Ig4iluuOdylthSPXBCZIsu/Nr7iuACTByGVcFnb
Z+38VCMilDGxDhwskUm/vKhMd0DbfnpkAuGedrT6aK56ZaDbmd+w6pb+GzVB1ZuTUKyinFR9bhaQ
MGE4ykzi6B3FBkFK57nL33pPoDexQo3A16Sq7JGLYNXmiOp6IzLqOV76XU3KL8z0eUvvn0pJ6PKv
lPYP/1Bw4Ss4wAgdQ6+PFcPU+6usPj2glDkbR8BiFl6ypZdf0e/RPOreCYehMqAnK8c4iamZi4k7
bpx9KKqFy+uE5r7FqQatkZ8wLe3ODhNB784rDagIPyvRqA7ZQ2FKaZa56AMMvjAg1Icx497FBKCG
4GkZxvzLVQCHv8uZo6lr0u6wv/dBUvucfEekTRmyqva3i0ClkqSqyj9qugx3eAkYOmQuAe2UdZDv
gHhT1GCeeCXvJYOCvLW997/ywG3GYgLcc6VJRNIyWBPxAnPvDHPrCIxcnFh0QJknkRJnPlW2T94A
9zb8azkGgx0alAPbmZ3P7/gVRHxvERJ7GTP4jLq/tBbeSVkgy5e2PIgYfd44Y2O5pT96f3GP71Gl
oqAVtgHxPK2o/DZX9yVDjWy4zmkOvB4OfWs0FfWNBAOFvwps1FsOXaB8eKSv/CvfC8QAdsEqBYov
J5EWaGgISKiTD0z6XPBVnfQlb3hS149pGQtoVLO+VLpb5u1CxO2cROHN/0uW8uKCk6+LcKK2XgUC
vEbCDP8zsPA+qV354rcaHSq2HH64AYgq+puVnnVOBwccBGMC5XaUmT6JcH2m3aZZ8m5ObF8XP4kN
mMFrRzQ4cywK9ZVMToTQ1NsaCoeOMHR+iLoA2Pn8aIHSQPJJ/h63Bp4LK7ZdLxmGoHOxI0i/Z/j7
uRrFR0eUErRQr2bFbDSNSH42t3YLEtVS/W6DgDpzp2Ds7q3rarLvrqhwXLD86btDcfIHm9hJ4S5H
ot4AXiD1DE27Kj3cgKHLMoPZPSf9LTJ0uQAWL1lCoMiYpnQ9Dsp+gmNCLhbI5y9ZAZbthXSB52I/
daf9CW4rgBMbU2hu6B4oM6erGjiJ50zcZhoNETiZg58aHDY7gPb50tgAHXKdyosodfIREddrr450
KlikP21kPf9DCfhEkVLXYCES5VLFWvb6AKJp50IHEneLNrcFrt9z6oPUNiofSrSdzO4ZtfOfeEc6
y3+GuAm7/O6c8qHUyMGE/0aAswZa/RqLBkywsqJk/XYUsbbSFCukvX1pWTTM+G96IjRWhDTTkjC4
r8BhBa2bMVwXSFhOERWpRmG0JFn6pi9RfPzEK00slswJ2X2QVWShxri4CHMK1na0YUw+bO+LG0Jm
fDy+0Vh2FOk9aSDsBIEt96zJXINBrkc8fi3l3q4CD528oOxyF5F16YnQhOI2Y1GYtZj0f3zRuRK4
28SpVx6DeLieulT32y2GNGZyuoaab+dZSwNan12DIMkVCeUAYTmo5fDdjaeII0bRD6W7kL4kwxBr
Nt6/DWqTcZ3XW9h2OTZPe5LW0RZEo3dOyJV67rFxI/xc47ZvRgaSb8CXywCPWuq16mTfwhZ4+NYn
X2SZE4HPAOkIPEZXs1eQRJ2VuUdUQmg62LRSr0dmA51M2PDFieOaCW4bPhlMIU/g5zBPRKRzNKfz
1glqYWvXuVXOPFjasdl+nEQnjt0FkXj5yNOppGaN7LOb01lHzjvZI36C1tcnXFL96oR4gRo9voGl
lzI4IsjPdqO+FgtFHg/zqHrPVXhPDMAD0ydWxi7cc82DaH71Aq+fkdPk1+JIMH47CZF+kZ4BT1iv
3JxDX5w+77TIPx9atw1vLphDF283eypakXJ52gj/M28D2poQ+j6FsGkAt+j48mRCBstHMg5abtX/
BKUR1BZbAr1dcwmMNALxvZibGtOud3Xi5d1bltI1R5teXJ5MVp4O2D7I7E7VBE9Mpg+j8sJu4J+P
Ikmgb0UWqAa8Zw5GyJN8r0Kv9IMibwaGnSQXVreKCYBQLALp4enVRH3eGf1UrVmIEnjM0ySsk7+M
IJu5IdzK0WAJ03mFeapLr/RXd6DjSlrP1rFDJgEhzInGWlrU4GNVdBVllvY2LuvfvDfiKrZkOjo+
XNmtB5ndsZncTkBf1AJ1d2kbueBgnH7A+32LRf2qlHy61FiWmlwBD29KWe4kbUi3gKO50kG34qQU
8yHq1iLfaQDmrjBZrhSQbgvw8S09XlHNHhrMmICus5i7TSkIvpWI41Ox+mirDvkl7P8ED59kpsEw
Pti2bK2rPjL/aVNjnKqnNPMu4oJYB2y7oIWKZM2jYLQGzqw8KQf2hEgD2xIGwQzajJt9skHxrjs0
DFpXzcKJIXWP9SHvennc2fuoI0Q7CNWEcsC8iV184nwJ49Hs86foLoYqtDBH3zLm29zvPypWu2IK
JwhdawlVjopFtefFNknZBR7s0GTylWlrCmP2daqAQ/3IJ7XyLHQ+z6422sbAHQg1hwUgkzrMFFw7
H1oGL/TDSqGnMo/b+ID6z+xqN3qP9a6vvl36ntjsezy3TTE1EacQAx691+QH0sNnGh2RHQOpTboE
tNcbYu78G2fw7q73SpWbLpcoBrkjUJuU53lyck8VHIJ6O/c6u3XKCuBcObTxZj3xMaLuHZ85x1Li
tTO+Z6rgCEANfyFn+IgzK9Pozebu2bnCmE2JuhB021jF7oTvBK62u3THgzfslY09e2Y83UiaXQTA
4jWoOH8d9LxvtLvvsa4iCwMfNNcXnFc2Vgomxd31Qwqq/IddolQPq2QV1cNMPV2tJEe3YmJfXGC9
AetsathMU8C6ibceAZgzBfu9OSOYWdcJJu3Kj3HIL0Rk7nZa4mSoAxGrYDH2tA6IQhwgcKsKQZ2l
Es8jqhyQQZWiOu5O3+WKEpVGdW15unhFcqqYilN6kFrIOoydVgnCPsuhFrcxEnIzIc+VlSiOGDxI
vTo5rQyYUgLXR+4lRq5cagoSyebq4z7NTNk1zDunRrUFKU2Rbbikf1Sn5xmopGTW79mVaFhbv9RG
WjGLnP0E6FstqSZHXx5eBgYuoeOcA0qcVSwrwv0v281zMNKFJBsGO/i2+sNOC1SXeehXOnvkgONV
dFUFW/SwEmDnx7vZxFO8VL9jgMewwwk6RHh0IfGAy8kKZqyfKcbPFF7u4IxR92n6nnuhG9Q52tMo
aSl8Ipl6gBHlP/kgFJoM0zXeHGA5NR+OBivgz+nll2QZHV6g2XNHnswuYJx4/xcju8xiY/8tClWj
aKVYSVATOktG9LXGGiMtysx7NpOZ0SR11a7PyAsHf1rY7ZKxcxAGLlAknkA+XTdavQc+R5M23/7e
XFZCTc+Uct00sBeejORPQPzyRRb5UFOfjChbS2hykmgAtKQ8NiyU/4nuCWdX2QmDUAaGsOe42Efr
aW6VQsht4C7PQf7Gx3swq7TGfKM95foFyuXnuvbrvo8+guPgk7dqMzs5m11i4pWU1YplPhScHAqd
kMe/w8s0us/LlNsEkKfzyrm3CckaWXjZUZDs2WZ1yWw60RG70VFuU0HPoVuYs9HhyhFmZSiMvJDx
Tygfg7GCsCIFSybVk1hq1qVipCqTjjfYsdBvASoek/EOS3JQ9rYvIJ+uelwDHUw5MhPgL35D7jHB
AvNODX7al5ETV2ThSpLGidSyHyiTuEvNXwU1LguESk4KkA4kudRY6U+p0Vj+1YvTA5OE3xU38rUk
TIa4BI9a50XxEzCe7BajGuVgHUI6YtzGF2Vbvnve9NGv9XCFDLVxpxgcroDJqZs/xN6/oeR3wxA0
9nGN4Lbn1UODVhsscircSKQ9Qc80lQH6u6pKGjX8jsCPuiT4H05J5gI2dDroTuyf4sY9AlkhnO3i
Oq1VJT9pWasc/Z4rUIi8FoIQdzbheuq6h0mU1OOUaVgh+9jNjbPz2lcTl61WihgoDvz8wCZ4svbW
ab9qWSteLW7LBEAYqINxh4Qe3i4lnmNBerTB3l23qL0hUEhelorUAY7WMGX6ApJBE7T4ATsvvleq
0W0qVw4g95XAv3kH68edIODgXxvlzgF8k0ZtGyLnrrKjuHrAUmsrUdwv7eIQ9PCMHgUeteMV5/vg
LRN3IMFMKu+iPI7wy6GdWzVFlGfoN7FPBcpBfgKn+j9K+HMpdwQdUjt3247HTlshmJ2Wle/Ym70P
TBM1VyJf94a2g6IuN2Ko3WKLr+vou13nW/qy2PUGjbrsdMDo4EUH5tISs/IUpWapl//K+5Im66fU
zjrlFo4/MhVMlhju99qgbzITS9QdugLFB4sJ6/uxU7kVz79LYNGkMoZasMJnq+RPmdsedI1Z2aAl
/ngZXb8l92MhCi6qKQuYm2XUoW/ClkUH7efvLnhgin9qlCO4QIXOpB7c/tswYuLy3yh7dkWguq/8
qkpMzCFnZJNBGYGHljFGAbJZzwUtDDxgO/YTmix+tqmrLVtgZ88KRflV2Tuwyz2j3+or631TX5ly
7aL5pG1AUTX2fM13MEKHL/E4z5o0Rjk0ewyyObAn3+R4vfOBL6OdU2F2j9BkX9Ov51pv7Ugi0Nh/
/Dzy0TmzmvI6T26yX31NstU3Eo5s2pQcAQTsUZ1GsdjCkVxocYQWuIuxyqD8IvTvCPYGhOVfyfOW
HBKxARp+mcoWCtopO1jzqMdOaVTdJirWDfQVSvDiF0kUJaCvEGQvoI29L7wmAOfWgGfpT0RqLwss
W2Ea/SrVqcLYH+ztUlhft/BytMFgjlNpqFzLh4OTY10qZq5s1vE9lK+NVhKKUfKS2O1UrXJ/7Wzs
x/flTvG378eFCHCXZUCuYZ1vgW6/U5HeBEM1IcMnQCNhNeJEiNjeaxCRZOshjVSnZ07lbDT8hFHZ
Es4DxJ2RxLgvTazTn5+XA1Sg6lxfmaA2drJOZIAzhQ1IvLAFWDBQQ10RCvynOKYTM4e24+sxiH2R
BQYJXFIND/RwLWbpTUqZfSsKvSunu3EnLkxNsW1uG1fEff8qd3BhWr7b9F3B/+ZF53VVWke8B5LR
PDGgd2H8XzZCoKK4Ws/R+mLT95y5uZnNlcZuyuKnvFfa6qrtQlmP931u+/pcgZJllHx5shIVJ1HG
kT5ay/F2xM9ToDrKBqS/ckePRqDrdvFYEdNeZpEcu54XkJfHZCqaxGBdRq16WQx4vm7Xu1v1o+ME
JHSKi1SwMAcqnH2lyuCqc4fiElZBH9jbYhdS7zob4hBkPPdY/54eiqdolEvK8Wjq1b5gVL6CwqXE
mV1aB9bDihl0jnl9i9ZOfVRZ97NFSdqG+KDxY3GBYexzltPT8XzkRv0kZvD1YyaYq441M7hkV0/V
k+7gvcdPU+ImiSuI/KNv9D2XpBKkJ+q+QcVA3CpGHCd+5nQ23jpmtSn9WSTbMC3bFmgfbIGUug4i
QawL5GgNjLkIGFdu9vXeSDj5hH6a68sWOXJBc56eIY/R8W9YMZ3EdoEQqhsv505nPEgaI/kRL61F
EQSW9kfBcwB4/QdtlO3bq/WwEtStRihlUynKUG9tcYm3ZaqJehr512KfWz3GGfdpDZGJVbgRMslJ
zoXA/g+PzWiq8Exwrnco8xGmF3JwadN2l+mw9U75D1p7UgjDiPFXpDzXksX4GnFwYVLrdJ4w3/YS
pfdSj61rgoWZB7K039SuTKBPe1km5rwtYB2o7tmj3H7VEnsM/7GsiessVUTKhVInem7a+fTpSS5+
J40Y/USIo5vy9sT2tmbg1it/1MhB1hPOCud9HijZu7Xur6qTfmfUYrMzcmWuk1ELpBNEHcTVVcbq
wDD7Y0k1xdDOOM6WCJme6EwirVTcK6LKnRiwtm0jeK2Aw+3eo3KjGxvJELJfD9PEMdxiNrXmJbzc
b5R6jnew++DQ6GkfUcDjWotGCxi7wZ8Nm9gE9Mj1jITMysukOKHVYr7fWq/OX3KjVnXnHI6k0dBi
1FVWyyVxPu+Rd2VOlDZ5NLe/HPNFI6qX7igG1L8Dm5KkLGB1a5WvsNzwDN9jZHVOYrTuXWtzEKD8
P/i87Pwsg4KseK3YklRHqXVhbSoG3ZI5oBsCc/miI0t2iOJdWHL581vDXxd9BUEBgoCg06Ai8UM+
FTsqzB4wcqQsBYDD5uLY0+KAx0e/WqJn2tFD/GdW3i2NyF/K59kxb/iCZm353nhBAq2BaDIesiBt
AB6NsGAy5pkguQ+Gu1GNfZe1epR8SYQ5nTptd247B5n22OeRd/61KoWPVx9ATnc7SN+vkq03C/OL
bUkIdtM9AygrTQA3GofwD3ZEcvjhZV3RV58Dz9gkCJfXwIzzqGTzeuHd95ycDtGi8KJmFVY78BXx
bcAzKTkXgLS6Lraa3weqyEddfm8+MVe3U17WtWF9h0jgy1jSobAtRAp0KD4LBT5QlQo5IxMJ5wgo
oScqeaUAvr9uVLj469cudatIi6BJNGTnIDXAUAMtV9WNMTE+oq9wCuiiUQKHxReYmhEBdwSbAq/S
1hP2cy3YOrsuFOwRYeUTpDsJ9tixjaQmz0rJriNRQIahQXbKx2nBssHhtusfWJ1Xz4ivVHIr3mmL
ty05V76FuJ2iOjUUaOtCcEWYJt4q8g5kcafX/ZjSPzc3pm/neEVthG/S0qPFNV4WeQ/aoVPNk7ML
ENRYtg7yLyNzr3YM9jiCOhcn3oZgnsky16CXdoP0Kjpps2xN8jLU7I4lZKbA823ZS+PWjYLu9fZ7
Ht8vgz0+GfmtZGzcmKho/fG2B04uUTgbFEdmoi4ackxSiXUNW5IrNEJew/vH2zhFOGS07IIe54UD
zvv3lJGAOu6c9pzSjeu+k+6pvWgqp2KqR9V8BxfV7hIkcFUPb/dUkcQKK7rxDaDRRsKOlHLc7GCE
89ebRp5vVJJUr1DAdpfhNhPMIaLmLfw4GBMWkt0nmYSiMofBaWtf3WS/H+6dGk3jEoD1LnteLKvT
DkVnwmNtd28dNeDnRx46Xars8B4D/CS5A47jyUr7gbFIeqyjNbYp+5MT+IqkpIv9fh8TQC74knp+
J4T/0PpwqTx9hPybY6e9FteH9GfcTGyO+O0qmvS5+W9W5J6n0d/Kl85VmWPKKmTUQi5oJt7YEXW1
VH7aUZi8REB5zQML66TSfeG7SHdtItPNBaCGywX6UlqJZjzPxUdCyep+3iuYa/eEAtPpn1pPwgkN
lDTjV2GvYBdrKpI71waK6NzdH2QKlhlaHxEXHqPyR7Z8A+1mSNFH/9xxActz+eGXuViYqbqISZZI
BfKPjEFryNsj2ryaVBWlHZMH4C8ppCcEzR9qC7bEogXrIN6piYHaQyWTPNednb6jyrzLCzv/l8rP
T436UUm9VG0vOPlnSRYXORJbHhCi5I7tfP8OIGBE+XgmcJdLXadXQx2Ret+8P+BWoqqneVWhhYud
rDgQeeDwrv1JvMUvbFQhb/3ooEHSg4hHM8YuhtvxaXanmfhU9j92kSoZIj8jyfc8j6ON31168hnb
1MC2crf5BhkRPn7noQZeNRRAo0CCYVNHUuKO6ZuJWMMg1xeMg9PCkEiskR8O/eqs8ux6xqkK1Aly
4OuiIAhGobd9MHn6yNAeg4cFCDRRBelNj+9Xj9HRHoctgIM3Aqcke1z8bQvebw3mzb6wUDturD14
/Wtg3iNYulhems5TkccVC7Y4R16s7dWGKIwfZioKuZycbhTJpvIRuNKIykyGnBgJHW4lWewSXlpF
TCC2lPSqbwyV1dUDPSX6l0u7K/RukeBZJIZ9+bqTkdIKVTRp/qAIsSqePtaITnfE5RHPudbjB1F+
MuJhmhoYtZqjC6HPkNSpUuBwnQMq+OMST+5nHXVq1fuh61+uY64lVBHJ4RYiMEjXrdXYp5Q2NoAk
HTEPmxvXR4G8pKcZeK6hrBd6ShC6gVfz0fj7gy7PWgOSt+DCeXY4NxUpmuCvBCiHFSQlPWuRZzIF
mrCsNycV0k+D1B4TcKpgLOFYUWZ1VnTwCiPNQsHH8qA2mVIeVgz7P6hbFGnQmEQYZmkcVrY3kObU
2+nnIhqC0haSk1BX6cSNfD33LIsxcZpfsnHzmfZG76/mfuxOlDLePtNuQnpB4YX7xMldUcOOZZ4n
XTGbJc9c3v6z4LMaT7k19eawzczZ5DbTOTYpC9zrgfjpnB3ttvcVAuVyMzXirNJ7cw85roGctsux
+vpmGVLv6WHex3Rp8JQl1eJIz4Jg1Dc1H1EYR1IPrwiZbFkDtOnvmGrJs4p3IFHdFdoZJ5SU99vD
k0ihkol+Xn/ukNi+qDhsDxTv8wMM2lX6jD3/PfDk74eGFg2soKgRC4WOEUvKPrzaPZVZ/Z3rvhCA
j4MRAKK/Z3VoHffXaJZS7X+TtfTSFRbownCTSudqw6fHu1WcgR2coaAWWyrbNXJfrI3E59m1IeN8
aHhVMTfDZlg5Wb+Ljxu1KOmtziRaktG8loD7bmfYKE9IKB1G0btkSEe2MEv0X3N599G6BfYko8D3
adK4FkXjCl8RgoxEWmNIW9X0jSE/eUMqesTKu8PyWpIAmuQApuicJqJsrBYXfJKG6631xryNbkWK
ghLTg1wGvmcPdBP6eusszDkEtQo4ctegGX0M7HwwpvZjhbc0pWTFTnCXVJnOSjSHkRJ7F7ouGdUi
C2gISS/ZSDp8vBNYTRdBmETu2Q1vbt2+Yd6bv0x0KOjzSQdm7dwCak4c5FmhwNTuWBfSDOPaNMsd
b5RDRsFOohTbmOzJ2Vakq/TZ0GAzP9U4ip+c2j6GkiOkeIRBwMWR0AvDXceG3+nIDedgNWmrc+Xt
laakw2zNuOZ+trhgiuoD0zoSZp77xr/NT6Kp1VDz/iCY8KSQ7dLj4fza7GmtDL8CeApm/EiVFoVw
a4OUvYDVwFo5+oL0VrLVnBgbEs57UP5OysfVwLXPJhI4u+RT/nDKdu+ZMysD8ryChGn0scMPpPxz
ayFnR09uCSag3jqUNOBcslxUJMwZf8ohDFu+XGu2rY+jKTbGELie7LM7M0e10HShxqQi+R16fw7P
YIN9BaASQjjInNFQR8s/QnZUGkQJolUxQZG3NOVLMLOiezGky1ILoSRO2fg4NZewYHPXrOe0AilD
sEj7trYpbKrIn+gvin6NToT39ooagFux6/L2Xs+rPch+Ll0kkRUb+n8QQaE4JM6uDuaIS8gQbLUA
M0RNBhdY8aR7dSc8bjO2ZwZqSV3s5ltaBZRIWOpD+zpsr+eXzYWzHthvLBkvVWpCbK3UloqbZ1jG
RAthXaqwB6fNHk1OnUMaAFdlRVXQYgHkh7ZbJf2CFLEnxmUwRcNsqo03CpMHbvawEefPUbVwn4W3
8EYHL2UA6RZnayjbF6VzpLKAMaae9bwMeAhSw1pYe9b2jAvJcVjxBdMOL1eHKAvMkrtfWW6mVHPJ
yyPg1bR25FOc4fsY6MN+irFM20xznkGOZrIhznjPFAwrRSYi0/xmMlQpipIrKslSN0l+Qpy5+V8y
uGM6gn45Q7jQVsWD5iZZN9ng3plaJARgPmf2Kx7pcUenIVW4pqWTp2jEF6hvfkVB3nheLCLasiBi
jmSZPrReyGR8EokagSXJe+Oqk/dk81Dz7zcXDkE9LxT+ghPKe2+07eWCGObAGxTlZn141dyFPcHf
hHmG4k8Lo1EYVxDWVIFURh7jctSp1VVcgr4RpY4QSn6j2gQk+KkdBduJR7ep51qPwkqjeoKmn+Xy
stJu6kNVEloN/lAeREf9+d1eYez2tloADSMHyPxQbQAZaotG/9Ov0wJ9X7JymGlNrBSt3vFxNUk1
osSuffSkA2bx7p/0RGn2XXQ4d1vSz0E+l+613PJ+6LRpE8zQlDchPVkpab201lKBds/ALNbPMWYW
aROiUA1R3uv3XF+j3oVejtgeNBZRQvP7MwlUv+D0Fe3fXncWbTcF8xMeYSGla9dsMMykbW8TMLgh
qV9Pjgx8MYjrF5j57Lz7fg0vSeRrfqwiBhgs6hxnr/XtBtdr08p4KjvzZwNbWIQ3ftsw9Ni4EJaO
MMGTFOXzethy7FkrpMk+92YDZr5NP4z1g9AaS+Myni4IIF4jqSn0HiZHp3sX25RWJjOl7k0ISRDy
p/T5SChuXqwcI+8wlGSm/FREhMxAjnzMe8CBpskud1R+J64buH26FdE7A6Pb7CsYVZRwlg81Wmrx
LOnMJpVjjTuqopaEWo5jkpqcm6O32AyUgCoZ/trbUt2Yu4aO8z386TaS7WZwxGyNuSUkD/WkBHGL
q+0dOwGyyrXETjqe+XHCB4qcN15RFY15BmhqS+I/O6/R07Y9APWy8xSJVVxfDtxHRI6cbJE/yzcR
SBXgHFCslS4QirZfZgVU3mZbAWzu2fel4A8rSnh7xWYr2xku5pzg/1fcepKfmajjq5pnJsOCoZBN
eNfIa1q1ARjaWdEosvCEYmt0ZYTehFXa/G50zK3tVdTA4JdiiUextA42kRTAfzjgrQQbBoo85Kkz
f9A5mGcPWVqSQ7jw6oOKANIfvWgWMPHgTYvUmHLllzQP229MMmBq+LS8U2HOKWIZjMJtqXghqutW
oKE4NGqaTW7BP89EU6cBnbuBXKcwxrC5XMcUzaphJfhY5ronkGnTBz9qiT0w46fRycHTz+nZdLSc
wJ8rRw13wFampqdJavyjByHm+2EKlHSeY6N0+XeOII6qXA44FWotGGQKsoUzSFyiXmyH+H5TehEo
BII+D2XDV7J2EEvlQWFfNrirGuLJSztKe1S5ksEh8rAQ+bZs07Iw2MTKs4+1LpZpzaqFPl2GrEUn
qDo4OYy4UKPqvoEfW3fpv6ZZyJGBHR/h8ftoG+7RXFcNEkEwr5M6yuTozlYxaQiAGWIBJOQJQZNc
Q+IfzmnPO4B0ANTrXK6YmzWSDaWsTd0mcMCnTvjpY8sB+rRGmi9kwkqxHjPNC0VdEuG0FF+k/IYg
Ce6n2d52EOAqaTqjnhfwEkuQkLalNdMjAZCbMq0A//3AjjB/volrhAeHUgEY4oEdPDJrAAYrp0zx
tqWYL1WralTwW0HmBtoOwfFrMABUzy1eeABvcJaArQkoe52mgCC98s37ir6Jr0cQJI7LZupoXq6l
Hhq3U3ASLUyjKxAedHDQea8NLbkxoUufaLVkKGFCOMQAib3Dci6M7PgFxbCX3At2OQD/j38PHP0Q
4NZzyVIBroG1+kSy5gJQaldIqR2Zqk1WKJmcw+hKaukt76jiPr49SG2UHxFOmk4Rtn2FhtXIIC47
2vEH3SHevGWqX8NkSiavsmbXYPgtGX8fZhDNToiQymRLNTugF9iPLByE0kGvJLHghboQP1IOBzrs
QlkNRPPNVANe7qN29veZych1+C7adMQ4XcWDKglT6EF+GjtQ4ZBkcRhx3hs0H+bv9/P2mACDM8ea
FZNGtJ2odTSuCBYsF41gNFiJen8I3yuh3uVTziu6G/sFhYI9i+mKvNEy90NZ6+OoFaTxuMmHjmXj
rfjMeuATogMhbXmK2h3kdSxYs5UAhvF2jNffBZIC73J/fWZUdAjmncI6IEhYtbOzG+yRe98l9OhP
vITMXjVN+n19FPkpVdqs/IfONUd/QEyNkUYx80BduLdgYoB8b4+DC8E7v8fl7mOePfVQSr/bqdJW
Ci8iQn6rgFKceUp4NKP/5Xs946nk4tIx4RBSAVsSaJ5Gdqopk77hhTXLaZWCCXmbqZk68Yrl70ce
UcrF9h4+KkF7Y4igbjG4m07ChxG9a8Twk+V4FU6QyAqHvrBwl9RjBreB306tQdRa7cmEN8AjuFHc
LaGTMrxe4V2xYQOtvLoHrU7hlZ/Ya0Y08tb1pJOtCqwSR7Rm0hqwuobBYoch2vT7kbwyf5/AjKse
knyKA5OdSQ7+D3aXHjHtU3q854KbselcG68/HEHbrc1gXSZV6sDesq4eTuu/RljKl+UIt+RZaVz9
3E50E39ozIH//azyvNcCuto5BSjGOzfKo4Ly9hH1yNFnvbnhAiiDLUXQ5N08lHEvCrWssCYnB4b7
vHuIdrdCOy4KbYXBChiX1zZ8hvZG7DXvOoagf66DU1JpZEC+2gaXBok3Rpo/rIBnDEdtyyLUga5J
EM5d1MCK+fAJe5t7PfBIZD/xPqhfT/ItoRyOFAdW5D8JqOaMebo/4I2yk1HJcs4Q7kjnF/UbKjJd
TTXJ06dV0Zeywg6eUFJ/6Ai8nvAcqa4d62RC0pr73/QG7XyGA2hi655jfKkgPvJyKGLCVuTvmizK
D4gaePyokDG/CzyZrdnFC4RIsKAbnjbTg8mVjDW5FTGf1npNAYmG8IQs4WyOkyQxM4Pa6gtFDqZo
1WmpqqvDi4dYT5CIwUlKdoGxWAGuWXeWvUjVXlF+9zN0nM6qodD3Z50b8rUUruRvxQQbLJTgbt/j
nPgUrNdVElvnObXISdEOjYSq8ysTMIesRoAQGTRyKMvdj9garI0Ei7eygjPzq/ck4BSQ5rbTlx/T
XqJVkgVfZ7ZMdeDEh1QYAKM77FEQ/iP9jFG0+f36eu/RSdhjElT8Q6iGpmTAlkkPicbh/j+y5iiv
Wh58sFQBPuBwUXghj3B5PR9B1Sclo+P49vaqYf3bJ5Nc1eRFcU2BbgvUO4dSGiwddCYkQMzjNAqF
Paq6a4tt4sE6hx0iflT1Gxj/mTHdG9ImIAPzIzSENOTEgpaLhb+XiAZIAO4C7FF/tNOQKwwcxFm6
0ArFjk7F49D6qGkYco9QBnIcxYiCti115kL58SJNLVJ0m1SUD9b7WuZ/9ajrQVDsXClgvMQTny8e
sCLEbHefkVn5pQ+PmVx0gg3rdnfQfCYa1oyuW3XifJ17IrRZwR36bNPFBjIL0nebrFncz7n+g5A+
JYymOSMDRjxllwHmpcegaAPN1r0/PIg0+XEm/gPZDUmsbl/UR6bMived+wD8UgHoSkLAaDN4/eyA
zotRd6CVAEUgi8hYJA8nYHaQRaQ/oNC6wgoINxs8yVSffC2RU8t4imHEFptSrysn1qdNjH9VohQi
z6BW130o7UWLCBufIWgHzwrEoVM8gNf+wl6SHrv/vzSaDKa0qfW7DOIA7sGjqRhVr3VqXSDcZDKj
Dw2JoyDuHJr/1i0J1+HJUKhJLtHnRPYb0EOrJpnL62VikTQ9lkUH35SzllCSmN/pxVun1wt1bAXV
mYQDO8T/VzSnFiSV12oZ8UAox6p4BxxBaXnMejtDaHwrNgHaC6er7Y7oG5Kbqs3Jx6BVLrssMk74
/8gzf64bYbcXfUEBmA2aKP+cZTBEDilDf+h2jimSPkfeO4kK8F8UvZ2rkJGtXtCekNwU04HVMzaH
mOkbYr08LytKH1fzIvccJ7ulXxfteRws/axPJCbrz81sfuTgU8k0aHf7DxzGCLTDKSyDf7fwIAFG
N/GmO28x79zhZ/GD0d82WoXo2RfUNcWkWtPm4QqvqjWWhrzGg2NDT9lmVAX4eorxtgvEJxssAttO
/69HSa5fd1j33qDjmBJri06oivolOcntTvB0qjiWA8JgBoJmwhAMzru9keoVhLXj3IRa65V7QQrI
SQd+1gw7FwiICaUoFgsY+lC0gvEWTMXNMXccuDHg0DCroGrcpJqfhQBVulqUb9wDOecDDHa+pm1P
xXLZcXoIrNayDhO5Twa++9XA7nVD3v6UUvKpMwEyy6R1IA1mTDIwq/ElgUepeMAg5JawB5bCNNsq
7h2b2N2/YDneCBVbZStLYh+0Kpf4teC9VvcEAMqQk26lO55QWtT6L0wGgGh3OsrvqWta+8OGr/ME
+37GRvknwkEk5eMTkVqG444nr/TNwpY0E/z1pMntKZxVg8owHfoC/+q12EQPQnCmWa0rT40rSG5O
U/VkI+q6nZs/K0j5b+mCtgjpUP/z1tSzka8qUt1SLL0QkERprhLqElH9SrRZX8qVsHvKUedP9nLh
t/qQI9rMNrMeeLQlsNr8EN61zVCuV9qPD/KRO7MyWggb4ZCVe8jllcG2ih7ajPV2B+exQErKrAau
ece7N42OeUwU5ASK7JVGkUtVvGdB+JHsb8WrsrHrab7LTLI2+EfWyjvCeiqQmeLa85I/SO5RwdiW
cClfFM3TYbg/IXmgLnNM2Er+jEnCYqI5ahFNyGA0por4ZitSuC5Bhr3B/zziUqyv33dyMPbTYVQp
1ugStJpHvgonuQJGkdoWuI/i+JTujjXZ1QMyfq6s5MbrL/+aAJG0PY6nnjN7aaahY4kGbrJ4Sc3I
7+8IfqQnvF9GH0CvOTGCIfPjgTOLFCpkU2do34D58K2XT8erAT0ZvzxZ1vfonIt2E91eDQIai/vd
8d935XHYgb4FXyYw5MigkYbedc1lQoUEcbke6O52tWpllXN7gODKz0Ek9TCsbTzZhGZh+oBjr5lz
qwjGOX7+zOp3C+dq5xSlZabjTrmVnyohkAi0GuJ7Stoi2XhrfnAT8cUBmrmAfH2cwfftbu4gK1Wx
DJlIOBuBJvsR9TdJSJB8J8g3ULSGv/7fNKfMpu05XzXfUijW3dSCC11tW7ehPhlBj1IsqxEK0xDv
g2MYXN4RrOMYVBxZVsQvcZsnRlRhdYLdVWop80w85zm/28pOysK9Sbeawc0ZMcDRePSlAKiBWWVN
nDwq/IloYpPg3SBmLUNv24VklMK3a1+PnXwfmRihhEp/qhWapUd7UycXek0A88jy5ykv2jdkqtp3
4WYHCfWBfRZu7CVvKa7Ouj+PjUBGEFirVbh8viWdjCPYndUATs8eER7zfevC1HW4kXM5IJmIx7be
uo8FAOeoc0+Tw/agD5zpz3QCH5uA2wdk5iqkK6jpKLCsmZkpvGJSW22QviDDJFMlbzvEAnVj1EmG
FE1oMbE6u+dJKs1ciYu32ITjES4NGU6DBoWMnE9/oLFaGZ5ocgsq2rjSHa4ZsN3hSRJ2Sb5FqtY/
Y5/9NWOiyZbrtGwx7ezSdcRVBta75IeJdYw+igkHj5gnpX7uyE/qji5TZ1uI/W0YT9R27KEAllBl
RGAF95geM/7sG5tggD6R6DubK5nnwQLguTpdbvZ031vnjkQ2jmTN7eIcTEeH4Dr1xcDVf+Dy2/3o
ku3j/xO/uQXob6xMKfjXd86tiAbCVXsfyfpK/hpHYiCKTQXNvY3Q0sw3eRbcrV8W60xzB/ZFdo/K
30N2JIREEHhDOWDhAL5PXVA6mEovxojPZu1pgJIrWIc3c/zdN7CpxL0Z0zNbTw8Hcz6ZYflAlFH7
lF9fi0BfWdWIrmljG+0DXoflpo7wNJp7ZZ8hXWyEWqwu8rWUl9Hs0ogC5Uzva77oxv8mn/K+5VMZ
awUViJnT8GWVAkbUHfvY9Zt0GiuP80pdZiC+id7QqtLaMLD2Pq2xpbJktGOQvVWlrUjEANaREDI/
yhb1bw33rOAgxwahKcpKtrFD/cbQa2JSCuEWvn+Oud3J0P6a5bKOwKFfSyZ/9XAprLhBdBkDTf8D
JR3R8thenqvIzVCfzh0Q8fEKQXpS02JcVmSlfanVhihsRpPPFMvDE1veaQN4Gh4maHAyFMcoicJ4
YBVtwSt4rfAX0/96O8YjZDZWyYU//I07dUGjmr+u7ZqnlRcJR0l61WZzdXvZAxDe7kDxqdf90x+j
fYe1k2zeecFFpSw6j8gBoiD3j9915/B2IH+GaZqNl12lilNy6Hgn/uLYf92/m72NzJDq2dUXZkHv
Ja41Q03cthPfCgQo7SMDKD9XVbfzYPRUPikOSQwwYLKY7PawQ/4cagp3wjCxHUYmKIUKKT++jRZ2
LxItVfMRWDFnOYchaAKGjOH340nRh8kDhjUJJ1T2ILP/OR9U+HbJG1IpRtfZmyyOgLfx8TCWzJrT
vW09gLpv0t8hdN4oQJc6+A8MhUbk1b53CfYRAds/U6Wsda/5/LDn3A1Z9+E3WsxkbfUaVq7wWrCO
OXFhFL33/RFGgo888org7Htkh/rBhV8hW1+VP3qTRev+HmMimJOpf5u7rx+3nu6Smv6QuNWKjNxH
KlM5SbziwPQQMEBtM/Tf0rjasVIqfLS/k5NJmqdf7KDeSEGXfd/TOcuGAxPK9oBWCm4L3ynTLV1D
e2xNHiXCskgmmVjPMfqznLVEK2pG9CbyLB21XFcNQrZkEYBK/g9wnvAn0TU1Z/aVRWtxv1/NrIkl
52feZ9oD/ZXecK9egb1UjsPHA5UvhXTnvs//4K8mKBDn1nuI739DBN5kUqWcyHIkkl57Hm7100xh
bL2aqqswS21GlHX2ljFcdgyR1iFrmOh4nduRqQYg8B+5XckibV8dLpZ07CFBlLFqVLgggOWnQo/8
A8Msm61o3qtYu2p7ItoVX9JijMzj/iJujYRbnS6bAfMUvZnypEchvfi2fCgMMtRdw0MIV/TiycsL
xB2U5s2mCEpE7IpKWeyFwevg/U6wyXhidXrkcTuPCQNzqhnKm3T2j7CMreJzEDJTlE+PzTZDVhdZ
xg3wzqTkDmjCOUKfhG1PJcWNRQ3aaZVcf1rGny3hVyc4aUt79h5R7XTgN3H/00uGNp8cehpiIVyp
CjmC0eA4Lkeap3cpQomIRUc9Cq8nzNON5RGXLZETxIVikbZn23iAo9Nlpd4glTr+6nLCzJhM7vGh
bKCpX6O6ntWmPw+iRR0iah20Njvhx4uRyzCjSUBcMUlJbbmgnzeRv1z+RCgwqxLFnaEM9dAhx4Jv
nV9xI43KG37ZzMNhcYECFhmtN9wy8nq9Osqq/3o1avHZ26Cd4PGVfe6r1TySVEDSLQ8uupko+1u6
asa3c2RWy4VZaOUS+khvbdxDGLq7bhM0zs9toliOmPEqLc5mWBbxYE/zEIiJ4SxGbOzWSNRfh3D2
XabtJf/uJLlsOzWusDxs2SLWnaubSdSHYiuEXtGPjUONZPRLTybB89TaDpLjbOpBMrYSqi76yVlf
8J0l6IQOJ36EP9x5zvOi/gLNvD5aO1sOQnk5SaEgApvDLZiM1aXVcZcXyEdGx2cl0E8uNbVrS2OZ
YA+YbahA8oMztHdD/cGoHNNWyUBcg9Qi3Nx9UfpnC3yjTgvXs1geR/j2MiHn3dFEoinRA4aJ3phO
PJg6AyJo2y2X2P5WAvI6PNgSFEL1eFbPuxbXrnNoDQQQPas127TkrwcX2ujMs8LSNItmFXF/tWfK
apGW7UcD537GeQftH+JkGVWX5FSt48/rBkHQXyCmyG/WenGMg5D1jJbgqUYiTc7T6GVux9jhsC5t
Hps45ComP+jIGHS5pFKwmAhzNicGfw58NvR8EJ5iHpLwr446Foqjoc0o+/qV2D5uogqM0USSwaml
eaMqhxZvWtgFeovuPgxaulQFKZVwgt2XJygEDYzur9awBZV+ZRBPNhMipJ/Jx3Sb8v30Pg4D7SFX
q50KQ6+04aVDX73buPqiYaCxxUnrUw9KW1gKvYV4cT/gWBHVc+77OV9sghhKTo0AeywKf5P7Rypa
3WPGtHjxhXXCxyVG5IvFjq3AwDNXwZjR4hWNuFTMd3LavqgKgWF9yWnq80nlgmjZjAJgQyuCib1r
2ZOQZUEFH5bs536bexmT/cE+ckC7MfF9yE8sTuGrIr2bnwF/V23nQoFvxCt6h5Shr+OhjVzUmfdO
1DR1BTcaTEeurXZ9YkC9wjGu2IvSU38v4K/7RcRTUupHNBdaFA9L33d1FACUaiBJF+5mSlKi67a2
mS7tKhRTPgE0EocDTsI4e761/DQLEsBYD1i9hRmp0Tu+i+sGVP5cuRtmaHYcNkJhUMWmmGJtxrnO
qshfyEhv8lq1S7lzNX2xw89Fq0OLMhxc0nXld9ZTra0ImTnsJNJJMDBa+OIgEMI+O4+FHW7i8mRB
oNZauJ+lBP0T7PdUn1ud8DQi40HKWvdjyLmdgAPzdwKyk9qp9if56qtGIGXwsYb2arHtaerHiRr3
zlwQH8rd8ppDYyOdXGqbZR/Zgsf+itBNFUYZ43yCB0E/8X6sVb28o712VTZSe8au8sStc6Smr9wg
LeVzdLjtJEzsF/kmqkrrLOEJyDAqHeunoSfe4ciI95LuataBNmK9a6xsWLLeiVwA7N3yrzmRc9mS
MKQ1sLEWgXOeMuo/xq9fTbAJRSMOsl7AE18aUmzOQd4egj0fdjde4rvM02pG6I4o8bfluk3XntBf
GRa7TaYExlw3kPGSpErY0d+9DMhhIN73Mrd02JZuFc0GkrEf8kU8nSpd0jwbTy6eD36U69QptgbK
9dHHS+o45XeGdq4+oiu0lvyA6ceMpEhDx6w/aBBvVXJ9obDRoYWOmSs4VJduJvRTe3WIEm9GNLBb
EiJrQ0zI5ZtLogJyDRSeIRl24n7zV9omFVrbGa39CctbcFGs/GeefdLPsk3icvJuRaiCkWB60+W8
uWHeYboAEwp6bABWVa/Rm0InnHe45C1z9amDc2L1qLaAap0qzCZeY758at6sI9zfa10/ArC64a4n
sBakwdYhy+EXN72dbEkMz7i0mrU409imCBRbrMfxIlgMmTvJsf1ZGQdaCCeq4vbf0ZjiQWw6Ff0H
MUzeA1NM2IU1UJ7aYVYZ4TYRM+SmN93eD6o7APDyUmbdT+1NieXwsa4nlmu3B75iVcKeKStzE2Lm
oMINVZYmA+z0lpLi3evqNnXLlrtdFJ5f2x9SEFAHMs3vgs013QeWeoXILY1ICBj+yYggVJB5B1Y1
Sx0pkxeSyIl1GeDB8eMSSVWX2gjgNn9ehMZME3v5VY89qmmfhNkV2qFjIXufoIXHvgK8rJLMRyMM
kh7ox2YQ7LOc827eWt8pywDcNefw35s1/VKT/RfsWccDjs72lbTPFrOessSTag/3EvOpahJsxD8j
/gfTtBzxnBV8wa4PGOSslUhEbdlqMQKBD5M7QkaQ+p1tD5FK87u/pP1jE4mz1j6NWuFywwsdockK
SBGntU1ComfO/tAYGpRTsJCVYv5Fl7PRcWFKdcrkjoSUR5aVPASUTRs2Z54xtetePNgh31l1hAIq
gHUCHFczLxWpWBCU/cpib6HGPAI4hqHI7vE3tA+CfQ24VlD9ozcsEUFjrHprKsnLtPUsRHCmPvbe
MUZi/srahZxO9LZnYozO0Ax+rs8us6CAqpFPr70uvLcUIeMt0Hp8osB7x+/xUF0mSriJS9rbC+ow
zuL/pIIImZgB34XuG5Av0ewFvL+S0+duWGR5khvo81rvoVhqNCNcDQ5qbPQdq9G3TatzTp5WBYOY
z6LROPBDPFI71nXFTs1VjucokLvYVOdZSDd+t85ZN7zepkjAzkvdTe3h8wcWB3J+LbuYOcHUk4G7
Bb1Q3tgUl8+CzKCh88ofGl+xoZyvlX3KQLYYpR1246OB3Iek7tXx/AXyfRPp9jLA9oUt1VbIfkON
96w+O9NZHeisqsaL5741AMjd1f7ES28t8A1V7y/uVGueyCoQV62xcNXVNQAQRP+RQWKGCgqZQTQl
V2Eyx67pfE97RqWEU6gwdY4/7yp5/WBuYaW5/k7f4B6EEvtyD6qZ39mrbkPHUwcAlOtMJpyjwswQ
P5fUmuIPItR7OUV22okbHbLLA31wR69gZBITo1SxmqWNrfI4vUmlp/UkfWTsudSHKxYXEw85/+h+
O6ly5CzQWWCVGcfA7n/YEUbvqjMfbEYdiQbocLzzGhIB8Pv+FyT1Ng2PdX+bfTvqM1g5Rm3gDGhr
BTTjFGgssn9YJ4M54YPReFtyeZtEWx/TKUzq9+rB7Pp/UDnzgUXZjrubtzmFP7Amii31q0GwjKmD
bSKt7Ya8IjUIQyfonlzEZmLfVAfEajmid5fvbYP+Nwww0pbgM/rdsFTtuAFO9CWQb7PcrsptWF6l
w8oeQ7PTwWoyT+jpQW/inAbCXEGcn64Fg/H3FVGxjg1Z16er4gM1J/2Pmdu72pIuNRFAsMlqJowH
WBDHXKKcBTHTuI46z2DqE2mRpOyhXRGbd27UR/p2hDr+tOoEY80TpGrZPmtDZTGOhb3Jl29AmjUN
z270LzR1G+C/EO+X4Xza7xaI4I+BDAyOgVqTgMBHPWwXYAXvkapklFRCFdZsfIHz3kOwPZRVPE1V
0WQIs+rWogdli31CgJpP5jhGuPl5eOUp6cfXCMdgHNN7v02NH7M7nNepuzKYUVUO/uatK9f9KsIa
RuJGm0WcxuW8a6zsHZeSLSheZLcsgRHR4/V3BQ2/aVU5W1uxhkrffi0TvkxqRqPQKDjmNSvQ3lLN
HpRA6F1HJQ0Y9bjup2hUFMIWy9QHuYEyobFVDdJ4UKxZ7s6CzbOZo3oyirDkafcyrVGVWRdbJL1t
X76itRN2z2pzwPSA+htykfZGky4HBtAy5bPAEiP3zYdaxW0cm6ILB9TySBO4NAq97kUaUC62UAjK
b8TpRC8wizlHye9ARlpT/xVkTLcA8PadieTUbf5lUzD3mhBVKyeVA4UIRLTqFkWJ2IdDsfbyip72
5rm163y88urzIzY64cX26CODuVEc72BZB+Rvry1Kr45ZWY3VmxI1UyP76Dg9PlUvbrO10Q7oUqNM
aKCY3J4SEHRBh8YHKbWvlbSm1B02FoDExsGW8qexenXk4BuW/iP0jAhFaRWz9mZsqBOewP/hPQZH
nxrOFG/37azlOAjQlU3WsFowTjcuw+DZRp+RCGwNLsF/kZXC2RHLUWQucsT+FCFnAMjuIZ1wveLw
hNAW6ICxfMw42zKUaCE/GRNLUgqPdtdOcWdosEowqm/taMwPh5AfH63swTnUWJpSbaB9XBGEviwA
jg7DDAbOJwR2RMJbhcO9i9MpOq7X9ejjp/sK0B7S044l1sy0G5I+oz8t5zbNBAjROKqzkzfwuDwd
SJFOzeLJKqqPc0obU8UZvKE+bqFlQqwvlvBHMbUBE8+XqcdZomXMPBrtpqC6bjLrficdTOL/Eyxi
Tisj6HKvtAMMPDQZds6UajRzxc43711wRcSwzsc16fgWMPqeyweEQXwA87zaI8fkP1zeo4UpDtAP
CWQR+F2Jiz6xr4Ix8TBaq1M77DEtAggJzsl1RSZAomye3FvlpDPPGjVHJWt3ywhbvhyNPoDQ1ggY
euy0Ebxfq/gUZ1YThzPv1Z8mw5QOcPS88HwJXnHVYqGHBbk7gAIOFgSEoEpeP/1TCy0yKJg+1zRN
v0S2zxpUBpUlelN4OUXfSf9qiQ7Y8IwLjWVOYOF6Y9Ee6L0Le/F+mcPo3yWy2bB7yE1Wd89bWif7
GL0ocUjiSV2QV2lzE7ZtdAFx+p7fSpmwrlQP7rxmi+3MS5IvkDSk6csD7r4iZlun6J8eVXNy+jpa
1HtB+Bgai5BmQUT59vZs5GjbUTFMct1I8tNxHTR1hXElQ85G/fOFDFx5sJSurDl1ktxZkMlkT65c
pn+qBGFn4z/Pnx6iHrdUDRvDPn0lN4OahY1mK6sGlQcTgmpP3li5zZ9l5ZyiHPZzSO56VvpoyyCa
OOA969uyLSO6CNkX2JWKe332NKWUS/i96fzmQhKRFUsIRGSLhFFUy42/BvfZzXbyKFGGuFJgnUNx
T+9g6NyzEtC90ksjbNau+nf2mvCp3tK3S54Yi3Qr9G8gzF/DPeWu37kNIwSab+F0QgSrVd2FC3VJ
s4n9PAPXjAs9nh4qbRqr4Ws1CEUhvIyTKeZERfS7YeddJrODDlS/rgVheTbmb3Cv4vUQyYhe495g
uMJkgxGO0bx9WD/5Yumzv7+1bkr3mA03ugECbpEvYM7Fj0ohMIjUGhh9vn/Il3YhxPvPgFtNb8BW
yWgux4QrmX2RQkD7YQfipj/XX7aFSuK4pg7PxMIBrMx3L4XQGrTIzhlnY19GruA55GEPLclVoXXf
mWQvYb6OkumlrhN5mTC6m/THSYSoRcXteN76jrCVi9OkQ4z6MLLXawsR41w9LTSsaBi6SYzZ6/1f
+6MkKhkx1oQ3bQX6yoVXKhEgyItFBXsZyohHo/YLG7a3+sdVz1pUG5HBFPNldT47dovEFxah9tMW
tVbmL2lHGoZK1Jhd07Lo3DZD5zUPVMl7ZG09DNX/0OTEShKR9W1JnONbiWoIyujSn5CtpwYIYlXJ
Yk1pVdFI9UyMnca0fFkvfmnibvBw2Ezm/aZ+Qft9LPBApabuxrRuIQBdyE8i4vPVfRgwurCmnHT5
hMvbFSAheJGdcYugQdFTHsv92x1XGARRquxQgmeQtU6O1tV9CGMMDyzyWb3yDYG3rt1HNG8S2Wwd
aYLbiXu/HN24E4RegyDKhYjox0+GEQvvViefyUj2KHw5X0RXrIduiQ7IfTMi1+NDYjnCA0Pas5P9
Wjrsi+yv5TxMs0nWV8ZsTFZYvbx8oSq9FyL1SJgohBOa3T3Y4HF36GSvYoMlimsr8J9qm0+Ze1vZ
oCLIRZZZ/D4kpO/Q528ErlkOJamXhE4twopVA4TgjjTZRlKM1eUGJb7kU6ftRy/jrfb5NebIhFfO
1mbjfDCbt0Y23qvMO72yCIq+52jhGPlSWgShKzm3WH3XUR9TLzjwQRt4lnez8IvclhWl0dSqeuGr
JlSWidcxRh7rGIzCaC2nBcR+dqCZ/wwoUIHDVDAGLilRw+lRLj/VyELkjCUIS2hA3yRTH3VS8KBR
qWv2ghPN62HJr/SeK4R3q8Vo8JY0bJZ48mGuyuvYOgAtWm2Ld/mvcSbKDPd8uvYZq5ftAfaXbeXC
l6eGiQnC7hxin3m0oGqdmW8Mml1QCoSGErn5tUkzAWFwbVKlnj7fl/KeHdw2TJ7PEKuQuPmhiHmc
8Bxe+M5rk+jzIWFFQF3i3bvWxK+qLiM2btzn8yr07J/RO+pLFlvTROXn9aZf5+5gX3rasZc7Ep39
oAZ+0lAwvTz4tJLXcLUkb/eLJeYO32OEYpYE6WjiUABCq8DEa/cj4LLAR4nID/j22ymfhXf9CSlo
UjlkNsqfhUmeE9K+bjYiQlzDX7jmzbcI3Sv9gUyh9bOm6tfofrnqRcseNvxONrb/VYTWMjenhU1v
7AXyR8M4+qyF58b7O2tkh1q3v1ycfmVWl1o2Bbkso76WvmVJkxlKtDy1Vgf1m7E101pko/m7S5in
Ym2q/a0NgKUDKepjV2X/VjSn99B7pn+iiC3cgJc/kBf3JImbNXm/GpFGJ/qh2WdYR9gVObubuoMD
UIISFhIN3tllkN85z1icMesvi5KRpvk2yLvNgcmgQzkK4v7V1T8rZcj+gMCd6VrWqWSMXbe1hO8U
pdxsaznGCCerBk/HJ4IRpeYuZZ7FRjb7v3n3Et8UvvEZ86WPPNAPOsym66LF9M+Cn3vbuyhknOli
xu62EbNgZ6IK7fFwk/2tgM9ygfFGYfkAb1W6uAqRwwkckTjjrT6f6B8GeaV9dUBimeAQz/fgD+kN
4N8LiqKnfjCl/KWtQ/IMFEH4+jf5UeDtr/N6+g+utco8qHL/SFbAeit3wmpOnYuxKtU9L7GFtV3D
DQlfh/qs2JJP+q/2DQZMm7ZO2s3y128ypMMdDWORWvr5bjgcEaVHXdv6EPsokqieubf67wG2UtpQ
bXD4azTFvIVLqMMCtSqOHgiZhd36NlkU44Zy+0mETolBw2tkEzeTF0U3F2u4zqNmQ3mJrP0b+A1A
9g8ybRjqAi0Yds9bsK9eIYhZZRbIy4iq+BRHOlrBtGKvSVx4iHBfixqWyKH5RnIKxAPYOXQlS3CJ
L8TyNMX3st9u9JyotXRRjms9gi9NYGW7Qpm4a2jok3JopuHVjxqpSPMwy+soohoEouwqveN1fMcM
rfaefhjPdG5kGgcJHmrAjrNFqttTsMFrHp5MwjJ/uerqgnAkjl340WqzlyzA3GBhrO0h0ksOL4sy
Jsy3VkqF5e+oApFJidL8lnobe5pB25rBBI0ML4laigkdh8YKQNQ6nsQ3FfqDCpscxGemB6uwTRH/
7cKGDS2bDWRw8b4wBiy536iLyctF61wmBlbAAenPDQ/5Mnw0Q712uYWdWhM8xWy43qyUFCVdiNKx
ERTZNlGK1sboZdAQXwaZOV+DR8n+h68+CKlCy9hYVg79Lh1BXfIOpLZm5b2IoM6A7iMl0FnVJe5l
iS38O/3V5ordhpS1iDU1FL7tkL69V7h0UBKSNP+TSjT1gdrMBmeDHmbMuZezW7w14DEEV6xu/J33
M2QEchwwqQMjtaxSJmkP9Kb8ByjszTI1F4M/D6kCkG3JGrp/5TqMp32Ia5TRdXUiqDr39ihmq3fk
fppJt99VEN/Je8yfSyOfoqPJFAY9Vde+EeD2o6Wkf3ri0W7gFb8wXYFZLMf9EG6/gCOuF5eJUAs/
NOMevN7WOnp4OlmOW7ohJifCSOfLn5NaOEYRigEXfPC3p/MwA+uF8x1s9hyvsP3HLorximnuuZDI
nHuBEQ390LnugB/LrNFMpxPYFkKEYPzE/l3k3UXUFz3z7MOnX8oy5ZBWrKEp++ZpavLdQLYnebdg
nbK605X/su5GT/zeQN9cPL/9Kact5eg2vAMg1iIDGApRMCn35Ttz954QQ4CGRZIggDQ75SsjqbmW
wR/v97096U9VEkPD9AmRALm3ohTItxxitwEZpGpRl1wmbXsvcGFSXEuse67jnMC5btLya9j6YGTL
FXjMXvvySU4561qM1O+u1iXay9fEuo+HwqQPPqrJGLlNdgpwv9d4tzHi4PlHBRQhp/UoXS64/B4k
/piTMOk+sZUHRAV0BzM2vYJVToZGrUDRrxOiUAmSjuxBNiTt+GU/SYOklAqG3oOYH5icgYqbHqf9
hrC8ZymXEj+OSvoSDgQVLxtYRQRUfmDx+G4/36eS2n9XzPzj/0LxEZSA0HIWJY5KmMkzY13CzoaJ
PISzCkT4YIsgug9X9KllerzYcQa9306c0odv9FLTOzHDs4r3lk3rBxIQiynjTxdsgKnTs1nLNkEb
djM0Sf0ca6ag8ddGw3G5fsk2cOGrA+ysoydd8T1JNyajR7uw0Ygq7eC2hpADcahSotehwZazHInW
lpu1+LOz64A4MG5U9t9slzC7J80ZG/LFQuW+9cayOnTIlLulkn09pOaQMVYoSEp+XWNIU1oBF3kj
RAR08ES8iYi31VBf8ABz4h642QDDnT8Zx573Fw5FsYTF1BvG/BAdToUN4LYUJ6+RgRCE16XQiW4p
IJwYkq6YdC8p2WbRvbUGV3Alq0mecu9tzO77ktpCboaayFkyA/9JrQWrKk3oVKeJOTIUVYk+KU+a
2l3LVdUtvbHwxpa9oAcHJpds2RgwuemDjYEqFbfnY3XpB/6JHsjdyhMRA4s1tOvEV5NHeg2RnAFR
jEQMKdHJBdPeLcD8MZnGjjiuZJgifOivWy4C2bJrE0gRXJqlWK3KCkfWIhp94kJnFdmkM2GYh2kN
ojGWevkAGl+1ze/Zs/QPZiKdW616PzNAn8yjA+rqIOs2RZHBgFVwi+Hp8B83HCVUWZTccdbn4NxD
oAEJIyLt1aKchyEO7QQ2gxOsbUxfKMCpgDBe55KFbR131v4d4i5QnjtiMWcVEbS+a9JAW0HFXZW7
XHvLPqZQnHjwpekrKXxMT5RHh6G47WVfCxoxpD9CdG3QjV52gDt2dHS5MIQxEEdXmy3bWUzMwg8a
aQTRuuAPqsIPJvzIepoadQZzFl7sB5friK0zpvCk6oHpFk/I5JggPxjNSo7IFSPgCyVMrsD8od4g
I6ubJE74Fown8R0rNDMW6zsRdEW/oZm1EpWOC9LNgicNSOYbSMnrG8veTlfYcvz86xlvnZsMA2Ey
ZuVdAYlf+MfRCr27+GFtzgRZ6YvXVvR4mCtXTr0EizkNqMVI+AGydo9XgWsaf3sKqYxNRLsViHBW
hWblkMsHE2gS0PGrNK2Qx6L01qNsi+MeF2l1tEme/Hg1C8e9/y97iRqYe4lIPgS/5kIQVA1dSG9c
gXvK/MF6z/5Mml4BI6EBPBB+8OsmOGm5lhyNiMEqoPHpLZ4Hke1tIZ5unBlbKQXwS62NCLtD/2Nb
7Fw4DMGSf9AMV2CONbVYV7UMS0LmJRM6LMg5TiHNXdNPu15d4+lC/bNeHDk3JVpImRhfTyAYbTFk
T5ujChjfVwOkSv3yoZYZBoa20WATeI3hh/gseTikH7i6NI5glQyRJZ18GPgoXlv7Cpc+HOOP2P0N
DnQNFhj1uP/M3tEDh12A1vfkUigy3euCvK8rg7qgn4wxoxfa+lKneU8nW9ELOXykJNJoM1w/NN/9
tjM1PSIgk7ZIReJkrFIEg+RhP4XkCIohoLj+OB6T32rPH8mJRfC9l98oLWjv0zA+LFlaRx9XG4mz
SEBUf2XYKk/j4ubforX4giGbSN4E8yv/OjT0GlDllpS4Ggw74t08QGQRyWgEK99vl5avG5HPF9iE
CpX3K2hBSQ6ggs7ftt51oMZAoRdEwv+cPjKFOH9Lej8Nj4dzKgCFDwa0BsCE1uQxMXZxzyHIRBMy
4KqrH0SlN4EmcjfAnyj9SVHLC2KWzOD1wKbefNQb7b9dN85XwjU9/EyCPvyw2laVso+buQh2iYD6
vxtlhy0LBFDIJnajZqaxigTZFi4HDISzdpLyfidDKF9V2zp5YzoBnjNaq+gDWhbT2ihI1Yfhd4T0
pmYEHxzKelZ6FbFhDE8NuT8XKiXfcEqmtwG6KSg4T1QOmgJIdJhS4mQ2n+tYJav/yl/Xi6m5MxuD
kY67Baghz8yOwTZALNr05YSAN/0P+plT2qoQQDGMSuugRezVQGXDpM4fI+XpoV9H2RcCvLLSZ57e
+p81S7NdcD6KtB1wBwOwsWuwH23aqra1nWocnbJ9EhPArUnEXtdFkVgEmj8Y6LyIQnKSJFgNvc34
r1/TxEQPniocgGEl7q2XR60DmoK3Sr5OwirtE0/zbr6Xi0cuNX3tscci7mtqS0dz3VET3lzsYxOY
odSl50QQqSGI9rBD1FInNu45/eVBARDGAQsPZ76LAV2pse2O8ODYlE9ksSdFKVndMayZgkXa6F/B
25jsi3Qc/5qd1jA5ynCQamXHhwYbhwyD+uBDoa9u60iq2HNCw60/Pzi/J/35p4rEqGshguZnNcVu
GFEE2h9aGjK53QyWeU4Ob3rtsca1j2VPRRBL1zpwX/XnakP68KSQkrzAEHRcbN5U3RpPuQaFheTu
CyBpWOUx4fGyoRzY0I7poo91SVvP0dUrErjlHeQA5h4bp5g7mpqNz+NZpiM012GFEtVmQRoGVVz3
qabyyYaEvT7+wR0mnhsRN1pKjTeJDZgqXH+7683SD7STlntF935sJFF1SjkfAYjE396YmN0bhkM7
MYBtCUSTYVl+E+wwRRd7GINxg9mVgEvkbCcS/5ocyiErJVUUT7h8OwexJYyPCB4YxpI6o4RTj90O
cJ+pU9BaOYSZDxBhu1uzNPhvaRONfe1kBJ+NcMu/gH73iI+8C48VnAvbMljX4k6DJ5MrXsPQa/fK
HGo31XVObybSGhvQdp5PchdNtYBiuaBwa0az/2GPM/PJbndgRkD7Y6wRCE6nup+xWWpFWOUR/4aC
RyelwA2AJePFOPAsk/76sJ2tEFd2iW0WlW1Zw8rPAvXjxECP3s1Oat/3sBewH9tJ3IfqQlSGsZZ0
5Mpx3OUXW+hU/LoiFFsnvs54TbbaCwVaVotsG7Zp4mJCwmZV7Sp6JUnXjTDTDK6+UZY01Q/RkpRA
iKKzZwpKrplO62RT+5oBGFSQA9AbIT1IvO2/sEt7gvbnwrGWr6S4sji5DZ+NyaT+rMMyrhOLT4no
qGWpM2eb7LFwwmXQGSKrTkASks87fWjLj+gYohHl4Qj4qGhXWlcqIwUdc4ip895+vG5tLCevn+zM
UyNzVzZOEN81GPvuLJ+MkW7DG8r5s+i29b8K+MvNsaTrtnBTNHlf8bHDQwnbXL/noZprRcNZbobZ
NeFP9N4hxpxVv7R22ZlMB24fAPOHRZ0hEXDPavmz8h/nDUJeYjXJ9mJFignOalRRBtkVpwA9a+iK
aJohIQouLNN/DH4U/q+qOAKyLyDSctCuuQpoJzj6//265DgS4oKUmYYguRij/5bxWoy/7EMqWKwr
+5hVLyF+3SfGijLTmYbX88QOhbdtY8pyV7ObUn8bpadrcX9N4uuqAstZXioFxQMGu45cFszzywRd
Xlz0z7kljH/WC1omQSAJYOHLMhndhNX4L++6zqd8/ai1nOFo5BTZlHZ5CiJ/6drHGE1b/QCgng2/
GC9wfRbhB5lUku/ymYSOYNYyHhelcfKLdpjdqmU1LjWW2l4cpWwdvVOeJ5I8wP7prF+7FgZUXtyu
YnacZeCz67Uf0WDEzeJs7406p9dNpNcO3GB51114vGOQFt2cNymsKS9JYrQlFJXp4tSwMiXZnQGL
hhp+EnUNTGCqCRZikO5LJHChxh2f58X5iLTce39VeEIy7vkI4HmWeEy+Ts216mhgz3pUMmvuDA8S
JfPUfIDCiBRhARG7Xg/PjjRA30Jxyl4JWxIYo0JrWzcFCH5ze0yoiN4nNuVoWPuDLj4VpN/8GFZn
/CRRbvywXL4uQ8OVv693vJRiqGhcTrPbu4yu5/tO5zMK6cemCbT/KWOB5J4i0Q5V2+FoMOHP6/Pi
3GKdY0tCzWFgDv5uvC1GjaWXqRvdZ/PPgebKczYi1tPcR7uSxxallhmzQ7G342ZSrmKjWSbXOQOB
WKaMngIsyjjdtuqXOfmjIlCF84wG9p1KnVtBoZk4BcIUVHFpynsgBf4jj9YuNzqkZYM0jPUKCp0w
pXcykZ75iDnozKpIryXxOevTUjI7AONx6x2FC9dYSWDTW3zqRmFJ37BYo71Uy3N0RmXqq9XayNLS
bwP7Om0S8y3FuWq8BPORxzabILg4dIRMAQ3tcDv5nmkaQBkQ+CCEyLL/mFh6X9223bgBl0eNDeYP
EuOfuoDIhF/7Loj6S5Xi6e1TtuW2SzoJm/ahWXsgQNCb25Rlo1FT6NkKu9qsOXqYb+YXprdi26Py
PyXgNXaD/ghp9JzsrOEd//dX46HCFXPymLS1V5cw1xaze5Aml3BX+b4qRMIrRh9wMDHi1TADgTFC
ZCIEKTM0LCWY2XVuUWtoAAD7AzzsxQsS1O6oc7UqB9SPnxLT7BI1Lw6IpBq1Efq/LrSw2CWfDOGD
FuRP6C8Qsqso5BHGuEbZXETera6qRDa6XhBrm8QWdFAJPvUnJtYC2LlbvR2G9aft066bzaZy+sFU
GWKAqG2wiTTPmNXSVBxCatX4gdjBj+xfaQNWyi+qihUFPyym4I91tLrfwdKlvqs+WpfT5c4L8JWO
OzMYGuYfwCiKh8Q580H5jw0ziJQZHE6VyouZlYt4rtBJmKbFGHYkP/kauSf/ETh2GAniVQTERs7C
9wGM6YURkwAUNrlsPCDfSxT+W2gTNSZl7R4KSVHf7Tl+hQO19zxBH/87xJruynFqNJHmP+92Mwbn
W+4yYBhfSfMIxnRQa7zjB1OOlll+50s38qwjBYjylr8UvWl8UvI737F0sCO6TMU8qN+d46XO966y
BFGpKIXOoE4EoK83oBjVRvMdn3UiVJvR/oaJvsdBlj0OurQb1B4+V/si98HAX8O1MIDVwfn5YepD
SbWds9SKK6OOrAVvOR/eVnwKvopAw6R+M01FKMVMcrXp4CA5GTwZCbeBl3sd1pF8vT1UObN6jsby
xzofeNlKZxJiIRhVwJZZL+6NtpltfFfWS8tEUXolskCCsFZjEAh7Jnr6ywB+kUyp0qwNdLXWaoMb
anwXjGXDALYIAiVybRbQT4UM++D0ADoGWb67lPsATLTdrObUd10w871WQfB/8wnDUyYouAdlSjE5
mI0dpynuj+qaqQ8ZG81hbIH+zLGNA2daFXqZgJBTfFYg5RuuZEqR4vg3h4INH+estbtQUQiHLnsp
yKtIk4GHtLCdQDvx07UEWq+fWmPJRyzfMtMei/wY/JBe1hPHV4kzFhY0ZSid3h4Nh2wxOoX21Kzp
gh3eGdcI99/HqAEJHeKYcWJ+8177mdrLZU8Jdm3uH8V5ci4tGyLaA4fbiais1/t5BXBKAm0beO8c
Pp7ZsatAj03RECbdelnwrvVoQ6ts7mc989f6KBD3Ey1D6GecdHcxDhG2H/78vJE5WXc3VUasDQdx
s7DKHPpG8CzPbTFjWSvU3M/gcKLKhcG/7behIJN/heiZ/4TWTwNw+Jh/bm0r7TsaU+bUsi1HrR5w
cYSfMbDvuO4zMVKMm/3Cnlg90e5AuHNFUeGIRs2qvxDUqQU1fK8rPG5D2ctZC9RBBS8X2gwRam1c
oJ/B8ETgtmdxktJXW0MWF+jCBCGvvLFu5x9BF709GJByy4mqTaWYRlgnGXeYwaV/LDQbh5vExYNF
wK88q3avJ5YMXicS5igtId0/W7Lqe6P0zLqSZHyziQtC572t4/H/APLT48XZeYhyBxl9NY7ncCJ/
4JGEo7L9oeepHbDsaXpHsYk+ot3isPmGCtgVvQju5NRJMziJaWXzHT5iIboWWPCuKRMBnBCX14JO
06iBjzO02rePX5x4qDdG8CVxF35FpR0j5TZAI07IDNH2b/adiWNywYBHzqUI9IuVD9ZRwmtkK3m+
5DkdjLzhOJhBm+ZZicqOeOu8D4KqBZACbVQ2+oF0Gy6fDF182cYlA0LECCcnjgpcZWUcuGu2T87Z
FxJVLQiK4U4MvubIavJo0Mo8dbfHsqCPex+9wO79wI/aAdt4Ih69E8OFsftPceoVXNkzbClMRJX1
o7Iefw8t++HJLecJAiiRvGiGZky/YlyReagf/Ykxov10nh3akxJNwS3BsQCLxNQkWysG1WimqbTo
0qXD6wiwTnt2hqc4EGM9sYW3PaoxuAjnoUbU1ctqeCeKrWSTLFapvo4bRojdxuh0ubLLq9zQnzKN
RwMMlXECGyR4YiZephfKvsWndpOPW/JcB2kNnfVBB5u1Zn1I0nG5zcA9iHA07gsr0dDAhNV/rEE0
03+bLm+k97iOGgq1zl32OyHEOiUYIpn0dcz04gAAjcBmhJLZHKggeZY7nuv1MBz8D9pMdrH9lXng
WuapzSm3l2FuAcBLzisHFaeVmtfpP5EwR/BOkHyp3nh0GO9yamdBI8r9vazQbGeVPgi9377y2n+N
2ghsTN3gkcH2rXMPJFTgJG2zCvgfDFH6M/0u72OGSvwmvB9Pqlj4JEKn2RaTQ3q9yXRPblbF5HkU
VTzbSEXL8DDFrBLdTi4EZY4gUaM7waKTqgzem4Vn9HdzVQudPq0ETN1W6zDn3ln2BHjVHdOFiE3c
PukBZ3/6ojkKGuxigcv1Eiq0Bo4trZ9OV78gcoNUK8TmI/wWhcyHBVag1AJ7vN+eHL7zwmcLJRMs
zVhD+B8rRXLlCwnH2FhbCblBvsQKultvbowvBIErmHoUyd3nZ6k+dIOoaJJulvdnnTEOpOqFY1Dr
fKHAO1HwYEPM3B6pU9xl6xoJonrz8Nub9WW50FDOL/f0yQkA3UleCiqMxivMoGrFkNuu9BIr7DCJ
t9r9zqvKKSbR2kk5vPRPewrbrGzIhYkzOexArSmfP9IrHyXOnIHjn8rUUrXr1awxvw9Ffji9MF7l
+wqJglgHYGNvC7FPjS6+qGMC7+X63DbhmLwgx8BPYJDMnAB9Iq8zy7iFHgLNaF9uhm/NwrsVghwl
beKOy1+KVLmiEWMU67pr0C9XenkGq4N1DwdYEQwsfpnT9EbdzfxnVC2oMT+AFOQL5IVSf4fk3dzP
50l4as0YmEPd/xq/Fz+QuAbAdCY97ueXzum6LdP0WtBYtgtzuS07RlhcykaBhPIiyg2c3jLnpfek
emK6FOt/K+GAVN8mq2saUsUHslctHkKc4PYJLpIVUyzQetzLSweG75LMpL9PXo/9ovPb2tZtAjQ6
buq4rahDQoFzR/EoyNkWPxNKjGxbJYcWj9+yLEABqqexszQq+gWYKkUBuV8uW//RnGeBVaJQlMit
99nYEY4MPDSO9D97PnjMJCOz2T3oBO3sJCQ1ybxiFrAMD8cJAkgaJ07/rmdCeU1NF0Msqz1hky8s
4b1PggMoQhmfaEKZoP8pv+rO1xOGb7dyedoIdKr3bsciGkUPut5lAq39PGFRwoeSMoAApgVbUbpI
QkDTZy+dPaz4i5myFR8dn0M/nCt16nc2rbc6o6t2HVRfcbD/q0U/JEKvWbdQ20d7VO0H909dityM
nwJa1yVgKI30S2ZuIv4aEeksrq8K+qtdWCLt7+DLyj6ZY7PpPwQ04ZiaCDbgr/cpQ9UeK8Wd3lHj
/DHrqq00eyAejN4h2fdfQzxIyI51rHYsLBqHDSDI69PrTtZ6Un/eei+t5ZUsZjzvWmRH3vxrprp0
SX42cGLlhXq22kBpRDn48HGHyN4/NaKvRwD4s9YhMMorR4j8Cm2zsxX2yCWqLvBZp9brATY83jMf
L4yDWMfoXtWmIQZIUbulWbpM7DysgzsC009FeyGdHNrWFfuZNKnxbXdQEZNEoNz+i8r0UNRzOSNK
ULgBwEPhTFQ+W7chYTklUlI6iLZ6cZWeDqC3+/dQ13Ur8eMoUXGdu/9G4KUO167X8olSYVN0X7TD
Tx2aloozmOFEKSRk+d5i2OjPqQYXTLHqOEoJhdCF9ljVKOLKoKX7ScHsyMqNllUvb1Zr2/+wT0EX
TSRDoRbwcNVrjPm5/cy22vMne4ch1PONbr3ANbzrqCTzKw7KSgmHEqe/sPzNNa1HYyOHZl0KBY7p
zujljoOPmMGKNfie/Zr2Rr9DvhGOEuxzqD+Dm74ChvKTwWBR4AG1fYPU2iayIniXfnGMNr7H+0hV
4lfOoajBot4WrYesw1ZQG3WwdjcgRFpLcer167f9kuQt2bvgAnKqT8vMsxmrbGZ1eN9lKTiwD41H
kXWg+FjyB8lS7Z9YUYLCoIn3Xpn44cnIaRv0YYVsmofTWQud8i3dSx2iliYsOArKlrVetoJ5QStZ
M8v1+IixB1H3iiBF0WgTL6iT7ANAiERhfLetikoraBYi6QEsJQcUTuoV5A5F1QfKoNG9yZ/oaP2Q
Dosu5DcJ+wlQSRyRoYxMspLQERm3tZPlLUG5bB2aVLyNaIbDDHGrN/Y8zazfXCsZz3fBdweWU1qg
D0k7YJxgYHCKwYGFvVWWWJU+suT5B/vlBI2GN+E+9kHHZHsaeVzKr/fgcV15RFQleDVf91M1T6XK
RMBqEgamkuR0HDPp+ggY6DowiOmLg/hJnreb+zVu/8gkY+PktHGssmSzJvqde3Xoa5zEHEgTxdPk
WJ7zXLJKJQzmdlturifuaXO9n477FxB1jCv6TN5eNjYs9buDidOuMCav2kQDOGtwl+6haHqiDFru
OMMJdjrA4uoZiBaVbZDpwjpP6k0Y9tE2HT5F/HsA+vokO4pRSo5yDyh/O2ri2cnssLb42JxTiJKj
amBFiWhguvZ8ALlXLMb54eVE1gucE931LNUxOF3ZglqA4YNqK9cBte7VLsmvBAILnDMOcO8VGdM+
/v/TIxCaj7FvNp2cLY/BTHiTFqIE6V3RaJ9BUt9zgrBMvcu0K7a7lBsf4UPhLrFf8C3Ex4J8fI9J
+nEaTPKzm2pLpSsIFVeT0NlzbHUsj9ld0CGhjGLj0wXCK1Y5spgBOsx/Hd+DhgQTtMOkPAfnQnN+
P3pgUI5UdsDng2T2T44QRmn6LhCNeRujdo2JlfjFEFqG4cxhnZV/QpKbIB7FSU6v42c5u2Pcmzdi
IcX54f5g+9EkvmnqIb/25ZPVg8qzh1pFo6W3KSsGd5UbcVntxJm/E/Yye7Lckc09lgKgPDQS9gvj
jL53oD5TjrPQvD0CNBLv9P3u5bpSLcblFegoTr8jcOo6qC/fPDfFOxd0HpNWnJg+GWNPUyvIimhf
vS2V8R8nvXXK7XvWl9BKOOm0MDLoFWj3LoPkdNh4biXbNNHm1GJsl+U8yDGmagvYQoxtH35NpyIX
IXpw24jEu+Bl1r87K0tCMIXDi0CS08DthvkJ2QYPmXjtmwimvj1/fByei/D7JbOMcAZfnODGVu0c
8oBqQtsOGE9jmq2SuTVl75cETdUKmPddD25aLztgeY+j2LZ4umbW7D8Q+wlKsr1G8NtefpLCQYDG
vFyJAgJtemVzW6uNhsG7mv5CO1JWoPQzEyrzXVwgWZeG7ht0DlKAX8doZYbkjP4cB8AvskrZ8Ayv
Q483SpnUAkDrNcyfqRopjgqyPcWAnteFQKvVXgFkYKALqLWwBVTfCq55mubhWbZXUtWLninOX7Pr
/gXwMQStt05n0USIPyZ8l7HhbccnUxgTdEdDOMiig8J6dQzl+/KTO61msyPlKHPi/YahbrM7msKD
UaOADawYUtPeKUVNvH6/PhpzuvUcO3SM8e1FfC6+HaNXzPME/YgBdncCGA2d44m9v7wJ4xBQ/iTk
Ct82F6tt8r3p3b+YPwSNYjXluA7y/TH8R97jwefYdqQfJ2GAtJaniq1vzGFh7zToHThBvYJAE35U
8TznMwVEDpWVwLiw5rnc53SzhwyPRYPFqA4pyz7XIlukBk6o5Mfg9NbYfB4Fonm8L6m0K35EYgNf
wAVTkf6sVoHU821oTThPNKFpWmEk4zvCXitXmB2b9/nJHeEZ57wTo5cmwWO0CiNxaiEHmNuTfVaX
RMqprYLiDFC7pKTnYSZ6N05qKV/v3dYmEemtLchHTrPsUok9/pPTbhiBKH6ULi7c5q7O8Z6gDB9Z
f2cY2XX1+B2FH4SpiVXFz+YMyqJX78gAkzOhZksrRp16MySPQPUsMymIs8JnrakPN9rGN4VYv5gh
6QIj9FSfVcehiJ/JrDvtwv2Ge1gdwkTjD8L7GCH/bEcRAbRK2RQkqMLSahDdev4MaVu9yGslQ3uQ
QwCtgj7DRJkKKumZS8I7ijn5QnEJWVo84y7ygK5zj0bs90I8QkSvEwUeene1nbSqzwhFAYxkEHHK
u1Z5d6Gqs6bsffZmVwbq5SkcFBWTjlZMcmK63M7xi+dBb+/pcSdJICO2TO+sGmAKaLzu/ySxCN5x
iGxrqa/NP45XlnjG4woy8l7FAFF6qflKWVmBcQkPmSn3QNU+uKr8tjcsOCbSJ1sVNl/e1/c1WctE
9znTvZfWQ6fDk8cHzXPB1Wk0yytilSltvlM096HBcxxKLAYQpgp5o1Cj08uLNxk84Bi3g0/Qt0mr
EuSQX68U5do199AhfKSQY2etbkcPlDJe+fsTdi0nnQSoF/UkcjxB+PuE2NtYjp/gPsJycxcxQCvM
pNGEy12fLsChURB4bSgGjQHDbHs7h1H3oLuZdXQYJhFN0HSoNLHwjNPrq20huFjSguFmro+O027b
bjda7Me/besMyV3Q3IfnU8Ms/GDJiua7uByMy6nnyQ0ydbDugeFQxO0VvVboz6E4bkqZoIwtrXdH
SdQuDKDSzVY6WUF5nd7/rp96UdTzw29oKJdgljiDCpWPf87a3xYMklX9fVEVLB7kwR0ST1WymP2t
PS/Y8JQPTLoILdf7R3DWE1TzKe44D8bgj6QmNPzLPIn6hIIF1XWDhSMdHeF8eA0Bfv7dRC7UZTGN
aAZucLOts+C72HjMe68haAMgExhVdJWFHetPB7FeG1AvPyu+WZpTeI1HYYWXBen2oWHLxzkJ+jZi
OpvIlI9XGyhYRHh8gpQwANNh5CbZzE8rrq+uzAVRXnsfx+w6qNa/1zGkk8TEoQNlByZNFd2HieNm
xzHbwp3C2SRkhlYnsMaGtsKpKh9rvAjcrV3NiINg2Npa+3+b9lZ5n5xSj2dkjZzPcEWddQd5w6MA
l2TLn2NRC7htwAbsiICC7y6C+/1oTYHjGYSCTU//Wt6Myd1HZNTQE67ZprTikPwuqqv6WxnRKZH0
QbUW4V+3UpSmS2HtZVs4RiV/UAD3Kn2U2idWmFTrnLMP9uwiLR+Jk10bfCQKwxovJjZF8z2comLe
hzjVGD+hD7hbMfz7GnTtLd8jcXnpHIS+9sCj/XGPXb0mtIi14YXUIUq7FZZnqwOKDSqwA1ROpoKo
6SVmQT90v3+5rBFiPBbVU+gf5vwb7suROrMAaOtq0JpKekP3RF5nCUEpsS1EHFtd8yfkkvKzZuZ1
xO0bXVQMS9JDVuB99c3OJ/71GSsEL4nTyw+/w7ZelGV3D+MbC9my/4XFolTtT5EmK7ixGkMQtQZn
aP2v7YXCIkNZUzxxdAeumNnRxpgLWS7lxzcTX2Xcvp/sBiX6voBtsGuNLuaze0AX/56bBtUv9nPB
TAmgwsR1HY1X5iAyBspfmJ1sgUXDK8hBj1zsTsap9XTzxi1TDE6qaEQqP+pUndBU7YtRf/6XQTRQ
FnKni2KuM98ePY9iKK93z+49ygPyWlT56vqng89S7478qCQ+o3rqZ54wEgOM0dXo9UUpmtCZcCU6
UmcepeCMNVdB/CXxvZo8bpYFA0HcASUPgBg3Zl+c5v9GPbL++W6v4QFhSKaPb1r7EdMT66jFi4Yn
vA0bEw3i8+0NYb31LGEfIBp0pwn7ing6JbUV6xGxDkXXje9877Xq9JX4LSJacIn/7Q8YVg9Ee2bM
Q9Jc1UgXQxgfG9yfRLLa4zaoOZRBfGoy37pnYwXE48uGkfxlJaobPVPTW0m5/kTRghfmRDtkXl6G
I5Yufe74sBtXHJfsFsumk+4PO2nWmglkLNNTvrQvDcCtwZj6uz4oPdRZYJcOtcJ9EfjY5jUdp9mI
MzgbDK3xrvmlKFn7t7gbmvl73eOUxVP9SFNoBx33tU1Vbbbme9gS7S29PLr4U8UKQBSVWYXCjNq0
p8HzxJGngO8Eoo3bHaQ/iX9A46cZ83zxWsTy5YwZg0etTbLgGw8eG+UN6Eg9Q6X3wthimydZIMhI
qiAPJj0NTkrIIfoSwbDOU7RbVd2zhI1i5xh8GwzNQa/QqlBOgFBipF+uP4jgun0oZ/xj8Cf+4j2Y
F84JdXpv/WLsGNN3OszpL5WtanOqSfrOwakcqc6GAbi8ISCFNxS8ssr4BlsTKV2Kxc7E+49Zc8+4
iHWDfwi+45ljUJ0hvdodhf4II1PK6KwAPxgVDStmdfZ5D3uStxXf39cbUisSiIjDz92bId2g1b6r
Z6ao8l0TIw8Klnb8CqBCkvdu9/0Mem7DTTW//pdrHPimZhCIbvG9l6M2MuXRqD/tUE7azsgrhuP7
8HwVfUTtDRa2j/j5/JrMphOUT2mEzEeU31Jqq4BhIT8pI3CnP79lzchyIgsBc2IESlKUjNP7foZH
FROJfOIwpvJHOeuUJA7d/p/WJpd28bDGb2+Hz4Big8Eo7SiwSuascKuXYVRxKaU796lYbZb2w69i
ppG/PI/JOTNzxGDZyIKnnAUpYNS3URgCg48CKaKMA6GzJv4Cgq6ytkg4lBvLewiG7ZzfKDOtu+6v
itaP3mB/UhI5Qg8Nm4C9UOOPmjdAZatBWj+eTvDSQZUleUEwK6Kg+0de+XTQ+madLRECTdKit28I
Wt0/460Vsnt6J6tNJG0hkoarCUxFllKcGyfR2VlUbpkQ3X7p2Ex/fW7YRRG/7iBM4MzBErfJWGas
EVSKCRGnEWqjfCJlOmJpqmUaE0OMXJBPHhIpJDTALkeOWir3rrH1isTvbRsRpnsHae0sQY+dsUz9
DbXlg/rn430l+nfupcntM4vOqEAgJyTGWXpppdjlBja6cFtE8Td0vMuKh7Bz8pzg7cQTuEozmE9n
4oDiH0zddDwa2eU38uNTjiK70JkWmOo6e6TWgTG99HqJfB44ixZKihrSLfT7T9LfQ871Q2AP7bfd
FTk4gcIpykWNdqi3rG8HJ579hTqd21pVdzVjCgRXOMK9mRaDDP/QrhuPbyJ58IPpKcOliKn4O7Ue
6E+y8s+11aE/C+1bRaCQyDI5U66KqJUFamihraadbw1CpuQB44ReWdiFxt+8s4Mqb+RWl5B4zTuO
ILjtSaMyCRcju9Ps+ptJbSN2jGdFFH435kLlQs770MoNY8Il25SUJeFqcHG4XWEI7ryo/DjjY5Wl
//p9vr3AqbVxjjcpx1pl65sot9GpYflFRliu/FagdMskshqvo1cbcZ7dbzssegANr5g1mw/zN46/
wb+3QuTHWFN4h8F5vre/KnaXyut1/iTsdeluk5gNVMXaSUZ2ZVmmo2vYhZH6EjJGHONMtl8yg/oM
zBiDOp/u+xND9817J6UOiWWW1Ioykqr6cgzowwV13nYAr1mELWj9+JbjDMCQE1zR1aOUlRussrRJ
6PRgWLAdrH5c7bv5MeZwR7ZHyQo0nL3KVJ/WqPKZVS1a4VYXLgMuE0enXIpubcIgYWmpIGQ6rJiQ
BfRE5DDj+H5GLaCiDforyfwWpwAm3iy/8Tal4VbmYXy4rttpmoPnn7SsOVSbXkwsOYyY5wib0uuh
3Bg4kU8DK1z0etYTicVSGf9O2+gnnMUmg0EOeJmWotCbiSZSfhq34Kq49SpFzbcDuZIL6JZwlrFo
upyp9dfMTYDwesDZMujocYPz+HCNrjiKHEwJeJy5L/hr7+5bDt3hkwWLShv1HgGr1kfOw4TNKnrF
r4PiATQ+/sBc4aVBIPHzCjGaCocoKmZJan2PvMKPv5MJVQbZ4JBr9kiMSGiiYEK4vymndZLRMFgV
2go6+PgzI6LCQs/xg0XHVDoyyL8W2OKWVBprueGKFD6bPHUTXL1kPidVDnksE0vqWyoZLHfsS00h
mCZtYzD+jqmDrhQKgf0ltiFM4defKczXmdo9i3BPDCa7zj5Hrc9iupnB1le7/cDd4pZSDEVgwk7k
1XtfyzG+wvm9PNpH+61J9UGle/jdbOhAV97RlxJozFA9wyQP1wzTnD1Ha6GAKVhVUoD4tqOTMsGD
U0fo5WWcuipIaj+uLpjbVf032BS8YX8Ku89+X3hXNZxleXJds39o5AEAPf2GolQv4nF9Xa3rMpxE
FrF24YaWQxO+cXbXbnA+5y/gGnHG/GFqC2iwk4H+tWsQXKT0mO4F/qAEYhXAzthpAETYplN9Lz6F
WuEz1BMhkvwX2Nc8iM3/QQc9x1vosk4fKqWMQbsVxj3TENiHh3i9L9IZg55xRPsJd/nmCZ+pBlpM
BbYNHlm//t+6IJpoTg5+lgggluhN/YhzdSXKOEn+scIVPxA+W5pdPtjpi3odTNmpPD0WVT+YcC69
uywVa52NbzV14HLpQ/lF0hx5ciPZaxyXdoKo0xFPiooaKoDea2tq/rkxUsjSg7yjz7hdEfoGrZ/Q
ODgSJw93L0tbY590BsO3qD1iUticUKR6f4sMIhIVbTV7b0mQtzi3sK8Z8pXcPj7tTC/f99/CRuYl
xTFcU0RkwJSMkFfGi1L36gw44l0LtrjGrQYUuEtV64p3TuBZzjEWK+/jkaUi3ZjRVcy02Jrmnbnl
pPSocDK9gO8684JSMGlW/f3rCITscbmFY/4EZJ0XOamFqiN9NGe+IpmauCTmfXdytlr5YArP8f+Z
toqGjCbR+t+Vm5ejAX8JlXpqiun+KNgpH95ThWR9a/DC0mggOM2V/CXnJZwB/nPXRdtcasLrTLO5
19mC2cXCejs24Wbij3ozZHOZ/Wsd1QnCxM9i3DS+0xjMei8hChgAGo2I5Pm3YXXN04bkumQUWSal
aW3dKAi3fsUbs+8Gyncey4ZR2Ep6rv7xeYjwGKMgg0PPzNfyx9rBaDd1AF/BpUAmcCCUC2yNTVJ7
t+kSN4K3amko+jBkgqo8r9hb6ZxUYdiCRspP+PKTfDUNwN5SGH909uLW2155TwFC+o0T8cbYOcIA
C/cGIjmPjuhro0RUHGSaOkpz2d0VYfQbDyzuiqqPQxw2j0w2EiGlE/QQaouPmD8BsJDx3vzJFTlY
KK//YdxtNOysueH8CXPIKmfsL4yEjOeW4jzNeCaSrTLlrzEUK8SLUsMpirDr2SoYwyrJuZpjP+UL
ADtQZZyMl1sbn3Yr0ZfZF4dc96BhM6e5tKYhVZkG7i1EbpUV6CTIzZB6ixksVDLIn5QBrbwdcQXD
oWmP1avdYVI7qM97bzAfX8BIvU/CxksJrk70clPzJgFGCJkNMRZUZ0kdxv9d5o2iEM0FdmWUjwhr
MiZe/3FS7n7TmggQp+1q3e9nXsRsWg2GnEA++uOmc5oZtmklLMOMFMxuwPl3D2T4xkchoKFHRnF2
R8tygng8hiS2BlhZ6qIX9rsZLV5s2NTSmDH0AjwvG9ghtq+Rog18Q+0UpJ6R+XzVwqgvjW1omJVm
XLWW5OLwOusWQxvLF4MW9gIKVc9dMVGjYWZs9YUWpTiDdD/5bsjllVMwz/BIn6iTqLvNbmJ/W4KM
rY/keo64MVQ5Wj/Ze8R0GYDFYG56WeHAU4/aBKrk7QUPkL6QLquhpEKP0PyTyDqUjqjVIzHGpzMx
DCFXGPYY1hNqfxcQHhW6s2g1/Y0XX8MlKN4PA7RLrFb4sto0brza29RRGNLQnbbI+ZtqWY18i5iQ
ZG3fhsuMFJEbDnJ8D061F/o0ghPolZl5sFNRlXu2GfMt0zfqDgIObN0qE6ieNs145nt72FmPzalk
ujGQ2ETAbfS+YB8+DwhDhl6yERDUsez6e92NuvljaUn8uU9p4/peQGDfmMHZV2wBZDBkUDyFVDYt
vUfVkWlmMGAbX9vSb1vWgOMrpGqoPz9r1wTRXVNLzU8piE1LNcvOadoQE1MyWALtZ5wgZSZiEwej
wgqQD3EOnWlSUu8Cl7bg5G83E1A/DBg1EXdOs27693z+LVsdmkRn8bryuoiKpPDdm34TmX3TSVKT
6OiZq5KV59naw8Uol0fsrmw77FHI9H7kl4/WuRCDrgAfoE1VU2UMmGcbnyyNJezs9exBPx1rb+Z1
Zz4nKEoAB9xMpkEZPgg34yZAlPNBZzwezwTNjQdBPsTkmyy12m1T1wbsqdE3VXmPuxg0n/kHl4Ln
XFylIrBxQ85u1jrH3YuJRQG4QHHCAOk6UfMKl7RPLWCvUFypdthNZcWFJjb9c8MyTAjr0RYnmB1k
ZKj6qJIPLat1aodBJKX3FjpR6iq3VUNytq/GiOgt8Kccj8Fu+G6CbaLeTvxO6ajuYqNQkQUV40EF
sqt6CwTg4V607P5daTl/UnqmxjHH6GLQGiIN6R684KcW5FlRpT/JKPkyGMYSyxmuB7RKjTfD2fJi
/PAEiBqptmPcfExazRZHkVmY7/ncStnhoT8h8RiaoBddkMC+wcekq1sXbYmOVQIDYAgFXW8wH4Cu
zkvlCnbWyYiHyMEmUxTlICi5JZZPM3Ju3i0QEn7FaG3B0hWes6AyiED3xfT2W9b6yX8Ve9Pj+mjx
OECVXeoPTDifi6tC6N41EjyB+HidnQV4pfCmiSZbzXRR4pePhZCRPzA5HJoncA+0DscjqGoS0GK+
rTOlksMMTpIPrq0Hwiz0+sQsA89t+EL34/QMr3PE2COkJ8xLl2+loxVvZMwcYQv4JuY13YzTq5Zp
9vhn39tad02CK7a/CWeYYQFZZ0O2na1ze+xiuoXfoEoR3XT31MtDo2rgOunErC5inrQdDs9Fm3sT
9GMkGw45d2TDn0x81Oetm4nGatYygJ84VWsoE1zc+zq4b8xyI37zdckwLE9EX1n4yPlydQiN9/pm
xe62kiInu0s9IOi+UVuqlq4gSLretOZFO/ypbLfN8R+9RjBSBKWuixU9L/Tj/HmguJeYlQ5Ym+V+
4O78ek7f7HLmuM/hGfiWAlBZXC4zf8ejnjw4tSMoaiw82pVhxwXH8dDrzO6vYj/OFqnD5nOppTRc
IRf427HJpfjEQi3lLocl2KNzz4cwMi/4RvMPlwN4z/yEgSeGm1KGmPmN9mG50NQS2JDFGvwqHOyD
+IAwXPYiNzLHZJ9AVIUtXqOOsCEBLQIZ9+v15EilWTWRMAWeYWqPZN+FIsujD1qdt+csNVQL0sAx
6lHsacxLBj661nwRvep5B6oqRDvW0hzBuk47PqTC8SZzuq5FZQa2ChLdjHi1a0ACia6aZVIc/qcg
zzHpkNkb3L0Ar5qYmADNqsBDr819Lzw4EsdiC7ZhrgJ+sjIbrSVmjzfUd30bQOxBDWOsYgfAb+Ps
A2qGgd/MxNMUX2od5h7hgYHgrZD6z6YIEwOm29b3Lrz6CLMsbjCwIuiJjJOvIjTVXyYjfDHUaiPE
Mjd2qHJZ6A6QFhKVmYIQQEcrw872wNBMh1lxUx3+HddPK519fD5zFgxBdJ53B0FG6olnslOXiRpU
GHPENSuzrcijzFnZGvpFGa9lESE05brrK9cuZnNleHBkFL4TTsslObOKg9gXNWs05wZeo9F7UOBR
eljyNVkJbNw7cZ2N/dzj2lUkDwDBxOt0E063kV/CYHDy7UrZHayjU6fkm46fnb6XyP0AyIBQY4JJ
L4vFyQQ8vLt38ChIL0WGcqFnaRO9vq/mNAt/U+MW1Ryhk4i0UFTgbj0rDT8UqlIDMZngCt3uZXjq
oKrPa2tSbepbYYpIuLn/jvEDRY5fITbm0Phr0KYUKKvc50rPq2a867fjoCrVsJ1/pOkEtKUqhwmJ
eSdw6T6kKUo63jE04QaeOq2+jdSCruRvLnYokmHtv9n93oCRHbknhxGG65o213H5OO3a0e+wBYVm
hh7Dzb/Er2s/1/y982H6icJZLuupEcGtXmSNbLz+dff1e5H3yMbza/KdlO0kJJgjfy5sa7eg1mbN
UBZGk+vUNR7k7wXduBVmZAr5DzeUpOKLCftWkt9oHvrEHk1Y4qiBYm1ncbb/ysmKrUHFVXL8qQSc
7A2hSvUEDzuVWPXnPgZwdXpVbonSw9z8KWw350Rwb54dLDsGZzpu2BJ2X1SFkEWYr8QQto3JdAtP
gH4X4nIQ3fVIhcwX51SslvJT+3Ko6bR8bWNasb8EqYtFaSu9cm9e2xAOmkiRZmXSNlaKnxmaRrKs
sELdUgPqwePIDB60eIqJB6ffAYESL8d6ul5pnYkAiCvx+ScNwfkYVKxdw71rKlJkk9prcAKUjHhT
w7Y8V01yqw2Xbgau7faQDC0zmiPj3RkDtGcaIFinDoFn1xR0y+fuekoYoVVQMApk1n/aq6SFveSu
Fv0gvWAqAcPgsLwQGDaHg9fzRHI1YECkGR1mTjNOQ8SiEMBv1HUZNBuC9xIfpOqrrR4dUtaR00Uh
xLOEvAZXOUiI/q/Eb8YSTzUkSPPMR1SvOD4W9yhnS1SP3fEc48l3/qn8na58jEW/CFVClLDl6gHq
inpS+3wvbWilF6M3pi/Tcg3Zzei5sf06r+UyES20PfurFzohXXgqHjvnD0hV1h+WWlYq1c7WYWaW
B2MpBCLAiwWNZL4aekj31zRvQj/O2apzpCZ8BQSG2CtJ/yCIVtiTD0P/r2xmGi3xfS5vvWQi4r1Y
DpirZAApEB6bQV8I+XlfoLBf69MEAXiO9qfKNy3bn+sQVnczbHo8ZKmpjWG5LWDDTejncaPrWCE2
kSYDnUYV4vb5klRWt7WaplFgvR2t4QNbCvzteR9DbZC4aMEJB6vqZO9XaTMkUIFO04/SiKx529Xv
w3siIlFTj0dDtH8bOD5nRw4EjPQqxQXPnErIthqC0gJ+upQ+GnzHg2O2oRbdUamHTES/eyuvbvVu
IdzVjPLC+pfCE+GueFis5J4qmHNShyroWWDneOfcK1ZF+gt/Ma9ONhuhJaL4un3JUFSFv2eekMCp
8ClTATCsGy3+zDQhWiRg47xFtKXIMYe/F77EUceOtyY346hg7Y6mAoSM4ta5RIsX7uDxgyyGSTzx
bfRcvawQsdvo2eM6XoUGJMXV/8poKlBz/nP6p0ylhgn/eTGnhvHxRI2U9Ujgbw3aAYfxP6q/KR/V
0z/TR1rlvQ93muyLg0k3d2sdOXy3ZyO8f2y1GZWiR6YfOrGe8YFs1Hx8F3bOqrtHz6M+0OG09Obc
UYQZ1dEo6aPw090Dt1UYAzOMTSp2ywMdjAdDBytUuqjOoRZhOscGsb5Vd8CXRj3vQMrioMkDQer+
MfEKmoejrO/1odontgRh26JY1nalAFvJfifJ+UAXbpXa9tUDxlGNVfJK9FDIqhehEx5CuXRjzSsV
81N8wgVnpNuOquc+0LtrqkU2l9JLQnU76xeyT4TUIqFXxYr8G9uqVaxj5eyWXkRkDDs0s8tp46B4
csv25BALgKQJa31mu1S3kRRyfUTTRs9KTnIAZzrU48RxX/WKUB0GMEY3Rj2JyftlKm35rx+uJrM6
hH2xUnoC3Xf9Gy7Kbv6KBbW3f5srm4HmgXsNW+FWZh4HdqY7DKvQK1C5DltWHTfRZmaDekZGbKeX
MrEG7bgUf7LO+WQ5RIsvi9GVwPOJyspU59Tmlls7zD936WVJ41SVZTLGzu4wU+gWG4+TsMnKUm7Q
jMiclqKW59U2OwS+5sgebQ8jRUjJuoMQVh4DAJba3tfthMbVcbdP4K0UOqeZAN7xrSE3Jt01obiY
pVGHsvSbQRmwYzRUsXJKSink+CxYDAY8Xj5QvjTUVDMaVowE5NTf3EJuV+4ny2XbWEhVcPAOsEz3
XLt5WFXlm1RsX+rMmMmReCMfMsmX3nV39qLfl74LjWrIGRJG0KX7u4PppjP/bcTdFZfHoY6C20sM
Np0Tv5p5pfPdGSf3h2w6+kZAqxxCCcDMErWxxmnBCcTSOBK0IsiEm0urwGU6FOJDS0Tbnp1aCP1C
6O/11I4z/cS0iH1nuh7Qhs1WHb3PCfb9VY9Duur+R/BuDaEiLf4zMfacCx7gIVece9CNYoADc2Nu
jp7VLQ8E1z0YloU1LblB1n/PXXkhG+ptd39sqkaBiSB6gs3lB1mDsP7i+D1s/Vc84ggTeBYxgDw1
skUI+HjE6LfGjej89NLGJ8UZWUYKX7DyyjSsOgs3KUopetnj6kkMw4vbT/CfWvXzWdivY+hb05YE
TIAC/7Rm2qWiEP1cb6BKbKiLJWpJxRQD6rfl7AEp8+BsBG0lFavciGYJY6L7HQq9Lc1Az+H2VlYO
qxRvYuAr+O19qinbqy+1AamV/b1pjyfmstX/neZvb2tXHA/2e1MQ6R2RVUAb10q/2GEEdkeMQ3ua
+8bdHPM6LjZJ18wDNQEXD0R0o/LebXHQ+vJsJHgCYLur7paSp3RHKiBVHloMVtFQeYWFDSkpma6o
HD+1GnPOKyRwc+fnelWJYPfL5QJUuYkh0R+xRZ5ZsLaXizIBE7jICyMOtoQ8SlHq4imU8tJdh3Ej
h2v+I/eWskKwKZvmGJyVnco2KO8xcLhrCRfkbZTBDNXEeMa5sdwCK9XqGtR8g3O97YAGTh53RHLB
Swl2/j5N6u/YiAKr3hQNG3ZIhdEwGlJfSbLxwc8uSHEL55DoEKoUuwi1xYdVKZb+CR/yM5SXg1Bl
RRx56MTtnQoZVAEtHHQOX5nYQmMDY41P09oTdJGC56ieTJdhheLEqP+LHIc1wmaQFlU0omlKhOp7
KON/aqt8d/V2mKvaaWjCtoO3Zx7hCo13M5dGsRtlsTWrfkwd0WUi7bG1c7xywBWMEBhcmKtJwOqg
NRFPFtUU/F9p1DGZ1mz/iSR0Ib8tVQWXDBh81RqNBPKZU69/pAuIUC4bSW82UXMW1jaMpag1PJ1S
DC+zWLqEmdFsKp7vqEpPfjcuS5jOxR66uQMHd4eebhQRDKENfX13gvibrdLXwxEAO6vbcEgBN2RL
zyQO8LNsh2s53wkYKRB3ro3bTS8h19FzNRsFP9HVNmgXeSgxzl+F2Ca8T0+I7TTr7xCnPh+mYVt+
Pyjh/xYujN3MxQS5Lr1oGQR2vDf7zDL9v05c6M7yo0jjAQcCxd8Y3sYfOfEOIXS77du1A4DM3y8s
qqaEByCcPWahWpBjK+V5aPgjHbMtjMpJzqG0/qoTyMxcXxUcdoMKf4xJjEpHOzLxKlxn6j6A5odg
cEbMp7zbKz4GappKmluDV+R4yO+GCNxUAUJACQPxk4LlC9UDi40jP406MV8UajSVTibtTXxoPTUV
9rN4vlLTk4k/d6qMXXq9FZf6vWP1NAqQcOhsDwwuC6OtDlOlNiFAsesgQuqipQ/2miaYfH1B9gyU
0MzTRPji9wO6cCgxDTp6LpFziJjgOfzIp4ayFYtXpxDR7b7HLnuVTM5LeOcKs4mtTvhkDTyZFkaR
Ur+oiRoh0LZ6hed/w6CRQfq8KHkJENemnqBSlykdGHq1zBw3Hnv1XqiERfH3SWICQ77tiG8JVhBn
68BiTYwdwncWbXcrGqrsDQpOI2fyCsNIBXqBZbM36nFDj7NCGR4EQrckaik+VUb4roNTMLEeKvc8
tbf8t1zpaenTQCxQRKunMqgW9g42YqsnpsbYOT8e7PViIKFswb4XbKDTOzEPegzxarUhr5EPtZGZ
BpzbSCBhMxNhN14TmA3w7j7DuyeEHA35KV1cEQGug9IEhsrsxkbqJ1Ee1LeZLZ8FjiN4Hx5OUof9
S5ISKirSmKfmgYPMRAxC+3g5pZnEE2FxLjhgLIAsPBg4aQR3tg6tnE33KqP8d/KB2HY16M5Jfzz0
1lbEON9S+/w4uQWk0wzWGmpBZ1fSSbc3ZaEmv+/fYgPwIA90UHmftQI8RAw0D+f0CxDp5Qbw+qxo
gxQ3sL1mKr4RMD+dgLcAtLVDVGtiVIOUzhVxx6b6qR5WgBer8ffZZPE63+HyZG8MCBDfZZMRyEQR
OQb3hEjAQchne5RbD1krZkEI9mX4IUwJzgQi2wxv3v2sGRxpUck1M7986/XLH3brvYfLh4NytLWW
FYPlwxpXY0Te77M2ojwAHmrcuE+xVaodJnjW7KKXC7cqSe+69+XzaFw2+l2jhEUBG/CvepF63HYl
Ryt1YgG1ybCMB6xS/CcGtmVnUnIJDsAv5OVu4b8kQx73gTIxKSjps6NSu3CHc6aNysRx5hcep8pZ
ROABegojW/tYqpNPXMiIaH3LmekGfxL0RMt35p7gwIALgw4CCDFA2VgQuvJd9pttj96XR02eIJt6
8mVODlqj5AQ/i6DWI9u/N6waFdsMwhh4+LSzs/mt9CBlg/i1vAyi8R1IHYQDX3s+CuKBV8x73He3
Z01OgWgr9x3emjUKx8knVNft8E+UcSzXfiqRlMNF3pd9ep1WtOEDuf3GaMI4GtICv36y1Ccr8hY0
MOut4UkbdCk04GLTYk9VTVGiBojNHxauZhpjjFJSBkTajvlrv54DooWrPbsukcOWyHz65MOmCwQ/
O7maBIrUn9+yU2novzogNXmhHNIWe56E/tHr+e+RuUNSLbrkn+ekIkyhQBJj3Z1EwGd3+ATimBkl
a2dswp3XLzsboWTsethE2PMXM5cY0SdgEqNqMiflziOwYAsVi8db88sAbdBoXMx4iKJGd4v3ffx+
/NP+6BYZAzWzPLPcE/uMyeoW/boiYNo7KTQ8d+sLvfgq8M4IStKcKTDI3SM6PL6JMouZMcYBTH5O
VcPKUurIcdfKhnXnOJnjoAisII/tHopsArMIvu5UA3poX6gazAaTc4UTwu0ER0hHbmhunQVjKIyF
XDnT7RbkZIWC9wa1FezPFPUmdkwz5Dd/xy4+weNrcOdQZsIuagxLw6mKWZULAPvQrdmzUrzZKf/F
FieHNFKet84JogDP1PdsfAhe0HisDyNk3dmbguBreZRkL7+4HdTfJ+9dxSs4EcXmmfKmMQKKNvfg
PQ0FAKgoe96DtrhDpx7MTgdWDjQc6P+TbfPwG9uswISgDCIrMNpHbEbXDsQ/GKaOyD9jkTEkma/e
E0Ap18CkFXY204u0qXv/Z9O+O37lHCnfbaNJkK3Qx3fVWn7fSR5WZlKUIjrJ8TVWd5vEx2caffGY
J408mTC/SgkhfUjuWC+sqkxPJoAxVAQQnw5vXAb5rZV+Sq/b7z8AFzRVidWbukFZJtZgZ6ba4xqd
bMX9dfw3XmfZMJ7albaFIj0JW7ytCgFn56jE0R2cX+oWwmdg+gfpba9UJd/yuesNRbxzZvg8MGZ0
BKCvBPS8WphTvUc1YeCbVLzM9X7HVRzZW0chrSlbcgIlxePBE0QxtrWOhrKfu5EkPYgLKkKB0Yf2
5rZQrTybIuFWfG3tJBfltLUDxdUK8FR1PdsxQ70WA804GDW9ucJz0D4jh/3kmZHupnQ8z7629RWZ
TsjdjnVMHY5LKgUrqWRFckVdrAFciKYgWXIJ5kM+28vjVwxclIKvP1ritFCrVX0dCxS6elaEE8Z8
zEaUwgb7rszqbi4Ng0wloxcuS9BKdUbSJ6GSNBEtZz+Ojs6DL7CEWWYBOCSDq6L5wW5Ms0jM5hnk
HVihTw4O5ELfN4CfWNVgXneS5/rGit64ToYaBY3cy5mqoIFCLOcTSkA7I8R6hj7kf9iPisdXKKbB
Nc8F5dJGgimgk3F0EfjNor2g7OF2LpzGosKvLXSGVmCLcF55dfHNt1/Ca7pLl4O4g1kNYIvXDNM2
mKGVoJrRdZ+i32tyc11Bx56G6z/n1G4kmjvj7asthrBtf2o04VUjBCXNoeGNUd9fMbkRDO4swiqs
E4MijV/aWoV2mqpAxf8KDdnVs+TmMsXbh2w/yhevC4ohP3nHonOEzgHO0cCc8n0zlUWDzVGHsv0f
QEaCgHO3AXPQbjFASUiOY0J8taIkbEhGLLBtESXDOpTh/O9+AeS/Hue+Nh1Ix8dcQ1wS8GLxkybP
prfLAUfT0GxGWvX8grkqHagalmdnnybjAGpX1PJ7c2wu6M9PfyxtqwoE21ziQVyzG4aM7AH8svli
yXnucZQ2DO6A18ojbB0VBp3htSYRswrbzt7rDSG80bjucw+Fxf1UcxYip9V8TpaZtn7uHhKz/VAN
rNuBMBqRAaPZPgu2SWSfAUeQJozO/rdTrjrdACDO7V2tjZ2teekWlZJWRwNtH4ao+7j6X1HdRFd/
icB20s+YHAFsllVNN+UEzTml1IyFb8OB+JYcTkRSwXPuWl3pjVw7mNPjixtQ3Nr/bnDp1GRD1u/I
R6Ze7DvFVk6nVpQ+kDiSQtFrujmFnZoJ9w5F/UdJ+PO5cjK4ZqasFz1PITAl+xEobLx011oiF2K8
6Z8/S6a3iOgb2pnaXiHl7yB3Ln2cDBxForaHGdNjgCOG7scnLloV8rGGucyp3ruvdNMV63IOP/ji
hv2nicO27iWVu9nze+APnTz6npvGxbnCQuxD8ovMlsKCasnJmDpux8IiMp4yjxABiGFnCyXE6cSU
aY9B+XC1jpBVGvoakAjQIvWeQNI6dWjelYtg7MzB9p4mRQni5E0BZLGbJZqbqiLGByqz8AXSYswU
xBlKsKp6NLLLzJG2RimJdU6wb907MHSzzaNPqRqGcWcY0UJgbSnVtT6meCCjOTRXBfrN03dQVQI3
t4QIllh6kticX84wS5+DV7kF1EpEYNdjequP/c5kZ3x8wXltWnvNSmPFJ2m0tQf7bfMvzzwR7kaN
bwry3FZdYhJLKXDoY/EgbM7XO4QJfYGSgyj/0qxUIB5By0ykSj/rTWmCtXVtbCpRw+uN7waKaDmq
q/K9+F9/X4bTXZ0tgjUbJll7e4wjIpzLxRyzFE2bc8C/COQXUKi4DOHUWloxCGOlIuWiM/wbwtst
sQhVTYLjjLFbPEbg+hgKRLFNaY+BbqV+/8bCqhXCGA7vB2sh/biSzOiaAoEVRwJJu/E7PuMof/Sk
NQ7G1/wxbiQPYegHNwLYERDTBZ2Uq7RQIdAudRRPvyTzklQSW+SAay9xkvPhdKrkjJW9IKB0Hai/
OYyKdc91qWKaBVU7rHW8iWVQL+Mrvu1t/nSBUYfdaLPSveDRZW+e4NNRyGfo4nRwUHO5SUvlQnIu
XpWMfKNsTo9ypRTq2tMIvz9ZyEIAejjFM/I/C/klhPzdhnJv7y2gW/rnIR71scEu2CuRrZKeFEF4
zz7pwptTuq6aC/4521BApopKXBKnpNjru76FC8CbkTkR9kARD9kswp6RPHL8jErfR1UyECAACZeh
nBy0ttBfmVD+KofKplcJZ7+D5VjJKxkSWB0TqVSKXGEL4MMQka4fAY4sIz9M2699LH0nfrVBRJSO
mAAwKdymkqmIlSWY1V7os2QTaE7BUmDGiCYjty6BDMGh7Y35cRALMJ78kNrZRNQTwddowDfbhN6X
d7UrcH1PQgaWIVTBTid3xS7wM2ICUSbxH4LtIGeJ2pLsYHQM3BFuqH2pF2XDW7+YtFpu9LOg6KHl
jkqyMJxCDpA52P4so/Uc+3OhqbKYhwkMn0m3SCc9KXAIu4TeKCQr5+4VoW2EBfaYi0l0Ctva/rn4
beBh8Jp3j4niFWkC3MS+oyuwdZBekYprmB1/jUV8R0/PtrwGfzJffo15iV+axIfhcKBn0EjuzU/L
zTopQbsfIvvBEEAJxDdUpgPAU/DZrPT/d4v6GBJlHjSxjU57DNQ5VEN7+m0XzY5XpEbDo//1EVAn
LSkQyjym5crFvSXv8sapejXtV7lldIR5tBJ+WXtonTWVI/5+FihEnNNpOOglFJnYwurMew3ONzf/
nPFYIeEqPZ1YOM6f6E91tNAabtMchdQr71br/qfIAMJPBE5KXnhT9vL8PRha+AEn5IshD0q91yaF
Fv0Z5lRtm4ncHgt2zM/DtBj7DzxIZkbl6HfOKpCb2pobaKd15vKA+HuuRe5P9S5gQaBZj8e8ba4q
Nkcmrr2W5u3C1Op2eSGv1lUubQqN9IAuFtxBECQomRTpB66AaWcBbFUAbSdcJM0Dq64wMpa08MtU
Hr/IevAqw3tK+04JuCEH04sgdC6yQ0FaFte6C/Acw3fjLQ8P226Mkr2hNuFtW+ulAENcXAIG70eq
0WVazWNAcQZ8e6wpgGDfnnOi4xL9DPAdwRu/ePL8xmuwr4IV74S4r2i8h9cNjOrR4NCvORUUmvSq
ZWDUllkifEQPrNHX1Ifkd7isO4Glnx10ruMrk+IsiotURMh+6caeqU/1ZxVSLjdW2vV3FqkCEs0l
xYqpncG7yGUaowsMbDdnUAo1BlvHHACdEnIszaTCfNutxtS+Y7vH40/GE+OCw2pf9Su2h0O4eRaH
HI/m3FyYxut5CV1N/w7dqkBzaj9C3vd5LIQOAOKO2BpRP/If06EiSsnMhYc5SN68H3DQuPXj7E/a
Yg0c3U4TZepQzOllnu/7UhIcG9DAHtBxfCEYuMkjiSoOKDhj1WQHJwFDPsNRSD4MnBLV/EjoBm9z
F3xpQbtks+j1VFTUOtQUyQUZXpT1CVX3tU80O6LiXGpFRriYewrvdfwsMJc9HI2U4ABWCLLRBJSM
D0ARbYiH0e61370/rnta9ngRKLGMZ87iqBVZtworoZMpdtU0t9/nS6FwirRNz1ZGfcbRVOAYBMCX
Yb/Z6Ue+9V2IbU4DWhi+FqcMFB9zfuflzma9edzhyO42lkkcXpdUnk72uP+VhqectD9PjIanbkQJ
NVdbmMT4p8roFTTKRKwq+WnWslG8KkRmGvyCYvVNtWazEW3As+zJ0amhAkENlBOrJtn7ioeDccBe
eLYL+Hn2Y2xpwwAlsbWpnewxXdSB2rdnMBDX6OZTpxp30+bFGRWeYo2PdpXnAqswInb4ivf/K5IS
zGe50fQvXywiwlBFp/v4M5YKhqowi1pez9vZ8FIoXn4pnHhi4IgqxX+na/P3mVjfDX0HpkjSlSjb
VxSqqPsHNmRoTrN+xBs+PpLbY+coavqFQagztQHpspnXgEio4pK47k3jU9C2v8zdY8aMwM6o1dt4
D8mgazNHiC7UGgHPaiMRMuH/+X92Ck8rLKshcKPAczy2Cr7k44UUfrV01LnkKMNerCSNTGsox875
8oFQi3o++KvTqg1kD7tzLhtR2E0ut7frTahV5QuSlMxObeOukBK/0ulBAmiO7DERaArICXExeakz
PQJNxFuZgpa6/VKI3AEgImSHEyvH9XNQqwBO0fIaaQ7RBmt5+mxO+sYn5d6FTuPg3Xzv+k8xOQ47
ReW8L+hMStT+d85PmESMZ9i9U9hpMy6eE38lOvlvm2Lks4t2Dn+zGQKBELH1JOU49N5L7jppVzXL
GFlk3NWB9Rt1LGI1qU3VYNuaFmQawMZf+yAEDloF8wgvoD3u4oEkVb5EIhgCN5+0YJ1te0efrKcy
JIWNYrL8o3RufwA/MiX9dSGuQqOnwfCJOPkwPer69BjZMQ8lfzib56VwGlz6Crh/gvHVNTM79tPx
oWCK96AlxEhWIrKcqKfCyeJnELMq/Ddb05CrlJC+etXTddbRGOJJojgSXoNgQLKXmaIf5lK5y6u1
9WdaTndQUWhogBPzkCA/TT3LkmyFa37nIfSHp5wL3kkjTzdFo+2lpZ9W1MF3FejK3kjFMzcb/qK8
vzilmnCX6prXK+VS9cvgECdLI6h+r+AAI54jydYx9X6vCinsuaS7lClf4ODGxuw0AJR9k7KXytzw
a6HbEVrB7YACZJ4TMD9fRTUagJSmiVuGXIlcPDC/OSUzxrecJih2ziMf4P5HkOXzzjR0YARmNq9h
Zc6h1BRj8njJJTjtMRR5QaA3m9x0bg35GTA1ecoH3HR3VSYISII7+xOHvpDgZBbD3x0YSzyBGVPr
XOANKcspoTthxbnj/Fd/TrHXbiZJ/avvJDlekRpc3flREY+s1wRrqTkDl3GDt0aWNe0tSpcwgUfr
0g3dW/rOjtPf/r5OFyNatjg9YrIBpEgdcqWyAzY2i9AKG6Q4ZWY2/x/Ct5FaCnfF2Ab6s9PsEaBA
DZvAYRvIQ7qvYBXCOZhG7fQFbF+fWRSb9xZEW8PLxALqvHsGewKBymXqs9OiXLGfEf0QQ5hwGjeO
ublHoKFn94dv/WtXMicLnYW83gAGz1SKr62AwFHl6/Gbqy3oDH67NrxA2pGCuNC4orsNyWajWpi9
6sFWJDwO5udMQldui/+tn/Or4/xdZrZFSnEubp4uRH0SPlO53QRuGbc5QIGq1VjY4B654ayLTdAw
Vv370Y7Mb8Tp+518t1oATSdyZQ7F5o8ykYodlxSc0q6o+INOnxlWmBKwnv++q6og4h6PPLXUF6ta
Vvt/piYDDeC3boHcJOvmCoPmy1TkGtv/TqEWcxTrYZ+fHCymZ455XbQtdLEivBtw2a0n1KBaeIbH
4rlCpqI0VAjMhfqq4iakAIEtYj3BjJvxgjfxT6B8updwKWOebSctW3zqH3ApWVEyEp+gytJmoOzU
suF67gP5jtgBF8WHixrDahtccVERkmoKBTUCDGCkV7WG2desAiSXaz5P7V4Z27lnaGu+POAA66+i
C9/tg2GAaJ4AfKiBSpzt/m4yxIlGjz4lbkIukfc1LIA+/7NkxwkVahz0TnXtbcVhwwXsZ3wWMS4P
ReSdL7TtFYZ5ZCZe6QJxzCVFwCGyx3kTaGecVZKGy0hslllDTGrSjB5zCZnToteqoG4mQ6OM2TuE
ZP7DZOeN8ppKOKOp3JBNaKsFaP4YifzhdTIrJsKLnqenFVVH22oFsmSxOqMj7XKSmiA1pIU3Xgyu
qEvvidlCNla74o121IkmkY7gkSEHqI2mVPWFM4M3TpkxUDQMouPBPHxg+z/5pv2apOHUmcui9kv1
+B0j1WcmZEitHpouYRAbJHlTiXKM4HXaGX54nZKVRycpriko1gB8mABI+c5qL0cMLILU6yXhVklk
1g5ecACQieU7wnD74S/IBxKwSyx+fjp6BmWhppg8lZ8nvRHE8Nz9d+5LoTcQefbSdg4t6O5EUAOx
cT+8me3tYXRAmUtbbHfKHlURKxeJ8dfudroTuVRkI1+PMple9ObvzNt7kepkOjGgBiQta85SKqH3
C6qVT0WgiOw4vQzlU/TceDM1MOHsMnYewSiM2udfhU3PVC4ssB9b7hWsiZHJE0WZJClfXv1TPCII
8bKZTwF1iiWXJS7nShYnXCIx6PSqjGf7To78k+6Xad/hX3sdVeRI55nGC7MFOxXYFHyde8YDqDfv
7DMcH2Yd6wSpfiiFUQzMwyJ6h0m9LCj87qWljqf1GNd1G4wJgVJzxHm6EJVtTVkZADQe3WOu36GY
F/JbvRESbRYEv5aSmkeMGt0LwQIsbfsdPY7LAzj9zymmgUx1+pDOL/StsANLphuRl1j9/u7ntm9I
Oj+dA6cCOWs3xkZrYdiz9rt8817WzkNwv+VvtWuSpYWZBTkdrSQnd1haTpGMGyus/X9ABNYPVypL
oxokh1K0RJa5JL4nIWHKsOCx37Ll/6p4pAGvmLxz9FEj4+KRD0jz0DcSHwu9HXg125nfkbRLWFTd
yMlxC1LHfz33vnv9N4lDXKP+v2p8C3UE7wRLtwXk0mdHW802WyJ+vrJnUQM24ZIU98+kM4vHqsJN
F+0Wl9Y7kBY42KiieyLCJ8YjlCiKYjOCVC4l6MQHnV0RhXzPyHElsleLSa1J2H9UGAWRqRV4gzT6
Faw4jQ8aFNNZ/EFmvyoB0qfujBlvcVTY/T2rB3nXGuVqOaujPSaj7N5jQ4Bab7onRa3VKB8Vx+dt
IfENGkzdAg4hxxIRtPrrX8BOV7LZ8BIUIX6Mvd4f+nhp2NqF4PRJQb4Id8Tl9r8pjmVp6Yj4XlFD
s8usVmEQ286C1kSTJnlfRUbpyuuhnmwjZ15RcYVMDO4FlubvqjmdlTe2+yHNUjT/57vqFe/XyM5P
EWvBBTCM4trfHy9heI6Vg7D35LXtZ++L3HVMDyYXsDadqxCdyGruxn9I8baPpxRfVE9b4/EQuPAZ
h/mzQJa/8H/WbrvKV2aHOpUz1YPN1mS5NIhRME51gTdK3FBKtnZOvFB0N4D93eQ0SOhe9X8NFCqB
M3wczsa5XIuH4AwMiccvDFrcnLqBuzC9N4CKgiRwgX4MNRLJkp/B9RjulTbyI/nGjkWsF7VExDED
DRH1zSXQtlrKEZHveQ7M6AwaVvE9bxmWszcQXgpU2vI8isTNCA/on8gDTBYl5TBbOIVcRBxLakJ0
bEZSSc0mVNuJfEVr7rQfdzNFiK/Puwg1V6AgojSakCe/OTXpiWaA0tT5z3fj8B/2rgY/XotBGeAQ
q7/cc8DXRn1YEyfN/dRXYUwhrL0FbiTARe/GfJ002sP7m98hMK7y0M48ow6Km8E7s9Lv2aCZO36o
KtyhW0IUH7UtzOrIxS3e0mVS4/ssKmRvpym+QMsJDqTA36CgVREVwse7sCdk0uJ5Deaa3gTWoMrt
rrn8N57pBPpwWeenYbJwK3rAMEsm3yEM2XlHi9vihhqx1HK2wOpZR0kRooWLnwx7g5Vjfr05VgWW
5g/GlcslpiQpJWs7x0rvv/Sas1h2tRfp7gv1xq8oem9xSfQqjHkhuAVYtBv3buY0bTuXcGC05yKR
NSPAPz0xmQC0o1awJl4vezUTUalnI6t0wVXN4arcQFwD97VSGrUUZe9ZhernQLPJtWVw4vCroOcV
9I5hfV43HaH3wCTQWS9OSRUJaD8I57UbPmFC4iO9rainepFf4M3oX0yXVrDc/4nx8tvvp0WY5MIs
0Uq3sVZLoI8UzPM+GoaTFlae/UuBbQPD00B368RxnDo3D9CXwd0c4UtqNCoao686a1kc0vPZbKKv
8YMKKX+jFTedy3rRMXMvNMKJPE9bPyC/dEYpyMYC+oiNjq0DKn4DxB/Jp1L9SjFHRxo1yOpyZhaD
6f7USjSHLOH8ywArBk2NYmcJnGE/eGnrfc7uv17nuVEeplVcK8Jh1691X9VqfmfzxQ/F9mGORafU
JLeCdQfVSQ7fdC46Td+353b64yHOQ5rqGFpp85/lAeVMf1LAI6WFQo9BcoSvK4mHUcdr1/ATcZ7F
GkRrtC8EbSTWlfxIiVilz4M8LuXfTyi3opJT9DhPl+Ji8iBzJPZhZ6gXfX9WhI1lezlQCDGAFmu7
5+N43ofL28lM38Hl1689Xn2n3e0tcnfhUF0vPYeF9DU6skudztkSLT6l2zJyHHyI3wTKZm5ljw9i
2N82gp+TQB8uxNqFqVAKD5sIiXW9f2gF5nLeVmw9IZSBRQDBuGnF42VLqgKbRtBgLXjqef3oRFtu
jWG6knRQXyjrT6LjzaFaBw9QNzh36tCBFxbH148SPUgGcg1B+5MZ1BWvN46ML2EyRgITJ9WBKeph
8ZzxXJynzmX9mgTnKEygnsppmZMH0Y76Hx6gf+gY3ryJ+4menlOFR+EmHmawv88Bp0ymspH72o7F
m1vqYSDhMDoN2ysB5H9SUB7jLp9YPsFQgeikvGrF8F1ULWTem8OhB8CfqGQxscyRB4KfpLygjSx+
SKIlHFxwynB2iBTCD3Tl2gKtaVGOuHmrly/aW8VDSajBvGPBgFzQwbPbAGsYBMnUazzgI1a8DNms
7LCkL8W6yVgNvfT+Nm/rYBBGbpy8IbaxafexPD/BA9mDdx8218iOnUa4+ExWM3EGfT6AbSPzQATL
XGZH1YITb8pE8nCuXTboBopvpdmteMQ3ssIaYlkjP7gTq0E8kVCe1iCIrQ5t/75uSnjE3jYtOK0f
G5IWKS5FqT267jzqeVdpGTVVf0QTkhjGDSwnADmAOBUE2lSRR5Ak8DUaIQFQ8Tt2s7wET/bzFWyB
EwAWVgdwTAbks0bJV8LCdbI1ndYyey7R/JEWDsljAI6li8OGXxHunAemd1aSQnkdCY5SXogLFT76
QaWlmd0L2eaVRAaDmpZoEls7hz2z8Rvxsv5baxC7pGa+fQbwDWL6Y4mMS8dlZaoqVquul4VVLMlv
dnTEH7aOIj5wpwJQLPSt/Xa+afFlg+LPetQEFAKd71ol/YKiZzqAU9rDNZQZcr8HyzxQckTkHpQr
jlu6y6driGaP+Q+qJABwSpc2a2sBz+DQlnqpwCUqcZhr/nz53kVOo1IvfGNQ4NR4MoPXbERCxdjA
WBVqp/skS+C0jLkJom6Kb6IX91haD04WWM2Tmef4CigWXbzDSGSneQj97FVbbG4+amrVLYSnSayz
Y6pt+tvKvomuGbtfhF5WZwmuR4iNEvG0+uO5lidMiJBY2ZfeqNKJg0RMT4+ReJfgAlBp88HVdJeC
ofGl7dKkZ6aUFv3UbfR1I/gwz+D8KC1dT8+hSUzoPJ6ITXfPwPlzwboP9+DXeAXfa/S6ci6xLZ2X
UWbESmxXPDAV82/B8rw3Omk/GQkerJPSvitnllcyChkCCXwYneSXCxZVJXwf3Uq+Dl3WM5TA0R/a
La9u35e5i1Pi0s5/n832GAzlbx/vcJl8a3SF6g7cl0oO3SyiR9eDj28ARetlBCAbarP0UlJXMFlB
64xsYb5BypBx5xfgxjNrnaYXJZ/cRyN8Hmz5yfFSHcm1C797lnsg4UK5Tu51ry42XPPt1O0y+DIg
MNAATIYLU1vVlXfja9x0j8Men8MsmE4XESn6qJZwvESG1ZQ2uKeAtXnITPE7mLnzOhqhLF1lNwC2
ehvHoAXUbp0LE0GxUFeuHbV0o5GTEpJ7hV8JFnjGoMuez0tFZX/KE1FwQUwLJlkjVDBluyG0SFeS
sQMj2Pb1EBnsBs04YelhU9cttAl9m0EehRI3/TNq1qBctiOvxo5dQp34UwfczkTIpF1p/1/ZJhBY
CVNdVVN+2p1y5RcgCNeVT4yLOF1skiIc/613cgx2ERoICaSLprtRRDKXx2H9z/W0Ze9RSqJRQcNZ
w4z4f9DBNfmbuhjBUCUQCszd0DaVMUgqdF8+Vi1cLc0CLOFCJwGdnN7MzzM+qCwtQPzGrOdloqzG
DghAB3+6QzGbZePC46y+8n3K76XchDLCrK0ZxkfLqsTL96XgM7kqzBaaDE4QIGKPxhVtsmeovYlK
wqIiwY8B1HaIsyucKTJCEqtNBatYRCvBN6PwZSHobVp15Gp9arjgeNicdwe+i4qe7VU7lzyrDC66
NJEQ8mW2IjXKP1QFMm2VnfEv2nsOyLPX4Y5ed2D/rv5h1/u8opgUcmdqse1bawQIGn68r8zt1heM
pwNgXc/mAJl5qY+b93APWUgUEiDraLL/cyw2D7aC7kb/07b/Y0n9NWE/fpyYBCxSYj7jVUt6MK0S
tB90X2DqeOGGI90WZ/2c4cxRcWO3j4iofrSY3DXPe8U1ODen0EjTSWdk9EQaik4Jfrd3YbDSIGzt
egW18gsGUCEeeM+GlcMI3tATG4Lyz/xqfAmoErpW5t42q1wcyJcGZeK8DC5hStJ9eKqV7kMlddJX
vVsJHapXLtf4fXBH/EonNZpjslq4NXTunv7aS8Moe8qwOONJlz7Fu48CnmgBS6+zVAKnsexuuLxB
IhoRoYH4HBlwUF1EhpyNc0KUADMoi5pUSzeMsqjjP34ZjNFoBli+7rtQ5wJS9bRnRvZfrYP+bDFJ
4dHUwhaJUbPKon8Xz9CWrY3VeUX/dN4d30RP+LfZGozJe6QQHN797XtVxXFoQox2pW6nnKW3lMRk
VCx9lviUWMvhZQLrgCaXZDjvi6yIPeIKPGJlFwdFF5JZ1pZDwsVfgjlT77xjl2j4Lf5ZRAJKtNFK
Itp2zZzWFFOLTwrhqN9rVODP8Xn84MycaPjIuSx6Y1qx4CAc5NGAwgQCxn6pLMfw6ZC1hpIrqWdi
Zbi8icJlPbvMUzbjoW0hFqLnG2Jo6oajq5pcyOllQma+Dwdm3raRq2v5szMN1752wKPWY+V7o5gP
s0onoJGzXLfEiFJDvlOWs/YINfANG5DmPr00oD4u+r3flkylhxZYv8pnRdpiPCCvFqqt5zhp3uWK
kkGW7Yv2L6QB3/SOStIVV557B5KdnziSxTdlti8aHk+XsyShZ9O1Me3SQoG0H1ATmX9dQGgtKPv9
7RzCD3H8rJuRNk6MHRuv0penvnbZyswuqhOOCa8p39zrXqHNmjoWj6fCjp/jzWBYv5vfXdEaRaAW
Htw0gEjx65QuSlLQE3FVXekj7DWEQVOugXu3BTOvI+HuygcwETHhd50Br3WbdQcVZc4Q7A5LWXDt
pz9WBExhk04luxQZ+xLV63SdqMDRV6i2j5Inr/8BEeftnbHCNC+PW6NPLeGp1zeTbJMRKSW4yUXZ
N60yrJyzTN6bmfhfV/D7CBF0JlDXikA4ewhAcV2XgfhD887kfcAGTW4rp1C1gSqJikoP8MJV/v79
ZY1ThBCmhh+v86i79nsbJ6zOhm0WDkquNnnCEFtnbgenXR9WJbJgP9VlKZvgkWmcTprxs76hltl3
G9adGjnHwtcvGWTngJsFFZGxnjFm6uNWK+nP1iQCSIKicfTODwKPWs9fub/BOBGqV/K1fY59xr19
YEZBT6FmwZNm3/tj/hdzhTqrt59jHUWXfO2Nb3c57qAf0srsk0G1XAEVRv8iufue65stdH9l9Xr1
NquU/Zo794fI66aDrjALa6zfm7p4Nrj/mzOuSSgO/ivylffDcj8l/8l5KSTcLnFjEa0XWy2ziY9U
Kq6Jkw4Fn/G8cLpGHccx8UaCS7o0tSaD+ojhEksNMxTBJu2I5SpGiP1Ngzf6VP0ovC86kqTvSTZz
FFY1uaY5YQYkduoLg4Z8jR43IGuOvSnGkHoyWzZUm4KHn8ogCUqh1lG1fx+aW+iQlwwpf9dyLDvt
sTa3s2XMDtwVpDO30g4VaREwbBzN8mjqhJjzc2IMf6vT1RZpT0bu3HqB+waUyVzYoBT5vIxdSJxq
LKiy7EH5wEk0YFSx0/+geLeBjzrn23CrJF6KIyo2mkD/iHuYBNvkvLPU6XRDHSM14v0mVt+M/4Vk
/BWGkE3r830QXJmysMNwDV3CpxkbxHzK1PsbnIMOMwbgg4qi0nB+5ZL65KD7Smm+TZxh2TybeOsc
SssCVRFHQLXvNJ6vGyITr7hI7Bzo4FX2sCC2/ofEKsP/FPFPqIngl5+1EgvjHAxPyBImWShEmonh
lZMUOWRmjztpu2z+u5JkrSuSAuL0jlD+Tun99CRQ3Wl76LxlvdfEjkF6xgDnQir9pEGXzceDHgCU
IxJWoVV/fd8KnyQGGBAIX1viiAKNhrBdq39ciI3N+rm0Q7GxC3WIDH7FbTRzz92se1w1ME14mNQ2
SQKs0/zXNWrAsY03km2Ku0dX4HUBeAOxgkgYWSpEfWs24mCXAbVmwhRVb2sG7Ua1Z59CNcd4ixWP
2cJQCJ5yEICWmmubFcqyib15i6fEk/6l8ssFctDPWlT9j+ZRRFpyRSi9ofRFBtRXUqSXS+nckK42
BLL5RTt4Ue2OfTQSBGPP1TXYZ2k4fmOZGJXC8FHUP1cghRji5XH0m49IR3i3H1Nj4wDxO8v5nyac
sePB8GrlzvlLoBGKKloOFG2O5Br1TIwkpDzPdQvtYl3SJrCUxrhGLsf8tSeLPC6rM+8dn/Ok6uFu
VelmbVUQH8zHzq25C93zyce4uSsjIf223oqYEjvTkqfyqSgz5XWX6qSTZlXkGCEbSfLnoT/JyvNC
Oy26r7MIujqIpLMM2fka40o835Pdzm10odYYRIY3bge3+oGy2Xcc3ajlY3FCl4JbQQhTAnfHFXRO
ZrY/6ZRBnZ1bU2rchnXFdupF+/7nIOX0OlTvZcbnjClq5X/ukZ85KPTPpnh5HUwmlwqtJ5BTAONA
7TuIIojht/9moJAx5dbItqbqv5wuRUQg88tVWC9/W+PyrA0HWGxsMYN8461/PP0UJLTLafSWI8W5
OAifPnsbiwrfhVqGG76UaPA/L77OjQsOITAOPTp2pzlna6FFET7Woi/VoQkXMMkVLhChTKG1lEhg
hMyWOiaNheJnOsG+WSSEEp/pM47kQCrBv1ylSwilpgeUWm5IrLw2gl4FQrQyAyXwE0uglY8dRZjV
QsXwv8u+B7odREGi1R8KePImWdFvSL7VWvC+dZl0qm/zHiqAUdDXR663Ck0SRIvREQzCgHBTPBPV
4YD7IZBIsaeOa9PEw7j0aBNPWM6SeUXs/fSLe3j53WpTbMhUTUB1tMRjObJrH/73TvSTWVKGGjCn
kAegM+JZG1YOm1QHRT/tI0vYjesoO7e8SLUT6xKDHROoCXFvxF6zGjhLqh3iHvT7V3rRl81BeKt4
gXetNCJEWFZNVi84B8PaqMTONV0VlltvvlMyWBwj7Ms4XD41EXesidaAsN74RetdI/w4L82dZkNi
f2bbIj9R8ugVs2FyFMEvmZbLjGTfRUafSyDu+c/AIvd6lm2shP1dAaBvLyCnxjkgYRXUdyS8LsmH
8KoGOf9qrBBaDS79gH5KEbOzD6E3u2e5Gzzg7m9GsOPb+KMR1fGeAKwieQcN5daM7MPFpzY+oAKr
VYfEZe2rTcCn8TJymjVG3sFR4EO9UBtDy/+W1YeyEktAw1bWTlmu43VuJaQN4jL35ZBYeBOis2Q9
iIjVBQrFsV3SVgHhKPJ8uABPschr/4tDpmvqjiNzXHaKISt6E5HZ/XVQynEio1tEUe46iEhW0WDp
sWYKVU8d4XpyTDoWjdkJqQnhCjKU1/SB13at9JRjjaY0kFqaaJpg7GTSxLX40fa/2Rv6cQ3ZDl8o
XtC0avTv7JrWu17dYlk4PxvzGdFfGGoJpDRgATBOtnG4xVoI2DbIDz64EE9PgXX2yZFTI0AKUBDc
qUl4pWQcVERNbzg/+Px4+4lYESaXZluq9S8kXWQOrXASQgMwAvX/pRJNXYsQoXeMA7m7mCaSLots
rXq2Fmux1kmniC2TmLlACK2tWhi5I5HQs75ndCSII3IJSIeM2TluaK2WG8RxMTyJwwVhgCRJLk7e
MSjZuogZTqGSjrPykKhpY4q/NLNqG73JqsX9jImPVWSAm3h08fbMxFt9EwK6K7S/Vce97hCrz0zH
7F71iq+LDyA51UArGzhAmUhI1J9/hzAXQ/UQmWHGUt+3aXlfNTMHseJKs0yWlrJ6bRMpwsR+qnk/
2Cbr3lCvUSJvrGLu3lLvQIGcyuG17u43iGMRRKoZUOG2N6y4sKrOw6dSgHxnK3p2VAD5v28O9zLk
7lMoTZH7WG3vdQMajEncLomkfVK0ZUOfyOUmgGpMmvHCd1aSUcwYkcpABGP6IS6M+Np2zTaRxsuH
CVCrkyE9linWqnuKcuA+xIK3a8GHHnc1d/4ScuLchx9SSzN4ViZlZ8IUYd/7mH0xWe2Sz2msTpqv
hawWT+wYqifqfkHMxncA8sggU+ZLjk+/DjQQzcni77+jU1zeKTdYhMJyrw1ec2OyBrt1YroPDdRy
GJZXS7bnC+IO/xhHRG9a1ipAT5EaZUXMSk8EuqV0d02Qs0PhJDCe8G75FTyd9kodKakM3lFc1xHx
9jcGsExMkr9kI3Ho2zLlZDqyKshOBFzKkO5jcVhMJGek2+wLRvHw/gc0lK3RuHJWQxOO06Nd1mFY
dM3E6TwiF6S7GSUdaaedKykc6WBJFWI5TRlRvBjAp03P5af4PI87/WQTgxjdppxwYKkqMCZENfDe
3vyy6tuOZkzDK1Mae0OiKOIwDar0ilPgufjGwhPMTeR6n8On+CzpuJhILGvSjieG3Sl0ZoiEj+TE
RNRKBynugfe5km/KK88wcVmao+XtkznVBajID8C+cYsCdJpMqnAuISCDJBXfbIoI94CSEfQdacMq
IIWpCxszftQ3lU6+LUd8Ng2Bm11p0YiVeKyHVhTOS9oVUyxdCtRp5wc5BwQmbWidOHCgjWldb0Pg
Ro5xX9NUBsoPn/uw4Abj63FeRuc3nH9qrhlOEDFqh+4pwW2MfjQeblqavjOZ6Bv1X0AHQLZS5OUC
Q3J0TlzpejQhLhwsCpGGLQvbNMK+GEBiUx0L4qTmu7pepU69+ZYOd582btbeBArB6MaNH57Zy2+9
VKvZWq02v9dYoxSda0HwySxf34OEFRDoF3PYJXn3T+4SC7yVBFy9KyGfOJZN5eCDoALq+a48VsLL
djKoHo1MDK7WObTnvNpxMEPIS2qYRDjrDsCFc5NqP5PmxoIhv4l0K8eFGogiJPlE9nOM1a2G6VD7
0ZvbCknML67+MMyWjXGkWlqwkew+9A7PoZrMqB0qu3w/OAXt+gv919UJ+IgW4NvWjZn3vDsxnVT5
8dVJo4pXqmzV3CjV7O1uAhJ79WbRsNcW3xHyIfJmTE7V9ikaz9svkONPcfTfeWc/BsPRIe0SEkDt
5kWzrc3eEye8k8VyXonZSK5USlmRL4hC94oPHW8NVzoeSWHNiFsGa7LbRX6eAXLa8EbY0kMCzabP
Hm5DLRM2xjfZSCB+dUyIjXq9Ex8rfyrEV1A5eJp9bgM273/af8vkBDBQtf7F4j8QCMbeYOOwSKJP
BJGvDewsBhcfhtuhTkUfLYDK8RYsDGR9AFejrCRkZv06PexQp2GkgU4IZMV2hZiZQ2oDU8ZVevAn
8kuxc4ygTn1I9D1J04jcy0x9XSqdvk4Emq4TwVbPzYvhNRN/lLCwe4/5RiIC281kBzMuhrxea778
TwPlYocvxjVZvfFiHhIzvB4AgV/RYo0fRQR9toulAXHT4defjBzIyAzi1sPHyjKDYWGF9zBNOPlt
YuAvA/F3QIPXbFdnafW6tyDfiE1B3YR1DtkNBZ0vg94UQfFe/xakcYGUCXXZyIM4ZBlQ1EuY9bCr
pIj5aZEkhjqIeMJ9zGBQNfdkhAU0DZLb4nYR43EcBXhoOw2lPM9XQRhRlF07rafy8C5MZLj8Wcff
7v8GDLgwON1wNclyXpv5/0TldN/F1qjNPj4SrwrrvoP8VF66jZsXzAE2FGJMicyEaro+Px9N3QDF
RdpQegr8rkpA6vr6GyuoFYtNqmznWgHX6N1cvHaac9oxtv6WkTHcYc6xwb2AWbwViELW0l2JhsG7
savRA0JeFKJNstRcHrdfnRNpYwoKc4vUV6nAEcORmN740JbgL43LTnYg62+Wt+ed/FwVxog37IG0
hBZ/1+7Zq6TC3ywgOsAUCoj0l5f+hnl5EL2aqecKoXinn4UpgHxh1Ce55yamUAZ8Mfi2zarvrOVu
uFiUy9/czoyipvniYf0SOZ3PlX76aQU91lJo7NNz9rnJO5fJmFxym+uE6YKdeJgZpzfvK/YLBTn2
631Av22EjfjKkZiQUaNCn+tdPnMKNCwuf/EzkzFwOKlitWGWH/mY0dm+wJLgxvAOPQRl2Xklq1tj
xqKItcvoEGG0X671um9KsWrNfMlxygzPG5MITuM8ez/8n4k5k9wS7BXZK+aKuJd2SvveRLD0yMWt
tTaS4WddpwlsGYdomVGuNe+rwZ/1mtkYX1t1SPTDlGEmei42geLOLc4S79cr5MMWiamMVxR96GPZ
bjve6cnpArmFchuL1E9vspYBcAW3NmK40gPN7rR3IJItRfUxCqdrQ20I0+j4vFNhBlIq3Jbm+05P
+P/I8+2HWZ5duOQ0uKUcCB8bPlRYfOSY0WKW10cC1/kmJco7SETnbaWfr+YASNaoJGTVOnMS7Jxj
egsl++qOYVUuYWFx6jtJyPEkXT/WcPDNK/tBAEnnv07a5YyMqGv0/+gi3O+vJIVNHC6D6p0yml4f
l/7wgZLZB+6CkzhdMOXozWJVekXqlmR5rvq1ttcAlmaoxAQ1i7O3ma2wE8hfn+CseqXtzCvltMfx
b+lLoTpl3FBdIzIVXE+73dKhm1eaxziXU2QiaMv8vdgwEf2MTEI5d+8dFgTIrBm7UK5w8E1Yp0WA
KGWtZs4nnV7QBU3WwiMxDFdEjcJP7Zn2v/GbkUSwhvlnnsrfFP9A+cse1/kUPAm72ePgoHbW+L6W
y5vyId7H4Eqg8+CxnjNeRHz+Vzsh7ekUdz29jXIA3GfWRJsDeWnQYG/g+JLt/UXBaKPzmUiYKNy6
nqFG5qGHejha+BM6Q4xxnxQRCUxUoji2B8+J7nKoCFsxH4EgwR6fzu+HFCKvFHY76IVQ/ZMDKAb4
XNILvRWAmH4rxi9lLjIILuhvl4ColnqPFub3UX4yqX9BmY+Oqr/+yOJ0K2wxnd67YQr5mcrmEF1U
4/OHTPKQBH5Q9hPhGHa4gyxWKhdgHNROLP8FfHXMqsYaren51XGDwwqHwPkb985eOENTNghRhJ6J
Qzxc+JoPxgb85F8TQim9wfBQtHbaUas2bzsl46T4yQ5iA6iYt/qV4e/Ueo4bBCdFWX2ilU29ziik
JK0HvSyUIzyL/CgF133skAGGsMoaQPz87fPbMBYHoXD+/3mkatJ28+03wIAxXT/tv0kBpKINJ5cF
JOLtRMHvZ+aTUoRRADTmjvio3HMTLpYwJZZhoF5FQo+cU8d0Dom8lzdhlrnO5/jr1+cTn1otIn2J
wnfe6uzWpUvWd5jMiOHR5WJPJJDN5b1QBjAFGkX3+RDgOyTPvBrWHe5TndsBUHJCKFBxpkte/XKP
HXzX6CWMJ8HaV1P4ANWQ/4b2Ops++bdW/VomWBjtJ2v+UYVCiQVtguRDGbZquQBY8RJ/xRY5h3WV
cz1Alf4gBPktadEluFhh4cNSxevL6OI1sixVonUk2UBcWxbGDCB/xV6Wm3OsxRI2YYPLjmIfvjxO
ZoujKzWM686V+FGgnFvWPZ376PKj+VGwl1KoUN/NpjTV2c7Do0S+TFCQ/Mekw6ue3ggodaZvfCWx
ozBkXXziDXVI+Hdnu6fSRhu5kzI5dgC6dTPMk0Ev6XCwP8if6CFEPEaxbQbqRyApy5T9HDjPw5eH
ilOsmewBbPvJZsGqwjUGivYZkb+snzUgjMLi10uY0+vP8eMG6/zo/A1ilja9qPMWoTj5DYz4lM2p
6cAbycnbIkQI/7ghnKK4UZbGmbSH3JX1MMKB1dVU9qvBEMpz7soyCXI2GK9i+quFeieGQWBSBfcE
8joaAJ7yq/U+Q5DMkt23jU3sQjYDJpA4yTZcf9XcApzZtos/ENXqrLnFKXiyqEfbkGNM66u5yLrV
PQr09Y+0IpLqqMdce1q3wPsuqQ1g/n2eQkwkxs3hDrl7ZSDcEg3WaFStA1410kYxMUsZa7TnO35P
HnorRjuhOUGcAxdyAWy5Sy5C0tl4wqSad9YvGKzAFvhc3hsLmsNOh/fw22X1SbifHYKZGsDCOHRz
Wmx+CdrJJ1VYcWH5+e4JJvjBsqUkGP+IdwrGdwB4/FR9Z8Zov74dkZi5jSsriAHLGMfC6us9Sm5q
vUZTFVgWAmYjXPWYmZXZ2718kG+XzCyl8txprVbOZWunxCAjUL6O2woO+59ENnraaOzL80SUZqFF
v8u3pMhGeSZ4Q1X3+1QFp14ZeAick18pwwkeoLZEslKgMrkLWszhKM8+b0FZHSHEWhVPHn2EFEqZ
gLCAiA/91lRPIETHuPbPCL4DeAMdZE7quofBZbAfDZge+Lgj42XZ45JnN7e83CxvRbsWloUO1lkn
pzykYfiw8v0pCQhf57YBrl2Mp73y3wmmSq8vRDE+vSKbwqeOuPOMFdBKOIUhXNTgXKlvCLzW//oz
QKwEawp2NiBZsDW3ScDic2B2rMNSGpflfbL/xx9fgwjyFaw7tN6fwblnFDdqlhyP9qa0dBbVjUCq
ajICtnJMRhaZaiO34YRZ6ogMSfHLiMX/6Cltob65aHrzmcAtdwydcGFLG3dWRybwRvxmpIcGt+r+
OdrhkQcPusI6X9xwlW5h+AuP1ctPK18Rd/8H5VhMTlxEp2QmN6VyOIuQ9KND41w7IjCOJWyjwacp
FWWZRe3VpD5SwP/E9+JigGlZOou02l+DO9793KWDLEpOkLlzL5Q8xJR3KgmiKqjl6n4v+iS0itL0
qF0GDQk/sdUvdJH37rXqgcTlQ0ZFaT6hgDlNRJtUyHiPQ/m899QEfE64b0e9+i51SfcTAK0IL/Cb
KXaZubJOSEM7WW/lQZYUqqJHzym0TkFJoJVPr48Oo/Ow7UnA2qPSh0XMSGeTtYTXmAvNiOBA5ezM
dfDatDLUglWOFiipSZQ0iHOBP9Klnto4wxP6VwiAB/HhuuGJGd5HNip86XjwOESw6BLHaV9B9rMr
eZV9LMrrqvzj7cUCEE6mWXItIXY5KqgshhlRnk9KY1swl+Mcf+tJPAk8N1kAfyO0ckw5MNIjlacw
Xv+aGe6s1HanCicx6oAxHjyUjVB5iul5wLobnrSeZ5rSQuFTdI6MUehjiQOHJNix/2MNtebLvO7w
G4DOmFgJXHGO87Ue3dWnZ7Q1A3F3WNURzEOv8ZnYzwKAJy01RDfbQb8BiQyATU9yBdj97lT6yl0p
Xj208e2ly1GCQ6tv+p6gjcNG4MzyXMlVdAjKsWBnRdM/5DdlW+nHrAv6nkOZXc6gapn4SEZTzVVE
5cPEA3w5nDvAm2WUg16FXwt5FUOnljCgfutAT8wm8V/U+UUoN7e9wBZotwRXf4G41kPz2wZHynTk
0mCmP7cm+4Gh3OrUEZkEKNfICBQ0viLGqMEkgd2nPwq51aG+IeROAiSQ6ZoEEltyoL+N8qZ7D1Eb
X/V+Aa8O4YXFzJiSUNDt+d8pvugwITJtDnAu//DCHqLWQc2/wx7ryqjm2UD7KFVbmvUjhMXXLnEW
HASKveZlJxYRkbuyL3tUR8yrFrkEBAvQ01lqYxkhUQ4XOTowUSQSiHhG3WIcqs9cbaTAO75BQXA5
N6jLQlqIk579qqsGXHSX9KHCS4xD27vlRrNJkpl9SgLCPz4vmulZZqvJHs5c9F7BVamCmpTIhKBR
aPN5+Zq99RxwBOz+NAbTmX87GTH9FTozaHmrq61d+aogUUhyw1VXZMew49x0t/A1IG12sq6ld9Sl
flbomGYr9OwTjIvfDI60JcU1qzb+uB9XwQd2LccHti+SbmWe5Y6IVb8RkozAsvr1k7GdufwuZFnu
PQR7UnSAw6OceYEwhlIr5rH10eQMNCMO+zpUfoNKbDy1EWWOrcp/U+uY+rtc2wvvwk8vyCNE7mbT
bbRglmRjRrLDKKC+lIOnSfMemzuyoBxzkAghiybAtxBCm11N2eCe3N/ddfN0spui8CO+6jZFJnQh
E4mjEvXrPeQgeDKeM6O8vJQ7dYCzWqcQOBBZW721c8CgQhQl18TObu1SaLve3TGJBQDbP/IGzgkK
bkpxmxSHmyzsj3b4252X5wmaDnvKuEBE7zhoTX3CEt4egT8JTK63smF6m1ztJkKPMrTj4SCT35+2
wRv5MujR9AcYUDwVdjDVbw4zATXVYc3NIfAysXJYDGHonUb/k8CdQoNXawKlqcINrUZKJlymqD2p
Snk1Uu7Ge06QlAs7TPa/1ZJDpKuL3CZ9ui+d846oA+i46VrVmE2+opI58B8s/R9W5UbrvO6sx5/6
ZF/czaqD0NeedXFzsXYLKdGC1IxQUBuSK10C9QUclzFuPI5NxgEl2mfviYLbuQqz4SbWhOiiLCwP
1lP1qPY4nimalP2hdkRkr3HVNUWCabs6f+btno6EsnijkX3kHrG3dfD7yQ39g7tVgePdJ+2omy0g
NcpORsZSOUUawxKXOtBXEub1a3PJtH+LGLUJIPL8uKs9XLtAv1rcAdRdy7vwLhKTVJ8XQw+SKPY3
JAc/Eho9XXZ+0gvFzLFVWYd923CieFTmgS4eVESPjvXjCaRt38NU85aHr2x0kkpQVL15TZZew99I
affSBAuA9xWjuv+S/+1XfD2b7bgC5EA0Az8zcOjc/1alGIhlcixokP4A1DzQ31zrrx1lcHn/JTw/
zZcB0eT83VqQaF6ZYJ5OfcAfZYJLboU18QebTIb/dh5aINfSWUEqZ6Y95eoH4WsltlPEAh5nRoui
Y+lTW9iwU76FQp+0VI62UUEuKyGbk9zxwW29MR+idWoOv0R1eEXvu7ryIz4DE+K6oxYxCSVj2SLu
gWZ84qHZyPqlAV//2n5wDi2SFiatC7a6A398tP13AKsYOiOexznYrDcqIeVgXQKf6iJF3Z00rm1q
U4LXKxfbZgSIchmqo4p2QyHVAmSPzJgHLIa94iw6BFqqdlUGmdFUQonND8jwy7ptK2oZK+z6+31j
OoOT6aADhBQa4WvgxwvStmtyevCjYCMI4LTBYSkoHon6kBGpOTrUP64E695pBwK5uWyBtqfZW7JW
Gc4QwanJ6VnQJAStzHYshsVRncTVxEv5UCBC8MBmg/dD1ZAabbahrw+7QydMUYS2J+Em5B5ALlb9
dXkgFk7gEzbVfvw9xnvLHYsyKkuxBB1Kf5++crzki+W18x3Olbe2WB9d5M2kbPpBrWllwtHOsG8A
RbSr5VfvPoPoVTEg4RaQFM08XGlwNoClGe6fk2n+pZa9lFLKHuZVhbHLhaUF5qy/lgceyHLDI4m7
vb24+CvIZHk13iUGsvcoVHxwDJrmLDDYSxSJ5ILFnnLcjQp4KLbb7JY9YnU9pnNuSqJXbzrFBAF1
Q6VKxVf9FmUusBftApgcBSy4ivkq4Swq6L8bnyiDMFMTJ7UPNiTImb6WMm5RDBNcaQftU82bSBf1
zt/juFI4NtqDvQPD2zIzc0SODhSbK+mBdfo/FerMaTFP60jQitfJENfwKwb1RDTrFFbbQU/HWcxp
HsxKKHuLd7f3dIiut5Hw67yspptCXl/ySyfqnjAkAz0U7CXYPV9CzzaOhjkKuH8OHS9yKC83S+DX
mrpJgA3L0vHKGESKKtbNXL9jKPkaozJcUtT8TtQ5ZQsJsZ3f37/pNIP2Uv0662fnvKv863pI8hlr
Yqp8lVUVUX6xB7y5FF2uk9oHhfPjNZHOAATryCh4QqAPGKPgHoNcMKj7qjjWtvxODcV5BBPjyrXf
Kkrwi99KTp++4vrmJgAkOIfbbeuQi27ILxiCkuNI5nbJ1OK6iueN5EO6l3kv87ce5rbGA8Hh8GAC
S/mvksjxgnIhzu00QK+1BQdMXzeclIuQSQYuGl6rYyBbNOHL1ov/gOTM2A4+X8wZPJIaKL7I75Pv
fndwcNFsuZ9BqnDYFer0+ynFo7QmKf3TOKuyc9zuadfJZs5CX4ery52L8RJmdjxZuwIlpWzjN4Uz
aNZMYwoWxireYHMbZCB3K6Jh2FpGgw+ZrNNqhU+OOMP5ZyUfFdkidqgDMJrgjyMZ+xj2Ii96gVg+
ZFjiHmmlPMTqWys/eeBVoDjWoC9pycyyVYULt3csaVZBHRMMIyd1buH240F37z2N9/XwCT8jsv5t
6zT9NHD8xbZYSfS93/h+UE7n8hNB8niXHHHlHMXFqb8x/0UxCAKXQt54NPfb68jWNW7EH21x9gR9
8Jv+bo0tH6M5NGIGUV2DMgqryYjIlKwWYxKKSmNMz+oCnmYfIYSuDE3GnNIiLaYzzfkF1X0V8lhO
reKntvEvu/CifiQ1P5/rqrxQGqkuLqMFLQl+vCkqY6ahdFyubielmNr3XMvq2LBC47cMhXFxyHEr
cO6sJLv8Ov3nJ9wrq3ZBv2sVOctxSzV4OrYg1pM/2TP/eUbDb98hya8HWMX8DWxKolSPJ0nyVxSN
GG0eJdn2JOogEmXVr+h3v6JYx3pDzhlP3ohGrol8cZ7jZp4qCQU8WZ5rqESQubZ9XrRiX5lDFFIE
bJAmRjO52jztbS3Ww26zAnXCGhDlHCylfzX9ljwLhjM5dipXKUaFpaTRcN5g9GmBUb8v3T3UWJ7L
CeUbkii72vEvpyKMkClR+6all0P5GlinDYPfIOxFl3YXokamClp53F9fpSt0iJuOEcD9kdE068dR
lth9H+5gU1RhO1CQar2MO2OWiZuQIMilBCKPCHexuxI80B5uaZI+mLVA78NulUPXnk1I1Kqcgl9+
yUVDA2pC2kKitHxzE/ynrCgey35pcyaQTlaz/rkaXjXPY4C0N8C19Ufnyd/Rq2tQ47zFH6+R9FWi
DZYTC0VttTJA5Qcm1sLRT9JFhh1CB63dCxF0G/I4TEO/VQQ++gQ9p0rkh7xjsWN6lMevrR8WtQG9
/9ip/hT1XFDp+BXZVmbQAx8enljlC6D6tG5ckmFdsK0IC2Kh7zZXZwEyDiKzjLbWT6jPsOr1OtEr
QAYT3hs/V+UPWycrokH4JXcGhQoWdfmByfOHyA/GFc1pBBFnAjLtIkgsDtWkwWR0na/mMCyQ1E52
gSr6Dwpz4ihUICPtRp5ReO3awCTyeME8gdz0XEN11XsLlKe+n39af/eKAp7M8VU79YID73t2vn+b
N7/Ypxkx/1xML+54OmrukopYZ8Rim8PIFr+yXdCkxKnSHTfM+HTtK5hq7WMug1w/khwamJsVHmF+
xd5HMxeRTj0csYXV/3el3daqGe4YK9KSSukidLuj4CsdyEc8zAZ8R/vX7/bbuFTInWUcYEL7ALfd
frWYE3WsnS1rodvrQITn7Ph9TmrLGAWdGkTrzbmrAxuEoD+nzYB5nxw+s2Mw37aXs261LhHZJ+io
xWEykfvURVsfrA4J9KSoBMrKNbdhHyLCr0WNNcKwC3NIe1VITDH/eEhzEpiuNi+0xEJpXFcW8Fwu
NvzIYFSsj5zAOcYdvkr9/cAgyKZvaaDzmlhJxfdjCsuocZSje2GsIfjzYdB/+PhofJPC1+NU41mL
8dIIaIsQL5xMsB7HOavtVLBlCconREg9ZWGK3x5HOMSOF4u1JXykS7raiVuxwfvfUH/lEIwnaYqb
RC/gP81kx7BkuKi7nGme9cS17TYznjAnkYKsvBp31hhq7Xk14RwQ8uz6UDfYuu2bMlzDGuxnKirA
tr+ueQdZ0D76w+uqvcEmRWjDhKsJQBHvML1LVJSBkoDmWo9kbTKCMP2mX6X7nIPhBMXpKXQqrQ0F
AsI+15tJFiP5e+sPyt4C2ahFUQ/qSbq8fyC2T1Z7XbENTTbvK4qdWLtC+Pni+VYR20u6jEseUWvD
0ztQTV7llWF207VxGB0A2A6F/xj91b+D1BxrjKi1rx+Y+6PnC8+/io+RPVBS71oM0L/524tV7JRl
txaIITYAX9YuwMHuAMKNS0jRm8K4/UyV98F9BtiyJICTo54mHZy+ksqp2peb/J+KHC56FKuC8drV
fL3b8tjpCl2uJRL+7YwyT8bvSv1U9VrRDK4zDW6nep+U0Sd9oo3brUvVriPcxn1SQbZoE1mfpijY
cRCrcS20hM68MiPydcPqFeCBLEkLDqPsZ4Bjb+h44kY7pmyxNiupTeGffkZg3NUIRKVeEh2/wS1b
lFTKc+2sudKtw/TMxgk+lMnJLnr5yyq8ORrnRGJkihptLzkNYssKlMHCIx59M6JS7oyNf3ke3vuZ
ikbpjt2fbW+aiCGqzXZ8nMA/E+8SJYpiotxjb1iYAzdDnfOssOtbQHo9AJHGhqxCcUawBOmUdJLt
bk0SE25dZPCMqzLEKlqsRu+a+8fMpPUYvmABafUsNdkAJgB04yWNUI/DXQ5XDcRz+M4RfUF4ik0g
BhX2GmiRlyBXCe/C5CK0hDhxrb8DTEoVbI/cAYbNGA7I3PIivXGQedbYoWEM69ousEKTln1HhaCe
B+KomZ8yDQDH0tCIBdaXxtIsRbOa0RbostJXHdPggUFqE4TYl8q9sv2cGx4XPP/LRvIRgCrRYl6H
7XfUjSJOq8HaB1FscWxRp2YKapHUZ7Tg3PQTJUNWJK9No+9O4VQ/pddafkQ0XzNrzUQgcWpXfuVT
GOryTsgfdJv8ZrkaADyvRj7axVREL1dj39J8LWlPpU2zSkbNJ+TpAMFISoDjWAH16xGXtKtUEKvO
eANBnjB+zggKZRNgowPejn8umJ5U12EISfOO0/VY7BhbhIaYE2NipJnCpYSrYVf2Bxm+GClVAjNT
j0aSR1VXI2FHXNFMI5a5vJrl/acftcHdadxJN6az43mpWfUA3+tM4l9y+3Gky4gKC78sOyxZ3dwH
1zEzF992PTRpbznm/ptV14xLJMcP8BRVxwi+XpxKqO7Z+P3BJWbRT0k5wGQJmkAWuStmm6EW709s
+nhe/BSTjoSwr+0SV808+HXmJvhcFXjHNVRDGKXfUwaTYwpc71G84A5WwByV7BUGwTtr1u2Mtw8T
nIMF1ffX8WgBjUvd+c7UrPGp+6t7gVxteV2vPTet+dyYP6kmEfqutPb1P7mJPfRPjMZ/C+j9ofC6
dY4RNoj3DTxKMTcOmTPjEyZxStkVL+KHinte8C2QJqb0BxuUDFzcMODPYyVkoLm+CyAir6ViU4os
FoDfnWEH1bEvLFgObA4GtVAl7WpSsP/k+f2NI07VAkKOT/dGnuoIWESetDG51W7tmnSOiqnR9t75
7jP3Ax7EdNSLsLQwV6fWugLVBbN9bO37a6JuN4hTXD4/6JyEC9lexbu1sO9p7+ER/jbUEqjolRIK
uoF6VGkW7/hE4If83U6eK3XoIVsT9SjG1WVuenrdoG5Ii/YxAd5n9KTWM3gcv3xd4Y0ZZ1+EvtoZ
H+pKutRDoQgkulYvMrno3sEEZoeEi6YMfGj4e5NYu5BntWIn+Fk3Qht3Q8C81KGoU1oNBQN3f6D3
+RzJ9W4sJiY5LdiYa1TwKLSU1n4XMDmAOZsY7e/WHBFYjhnY0Y6ObZxBF89t/oWSokTKa6hXGPc2
IKbgsiN5BJesjZ+1j4VrtsXR8xuhjunqGLXCFjab4msTAjANaPQVX+5ULcrTZsHSh3ui56w9Iy6h
WhLQbGYDH4tZmj0wSeSgwIIMWOGwYid1eIugO1TKZEf3vFX5YXLTtKXb1Hi6HVZS1vprcuKABXx5
SM86wjoCJ1z1qE6fP8umu5jfExBQrBIBDiwkm9eHXbWqQNEenvlZRzsSJSTu5yT5NP3isPjEcuOu
KJ73moBFPTO03TdMF9qvXAuQp2JCC8S2/B790S6WTIWBAJ/w1ezwp2BCIcKLaEfEXtXUq9JqLHBM
HPXb0d3vTnVxPiwenXw4UWorp3sfBTpePND4wc5tKEt1dkEM4pDj8S6sdX/UpLAjS5yaRCYtcEdB
gKJz2YSIZ+w7cFp0+2jlVDhTW7ljiM+j57KO/g5PDhnJn2n0K0Ig9Pm31N9CM2tB4U/il5I2uDVd
2telbC8rvVVN5rBL6amsXRZUkcCrLI2CZ/Qw1kUjXqDlU4YAF8hb+stpsF9LPCOSe2duc7JBj/1Z
U8YdZ5V1n6qZ28HqGYrntzUG1tcKwg1DPz48avuD1AXr26dZAZF5tvFJ8qNq21eum94+9y4tvFFV
qyMZL0TS5GnrMThrz9eyoml2lpxic+z+Ok3GqCo7e76NXSNeM4oD8ujU6G45pz+xeDk9t57UCtdy
IrFte96D3xhEx/K8wR2u6WoTZzr4E34ICWUKImn63Yr05qOjbLuBN17s5f+PCmRe/mbX/Vl24WSH
7iOrDG6tyzkEdnlX+dKT4HdXlMNv6XDdYZ7+hS70BKfOlqcVRx5SfcGIzAMBS92+lBLrcfRYW3Ls
+80gRpMfe7UsydHr2Dtw9IjbMne2RzNG0ikc6Ss+vpguyPmnPGO9QB1kcWYJLdcS861ubfaWvvVk
5xncjCA6D/GgVVyAafBkqJTgjl/eUiBAqoyoWgn95QkTlwBYGMzGw09zvrjLMUmd4QB0pe6aGH6I
QkiiIN3kaT7ED2R6CyWhtPbRYZwOFDtqEM4ROcxo1GP2QujsiYRGEzcrQac/qlyN9ljFVuNz9v+7
H/ZKU0kOdrq4qS8iXL8OZx+ux6SZRz+gZPlcb1xrBqtxl/jOgoAaNPPupHUZtiGj5pjESGnLqFeW
zret80ld+W52u0TC3ypCArCXbJOQaw5pN7cC8mUF7bpZMWo0/yTht2ezsF5HyDaeZWgD5guPsACR
t24MyAxD29E4smnK5GCbHKxM22ifiWRxKE4NRSnXyXEawSIjCV19G3W8TzG/GX4SUcsaNHIKY+xk
dhTFG3X3D6tb7ZS7DuULcRk51YECdgKknt+yYOt7kH5E94NsrbJ9FKvrBw7gQ7A0NahQe81vQNT0
HgBkC30YFoq62aYXNyMKJ0ZdYYcyyNhDagKtNTrnuC6Y5I6IuTOiIGxovcDK11P0DUrOEsQp/dY4
hwWq9tLJkDOZ6gToK4CLFAyug+k0qAeGqRxMHmeRoXHd2g1uNHG1C6D/6uPk8WLgtL4KcnXyTZwS
qd3JYZpY1juBmVCmND14w5EVNoG9/LlqQ8BhzxlGOyUqFfaO03RFcjlzPfLAqOiHniczGdyVaOlS
T5wLxZR3+h4mfcF7rkDYhYfRXSZ8O4VZkqU3vHNBbrZm7BTpzuIm3nWzRUIpwD5CIniJJT81BEJO
RkMM3AUOO6o3aaVQdI0vePcTZXCrR3hv1pO2cIduA/0hUrWeWOX9VRtr3CAHzgvlaS96IAS8w+Xi
jzQBqh2iLDWIk6XB6B7BsjuiLokFrxNiEN2RN7woc+KPQ8hDC/J5LiNZBVsWb4GmYrdw9Ejt34/C
jJtEt9c6iMZakGY0XDk9yhCpnNqB6+6m04LUYh3NpzEDTPbIPy7GHNEUKQXe0Bi9bu7E4rgBfrIq
pp21TdQkMefpNWxwEEvgkrgQ/Cf3211Vqb8Ow/7aGi0m78dFFVIg6h9anpHH1rdnvCswnFTbmIQL
Pj4nRAf53jCAKGXiB+PVxBhsLj3mFNPatqw0tqWA5V5vKTr6drhGqYso0COHctUBn1pnKeHN5CHr
8VqYDKO0xi/iB7QxGKGY4oBnVEuewmBEpWVR9hAuzjvjKTBQ7fNNnZaAz8cG6sWHUE4CM7NlsQ2d
H/JeTAvFN71ItRH+fbDRlX5VJW3y9uHPnyjJaItkmkG3lPx6pez4DbZzY2gPqlkP4FGvSMXnITS6
fJcrmt/CvFMLKUecaPg64jdJj4SlVa5cRO6S09OYYUFS9XGUFhc/qjh3d3t6guproHiDSZPT5Quq
E+NkeCGL3V6iv569kBQWHmghk6k4LL6edtVf9KyZQX0KGiGVChIqjqj98k75p5mU/FaSzBHFNXZx
eF0oTbEGe2q5tq+5iT22rJxjZfPZ4YOXkmwr/8I0g4fRiR08v8PSQAKuddpl8Kx1/TyldS7Foatr
jv8FPXyBrYB7AXi4t5i0FrAKod+AWNZwUczjYzEcYK96uYTy6HODtx09lqxy30GYuEJ1UqrgnbZg
S6tQ7QdJ9ATgAeF9WkokApZilTBWKW8GtFipjGaHfWQANLaOgG47V9oUZCaR5xzjwb2eOcI3QuMc
vuyZr+b7OSx0qJYsdk7OeH/EyEpVpGAesLJUq2N9LuxI+tqUi6RwuEuJ3HzokzdbL5+vk2Zg2OXK
bS04XfrJ+fhEukeAs2+UaQpYvIS9mmW/I1e1Q6OqF2VfU4eMF13G7Uf77a7kH9LYbZSVqSYzSAcw
0OAalmmKeDuuTXScvRGfSUInUbDpytLLxbx6GPi7l/mLlFNc+PXjhLvicHLsGpXP+jvgrtJsaQTe
v1FUgUAUEvJsntjfUPFhmAmf/hRdQwGxAudROiZV2RvB8g8KgozOW1LfIDe29XW157A6sbERITOw
E7mtwLW6aWEX9J8FJMgNQygPYt4zM27VQP2S09Gj/6yAarXFclyW1LAyAt566lPXG72J3DRLThpU
MSFYbezQU5DAOFNOSc+4zPhOpT9LYtB301EP0sH2F5rH1JLaiBrWQUVu2TW1oyM+pzVU6AwAqYYJ
EmagoOpOYisJdLk2loDyGyVdmeaJgOfyaFV6QxKG/aTMcBnQ3/jjia69uPQQwTuB3v5aU+at8j71
9kng3a+g/ZZ3AHwME0REf7sffqrRpl7qd2Hu0yajX9+iq1GYYKYRl7vYdr9Q7Z4am2x4x2aZp7cK
YDw6ZmSxfH6que/vu4g8YP8pTDb5RHlujnoC5qend1+c3EbSm0pK7lqEVstPWsbAC9R+qXFYu9/K
XLFSVVSNg66eAfzlPeVTZTqhut40hfULZHvsd5WfiyvGTlGRneA5xS2tkZyZgM4dxYJhB/Tj2WI8
q8aXVudr/rxJC6JSfy023PAD+jmsqvOjnVFkQb++0y1qMImUf7bJMeklJdjDAnVTqMZR3WtP/NRY
ttVNiPj13gw7R8BjbeBMZyFA8bJTtmL9S2pxG3tY1EErkuYPCbhl3j3LNrw5HB1jqw3R1QAmuKg/
0Uo/T1CTOG2k/rlDf0AvxgJjsd9pypySZ8CKrw8b+CE6YtPIJg++tlor6bRj+TW+CsWKLMIENufh
jEyU8/ny3r7W/PesOD1ZLoXLo3AJDbt9rGJcpANLg1xhh6+fcTbOXp+/FBGDuNZL3h/AfcUAvt0X
GNXzLAdi9+9Pxcijd5AgJ6eh0dA/89F3mdiI4ag/m9P8d7cFhzf/W+evmaaPKMB0XMSAI3BNjsIk
NKSO6yaXA/Ir0o9JanplYZkItgYUMvGxwSEXsNlSZ39lph3d3zUs4ieBJqtcWWvEFkxxFO84ulyi
kkAzgp1tfPd71dEABb2QvdURO4V4pyCPI6Wka/mBVAJxWwpwwYMLP80YXSnU2oM4CUpUA3bwpem8
Holk14HFQlHZ4vjIRm0w6V4a26mt1mbfTVq05E7FaLk1i6L1gcoKXaXKcFiQhNfxBqaOuWf3l24Q
rgIbm6aRrIHkLLKpgc3n1b5bHz31mnBt1wryfRj1It3yMEl4SfjmCxEOyMUozPh/wtqY3Qz+WSEV
dcxPlDle73Hm+v+QzWCUfOKhnEn/MWtO6QkcO2+X+2ODnXPJ0tuibXWvLFz6OULP28AqbBR1mVx3
fFxQPssreyQ5owdD5lXy0EYciar66yI/yulJSzTGpkfnYi9huMQhZ8i1QNBaM4SEf6DbKEyTyuUt
JcA7oL4KL39lXp3yaGgd54/tIfT/POFm4g5od60dEO/QYButfG9e5EW2fdT6MBxGw5mUZwtpDSMP
2JVwTtW3i5Q1kE0g9kWii166j7RrPigpnsXWYSss3Ek0Rn29El0z2mjh/28guSr2a9gws8XwYbsl
LGFcMU8R1prcRlZRW1D1q8WqTuWP9q0lHKRrnY5p317bIPcd9i+1BkeCfJTYfVeYm6p3TXMCE0Ph
4HnEKKfuV/AqU6hU2umvx8igg+5xOy6dJgHdarkX5w7dSoEs+uY0aif3BPxWVDrmX+J6NsGDPafH
jJFMgSfi0VtAoxrgxPPuA6RJ46L3h3NyZmG7ZeT2VLlndTD7E11vf6hN02PMk8wSRCW0OpkmlJ5d
ZcGeM1vHXytUTMsxX7BF4CTuYu2n9bzZNbYGzjzfFk3dNypOW3p1FUmbX4OybCrB+Nvx3esRW3qJ
5/DekrujpZUYasnF+97EbhzAtIEwrEXWOMlLcofzh3VUkeh5fdZZWnVmX8f/isaagWH0SllDvsEr
kNNXU3huumtZnx61ymkAAf8IyUwe9B4OeXitVhVRYFWp/NLE3NutnxsO8ak7QEKTZSWaOnqL6OHP
5Fq8XZbKXO9u0C3WQAfASXIVO4kOcy8cyROiDmBC+awD6FK2JJBLRp4amkii5nn3nQvedrVMZEkm
kCTFXxTDDgmXou46nJwC29Xo//AxU3IREktVSjmnTQsCp6KrRfO3US69whjQRyS+jdwoYg9PWnB9
hjIcc8Bu2e1xvSCVonXsbWtWdHvemOFn0r9g0ZeGiMc89sZJ7I9ogXNuCyrhVHbFR2XszqjEtyBt
ithmMwrt8k3qyfqml3zmQSCuTTgeKBe19HNzDQE5BjLtr0jhoQbplQvYZDoQS7EKlErbjGVxB3Rw
7+EmlLWaXIsJBFM6K9mRUMDUdRjY1ZSJwWuYXlkg1GzPvjbBTStCBMepTuZhWFQxamXA/w51Qoi+
FYN3fKtsjs92LpDS1hCXEtf+HpfEJd7QJ4Z3GM6vVJGXas47SqJhD9tinfbMIp1s5j4m0+nhAwkB
ga0j0cC+PZg/X4721c6L5OaFEHzrdr31bwb8EHd/mpKjAT9dBOtLBhNkfZ6Tt7vP7GTLk68Y77Tf
9POjrYgSobQfaJMtLQp4V2txNknocGVuhN47mBCLUZij+4NnhEk9DsJmvhiCh5V3Kqt9XbFhJ9+D
hdz3gTqtexrI7E1v5sgVUpYrI7yqxsIpy/FtUDAtPNVMN5Z8RGrYR2sVHibo59z9AzCIUgXNBCRf
8vNhati7p1Tq19usSjoG+CNEGWQXvJRJD31ikR8VcWWAd6i6Iy1y217HRs3QtiIOxh3ylSaKNyMh
1aLt05D3TGo84vRbgu701owGuM6lnF2cfDK0u0sLndgFRS4SfqaMWpDqwApnqtCsdAeo6VE2/upj
tr2TdbkJt6rPQqk1E+iumVW1UYOen2emRNlZAcsdxzffSaP5Y35km8mCJCiCrzbd7X1ENHOGX7U8
0xFIpYCllCNAoSBn3GIsLUSoDmO/q64z2EuHDrZL0fiE1RcIyumVFMXn/hDTqI1vMimL1k4An1dX
gZnY9A621HiCB+P2zoyvJ4FXjIJvUKb/MLLlNPeeDTWXSb7Ip3UlurTNujEsAfnSrqk9vH23Hr44
N5uL0Kio2wmR3QLugNySNYj5uyb+COQ8un3+1v+6KzjqG46+ssnAofYvhN19f5ZyoxNLpuPvH3GK
h+oxMxAhlyxntWCosWV1pxrVYJMZ79p0uytiME1UDSRFi24thWBdg9hw2ePu18lGhxGtP2S7jHF3
M1a5bcB4gGD4r488CdOlPCxwP1cg4Ikvdadj4Z44NQjZ8mtttO7TUcoKBZ5/MPc+GfMH/Xs0QQIJ
qWuvOU3/USypEveoIyOQoyChhOWp5BdjXqzBaFYNj10FBo0yGW7cikg7WQk1DS3k8djGqY27zpQ4
sO2C8B159VoVPKJ6AwrbuHWKhdey1qcDDwLBOAI47xJd4uWKOMI+wYSo7Kg9VMH6rBgdAYOCNSBf
3mfcxpsGFjiEb/ruC+5WwaCgCx8hIzOJDapU28Z0KF9WfCOzYknyHCE41xa+rhBkdYCN4nH75yLo
SXe6eis8oIwiGWJ1MiZyR5sI8I1TjnVKv1xxVkP+pAA8mvp8xqSz41j+V+ZzEZXF9tdlxrowQ+ui
4LrWk2GxwqMUuXZ8krXxs5tSZ7WsygFitv3XnC2R7ObWigS8qeF8FtzYqYBYS/tXQSURC2/N0vRB
q0RXJAIvEhkDtsIWljXi+zjSIQkJj4Y5UfvGE0ocBq1SQq1NDX1HPTUGHn7dDw9nD/RlU+4HVGfh
zWU3KtTonC0R5HxhxuhC6MDL8HckVk0tYS62BidowKCAGp1Xkkx/YVQK65np4BBSQfFkaMlsZ8nw
Q2oe3vTEItIhnUxukzcm6vQrlmDT14YWz7EXUzhVaCCvpdMkI0/oMWTstyyGW+ZWUsVAnCR2+ADL
fi3owo68lOMicQeeNFcxFFAhegAI0CT3qBV/24jWZadq686BIRX9bJsLknOrV969KVtbwaT35+as
Ti4+MTLgeW3HTCXb8nZby4+bXFv4HOa5lo6nzdYhubqz6NvdtaydpfwgPRSzydAm5vceZ/aPIiEy
XuntssWCpzE3+fgNYeGB2gRI9UN0YH1c7LVB8d/WFqboboAbDfnkEV3+8sjI2ns5NtZAzgUt4NeX
EKte2kX2mlllX45US50fWjQ9RY1+nHjiIRY9bNgZR1fJ8zI9XzKri9sgID3Aba7i5WD9Cy0jTHKl
82Q5rgtgG50XNdWX7T3gAZF4XNaWuYxp1RAYPx1Zp7pwcgcSJpnunplMJW+2FThCOilmQDv6Cnkt
XONt/qDOe2tNusM0Q2XrM6dtRpmfUTGnYaOClmZ1SWzGctg32a4pnrrRh4Sy9VkmaRBc7+YxiL0r
Gj9/kHteZZ0U43y8CG+ltpTGQpAhoqQNeAvN3Q4ORkUXhGKpdQM06HT8Zg1cswdM+hlPJUJD1/SB
suyBU1tChlyGjmSTGlD8pAaaN/ilkql8KhC6950quxyMVPrhszzL9wXxuKsP0rB0n3cMgOK7ia2c
n6JTebbg+RD7NVNgx1woApCU+UIbvdDprd2U891nVKkgQD0QAQIteh0d8pMWj2nsLb94BsTz3CxX
x2FNiwhVeTqDcrdP/Ad8UOgj888CRMK+3fkcWs0L57mwVBTMvnQAYcyx8H+TLHOmAzfvMNAgCLpx
tWgwNSIytjO7qUsuN/0SlFXcXqJ9Bv1IE4bEqKu1g02BJJR0sBDhRQnKxQ3xxxjQXMaPKaTPsvJ4
rpLA0FyKJcbAlsOEXsYDzZnGUZGfGMVDiOwE2oOxztNit2wrhifpq7Lk22UdUWouMSPcwTcIZbrj
G8wPgTKLbLXTcpIlyZYllmWUObDN2o5DHTwhocYiLDzGT5n7Lo4VXrGUJ/zs9doaWcCuAJFoBMYB
J5oJZOLWmnlaeBq94kgVjHXTRVSsaBRN1xYq0IqyDPRFvp1C0st/Yh+AT6VK/L9DcDhEcXfO9UDH
gquEQHir6+pXvlpj3rEaPr7JH62zO+yCfvpabJqwNlVHshLSpIqiKMk1ofS5HGT2Xx2nBXcij3Lb
9li2g1xAvVumMdM249ZtRyGn1OXETsaf4pC4i8N23dxz/sj2WoGmWQ6HvWqsGIReueZfmWdJ6ZJt
cVy0KanBoy5QqHJbPIl0dslcmpTV8VjYPnFsYdWEnYI9RnzStcSBg0lPaXLlwCch6HhW2zVM/JyF
c6eqjNfc28wyNWlULIOUQI7BIUSQZdxrPEvyjBgQpyAIu/IcK8ieTMngHLjxsenytY3U4kYKMcr6
J8S091EeBnimBYjXa8VUP3cDVyssNCZUObsowE7hKLM0FX/IsSeZYAaflG+5TTzpnilIFXXLL992
VN4uUsJWLKKLCvjG9tLGVepyUz9UqZz718u/DdsX0RvnbBhzZEYIPKQCzxU9tGYI1Xc3Nu0oMBjV
TlNZIetNemzZcHurpSKjGVBwVXrK826qe/QdEQ5HLwUMPDyIbrEWA7dGWcg66H4ZKUvQIcI6txOE
LY6kRTwLxetK1+EPk+zHgCJqP18vVrsRF/q7sR33WaGMJhGKcwb6m4O6DeVLrAp36uBa+gu7Szub
9Q+OfVAYwZ7TjatMQ/3agoO1qT83/FvJGtwaql+2uAfZprqvIPElkXfgvCFoItWMfok1ggeiH9je
JOAaCLKx36II/nZp9eV97YIrNZkO/vYITKpZPUZ9rawJbVekaegp5Mf2iwXuTfXY3sMM0fuNxm7Z
zsIGwGPAuGY2hfngptah9gi0OypE4PiKIvjGwei2LaqzGWGKxSB00EXF94LBrm/jNrNEf2yYqTLO
ZPiE5EDJkC53vZnvS/hWcvKU9pUztoXAYsM5Lrut/u4rkrRXBfHa3RdlBsnctGSmIkf+/JPkRzMN
U2TByfPCsOC+TkoTg0ul6k4wt3MNbt7YDbEn82ojL9vZr3a+BLSVDihBS+NcO+eXRl9bmM0W+pYC
Iht+M6fVWaiUxMH03zJpYhORyVODcFjC8GEKKb1GB8TdJ6aGRQ+U/X9KZo18U+3Ngu02HEQsMNgc
noxNnioWRoeR/Z0VxYuaKDGah9v1f9CRdOI4HVCZujMRmW1P4aHiRzl1v8ZKFIge2fRYCHKToUis
LeOHpnK4VAEnkP4HghGC+SXJcgDB41IHMbq73fBrxrIcB3X7zidxKpeZPFFsF8EsahHLSIlHe6M2
yqO6M9+dFaROc3hZGwRkkGUf7I7/Z/DYmm7RXalP3Qh8tiyo9jkZNqS09pC39EvcdrG/6aL1LlPD
HdUpzeF4gJL49nYRTUJoZ+ZKVf1HH3rUl+23wg2ZgVAzXqD9U/c7AQr9zDr02IHhhfJAhbA1jYpF
XtoAultueFcMOmtqH/ZHJsd991ic3VFreh/K8tO73Kzok8Z3BUY3wDRN+dHtGQDEFtRAd6spTW5C
DlTFtbFb5YcpU+CUXXhpeE/S462/9HyQH0gqa96QOcXpAJv7Vu64/dLRvEWN+RzZUPvMFYroW1T6
QqjPmm2IjybCwvH1sCXjyMffHR/6aGhXBToM9tUcWBeMnrnWfPYKT9M4NowXH8POvh32Agl0Zu7L
apw0Ufm6mfgscEDhnCiJru7b1h+bwY7Yp0hKBTOMe7synx74ILg3sU+bm+f3oADI2B53R5x+yQEh
5XgKgUi87qQXDaolevrcwfNiDMhXx7L8UuCMg7w4+e1zUDiYlT4LQUY90F87YUJbv8u7lBePwEcv
+jJPRh+okHQATCkVwpvIP2NaOiJyRI5fvDQwnG3oK3/xhZDisaKbsTAieFQ1K10QpjWyoqdHD98q
XkHivC4y7K9Jw2u+tX5LD/Em60QNnrs4dWSZzOL3T7SDoL8e8ksPg1S6V3rrPejw63Qb/fkGKsLa
2rPvnrGtQ7aywJ1h0IhKuklbbccqmzxq/8U9+5WwWPrppnz5x0/OtDuslN73W3uuorPxRpeV/r9k
ZtLD3O7FypsCkzO/r/U7CdP8sTYiEdx/DVloJ6QwkVL0w5OV4OarKwFSUGwpvHe9Z4976qMD1dfe
3lQAmoKcs3CDA+OCw9prKu7eHBNzHoxLrCFzHiRa340Ts3z2KuH/grnaEaJxv0U5DLkYQon5bCbU
chO1C9kqgqgL22I8Huwq/vd0SxLBjanExEbVqNUNMQ7llNBQckzwnzMytiFwKsItQ5gcIBWz9n5Z
29NHDDDvXjo/dzv5z5x8y5ezMkgB2nJ3kKf0+Fb4HlCzol/JIjvSZvR396MugM3f92Vw8SOsa201
DMG+/r9GWN3nnWDI8yuORdjsC0Jj2qo5eBAqcyqAxQ2l129whF98fFPWMOxwk7yy54Z03ifP6ggJ
KtnF7R6O9oISqCmLTk7WACVw1Ujjwt9/suOhuhy6+DXB6/CPsnEqXEr2uvfjb9o8zhVrknx9x490
7LpEfNH64Q8g4S1y+/o9RzcFrTtYVJY0FNzVRj4V8kolgTOvLvTePHJyGacLMil9+MEXE5kzac1M
PnZg4G6Sm2QO9DAUvpTQrrPr54qXoilKLCWfWptE+0MZPiNwdpiLZimnr1CQq94s2wgiuXMPUu31
z0kkd0x6J30rmyCgtRxInDARqPO3yTpuSDT6tE73gfeoAptHZSRQqlGFTNeZnhpnOXLz723ee6dv
lTv7n+0JL/ZOrN6gXcHnrwxroNq9/ZOBS+h0WPO5MwlHXe888dBaPMduOvuhOYwcHoAgszO/Zz0Y
AnK1Qc38O2CjOnZSNxnW3rO7e+5ZtPDkwpcm1lTM4Vae3VSwgJyUX0uZctbgLLpwd4A4TmH78dZ0
FqNXddNxBm0ANTqzCoezleuLXc0EBUj3MiB/TcagCxCp8IG63nDgjivxeuYcbhgK/DIadBrgCelO
fyBFfQxPBlcE0lfAI/N2lHntRnUvgLF8mjaXLosq3DObpcSbFu7sueQHdn59IW7rBFZPBUVe3oYP
WWZOd7HSupRlnGiD9p7zHd9LZFtvCtSGwGQIpv8UoCZcRtWiat4vv2qa6+TjFaIyk3WQ7u9EcMl6
Nx4/B2Cy9dDesePcd79ZJlJiVCYTLeypZ8iieFRPNVIH2mEhXgSf8k+an8xTn7A7fqtsZIYJuge2
rD32lV/78JyRGXhb7MHvYvh9k/zU41bRM2PY13+yw5Fg7VH9wce8sf4B5CmrcqG9kk7yWeXVV6MO
VV6NeR0hWvikK7zmIaItuZAB7ow0LWUiVpwXGAutqEymTBwzzMVk7HlteXmnUWCIkYvxeD/Csn8s
FRIe3NfKIdfdzru6k5KUmIXicRLpr70WQeC2APuAxCJesq8/M/gTwiN0nBh4Jn57DbjgtCpwlE5v
bqUrOXJukQ31eU/26VuGWp+34LpSNWCoteawUjCzuDcsb4u+JVut00uHicfNYHnwoJmf8RcWNK15
+C4Px0SreA0fMd5b593j6Mvp9HejrcYffx3rn6ntjrj2j+w9rr9W7HkFQ7ZaFrphrXCA20xuIc1E
d/Qt1pbIpyWZTYb5mqJt9xox2MBCXA58UJ/xbjwdm8N/cdZqXBw8cWZaGf5JGm5L5RAFN7gh74uk
PmAuRIgplGI7MBF1fkIkGjb6/szalJyMTeWT3mwFQEIJIYQdm6BUiVvsc4lBl2hvjb5FxnhyiSlF
k9ET7zqFZLokHJD3zqpR3o03Bx39G2WppibZXciJuKB4473+x5bDnkNqaz7tLZgnR9aZTjwGToKR
DdkZC/AXss8dURqo2HOI9mM70GQ/1YddmCXhf0QCXBrpgZqPqT13Dlh4+SJesIMKVpGvI1vg1Ih5
liwtVnjifybpigaTmMBrWm8Yo9ZTgVCVDe0yMXJCh+TyU5LgteInljDXCXC3Ky4xNarerzDsB16s
hATLItoHPYWiSWzQaoQTqaqk9+DJQOPhG1j1jmU1irmxYVdnCksN3MhgDzZnzwxnMpr6s4pxEb4K
mtV1MWv/uek47fCB9J46LOgBT81Lv6U8MsRxyoLVLdMESTK7dqGTR8wdpPOXsnR8IrURCyTFL/zf
sUNAJqhEvH1mxACtQLz3lUcIGY2eGBYgh0KaWG90Z3E2TVLFTFJ2g7tKhBWCJUoVcjrlhDTfcMkz
9gAY4dZaD+aD8kDssShQRTTOc7r2rGZvcwJ4N1sII4F+yycQM05XGGKJJMpwTVJYlKT9zjM5rkja
Kwci1noyZt21tn1tmGcI2anEiQ4J2WIiK/tOU/LFbqO4V4IkJPKXXVX6nEUBHbsQ3J66cART44OP
5UXD3GCqULZgsQ+BFCNRI08UcHaYf0hFHpzqIb56oY987+f3KmGQvEqqiFj8UVhn1C+7ag2CwZUL
+NbQCWsu0MBCzlIES8AhrUbBli788d/NQ+UDghn8dC3QpwGCBKm/Movf9mx7TwV820JsGw6AD7OB
Qu/W61vR5RNyLxyrsX/jAjvgVA7gKikyM8mCdWsdoWjMs7ijSh850GBV5yukvVSUTncrDKOJ+lkj
nuPYb/IX7Y1w0e52q0gAp+Acyw6P6+0/fHw/YUGka+RWSBtlef8BycxuMyZsBAhIUTjfF47BiTOJ
zsMi5KOXr8fb6TugLGU+QtfA5Lz7dTV5iG9Fi2F3ELVQ7EUySmeXNqu/jqiXIpiPPX8jFlaZkj4E
sm+eVWf8oZDHXARuahGUjaEbyexeX7Fozacbg5Zpws24ziDMiTT7R825pjstyKx40D1l+HwHbL50
x/9J7grOmu7vWANNzTAetpXJofuBpU6lu5CDSR1X0K2596QVu334QyAjr92xYJodzWXTq5Y58KVI
gX+BkkQKRXwGcbHNUpb27qe/82rc/tWRyAcuqO3waZD9rpF50cSE/hr2oSXP6epa94HZVg/tVIw6
34GtDCd9+Pi/nWmDofxuyJasr6qGqnDZKegbdCoQvYNbp4k6JKPdEZE44V611RO6R10/FzgEPZRr
/rfd766LSeuQS5YuE06WlOBIdfgPuAbVa/fpzrrAdjgs1jfbouQBWZ+tOFmIwmZ10UmH9RRXmPKE
MCOSYG2+nq5yqRaCFMmORzrc6Zn2b/xJJ5oyPBtzxLU4jNTiSvLgrNuTMWYtQB80TU8CD80Qhf6D
+bxgZtLlU8ye4V77sEildSI4EQEmX2ypybjw0KmDaYMaPAOuEph0W4aegaYwSZgxX8nsEPqiaA4e
y6DDXApRNBT3SsxHM+T42Rz/LaUsqy7TDMNVqy6btBaP20FMW5gTzJaAEuNNdiAAQUWe0+0Gq5aF
YQfjZN+2tf5oxn0ghTRAdO6SDZq5IK2E15shGpJIpDqsWnMLKkzbd+u8lRTfmxS/kxQ1CZ8RRObU
/NHP3bHlrVtWg+s+A7ZjyTChWfjRgHUYgoML5EWCHOaqubi8eWAV97HOZPhV0BKBjZgQkuvvt4aY
GuHpNpaHdXaa6O8hANOzxcJRtMLfEYX8ZWBFj91Qk1LUOVWoPIP/3qhR8hSY5E47pvmqJsQC0dN5
BTQ6uB7SX5BqngSfiHA2jIAc9wY/J3nWms+wp4FS3uz/HiwtQluG4sff91mFb8krvPilDxhith95
LsuZWiG+ZSbylZlf1pOZTd/MLrz7MmN0ZjgNiFV2KfJSm2Ou7kLj5zGFY4vpsSeID4gFQSO0zSwE
uC2JKEiB3iJyvsorsKIUtMUl3WJHQ6MnA8AJmDs47y7mNXFPI5G2nNq4XbzzAtL6sQnkFJIP1kNv
/07HEUVoA7GQ5yLiJCdcU1kLsJoKW/ZbKXz7xBh3jbvRtjCkXSnwFPq6hzQX/vUUaJ/edDFVV7oy
uUYll3Ae9ALbukG2AM16WrUW36Zb6E+ZcfcUSglXQJiPUEQpyes6q0UDd7x8pxOyMghZTM0bpllx
5OvZg6VYQOaY/bw3kkCFqq9PKAesG+23PI3pMk7JmqI3THGFr3i8FrrRlofcSeOJvWYuVXuwuBpf
gYVmks+a/M5wwO2dFcdIX0PvZTy8gmhsxxUkx2oSt8/42AhFIdo9b2jLJ7mVLadpYcaVwbgOyS0k
2+d2kWB+ubE5lJJMraeY200YnKZKDAvhJH7oAkKYA8yoCRek4KN5mH8IMJb+q8iZvAKrRnk5i9iz
nDkN35Fbu+HVJfi0jnLodpjR0bCxkmAavyGN7GlrvSSOOJ9IAEdQLWGz/4odEkpoMZsY9F+W311Q
cjK63/1nTxXr7/ZFdYIuxHlnXfXqHY5zO1rotVUuvZBWWNWfzYj5lU2EMbH4S3Tz6Or8TX3hC+hn
sKcgjQSdjVxsqMY7j7q7uGooiUhs5ie6vhCdhUqCQLI1Je73c1nEsN9f+SwBpv2AFpK93JK4ooc/
khp7+5vzIFE3sxO7+5NNRi65N2JT2rrtSZPKSd2q2IjgdlnY4y0G3oGeBGH+VZl7oiNKPuRWVPiU
86tsv/tsFPhnMoSad9YOHoHIN4XLE6pF1/15UWCm3dUXoz1/Su6RbeW3iQDZI6aDGt1HP3KexnSN
w9ezrpxb/AuIoz5uT109yuIRaO4LZDp6Vw6GgTq3HKRLcFXsXN5thkzThdocqXil3gTujv1ndQY6
FhDMRXr87gmealgeTlacF6TQjq3vIhWhe3PxDNaB263U8PTBUZo1YJiexmqilcDTNLv5kKuj6mUL
HRj7cFuEeI4tof4Ot25YyAlnKamsX+tKVqFcj/v5X6NtvygCFR6IUYkMTZzFUCw94pldQS3+WZpi
KSQ2Rv4A9kG0rAnm6dKmdGBF+eLA8/56rCMQ5dTRhgHtCBpnYQJRIXIVgg/avQd45ULWNSTYyW18
y4uBQ3n+fwxbl1FYhgRFTXEFLVdY9YR35Yph1LX8yETakX+t/ScHUcrYxXxJbCBX+CUo7QSvN87r
m1suLRh23HQ9QSCaVgJvppzYfS3SN7eMbbAvuMzzbiZtpHUxkZnVc8Dt2ceFCoai+CyU7dnnfXEo
7yjBa8ckIlFLJlU2lj8Jhepfpi3wnW4+F61KAZnrA4OWiFRt8LAGhAb3ehNMJzIdF/T8NQlK6A7A
1s+rJEFpLZheGn49NhzVcoV1p+WU4+/ubLUvvARP8Dzfj6nMM0ZaLQQVV6U9hxVGAqn56cCy6Fi8
/0za28VBxAWRLu8TxJNwkDJuqvLI2dBCiZbk7LDI1S1v4VMe+qBi2mak8bBK5HYsjvbJwD8OZghY
eCFI6AnaDFLOvcf69egljUhRNd5m8el6TlqHpOkyDd5A49A3tb4WdX67t29yTmjpc1x5c2ZsftN4
u0rzYneKErEeqJXpxci3LHXBzcCC6Ge4LOGDU2PIM4YzgwCdSg3ymisS9Wgxqnq8dI7RMetV9iZK
y92uW29h1B/kwXVNmgHFGPWoE+GQcu1oTEIofSUrLiZ9nVRPOzF0UcFhBmEyuMQFA11V/dsaujr2
DCd172gSZZ+fhXRJWcRFZvkOZDPoAmq4NUn7MBRzmD3oXwA0G9jRL4sdZNM6qWiApYskxBtnK6bm
9vHejFZq+t+Y4UjXbgvhbVirbAhe0pbVU9BTzn4m9J7XfFOwvUxOavxbmIeIDNIxHO0RWIAt75M/
t9CfgPk7m+bTzQeouUjgF8YButVMHq1RWf6YAYzk558VBz3lqsVGBOP2QSdpeGZG/bbNUwFEzWnl
+EEw9xTG3MAsUBmkRiDTQxDFF9LR6O3MGdR0L2GRtOKGJj6bfF6mo5RHsv0GBoDCqn1y35BSW7m6
YWFrGM9Z5Uom2M+/QGZgdSbvXumSg1a4o9/DZuc+yLo3jx39nTGLQvTl8SufnEh6JGKsvRDomJU4
PMOJZgr0uX+W7xsM7oExR40NK8ptGZcx25YHD+CJD66kDxYvRV+0HqR+bAUNUxUMNq5elL/Pppnk
UKA0dF1WDem8/jHaRxfD6+/Swxq3JNNPMEM/dcaEwfu58mDUIfNFdd/7Pf7HifUdOc7bVrKGP+TJ
rn5mP42/U1o6S9Hzq38NW0EWg+VCUX6MZQne2QrHfVU/D8P4Ot62KyVNGmfhswt6G8RoYoJExmNW
o/lnt3JLALMWp5rO8VVfyGM6MzVM1eD/7stny3sWZqA8bg0a3dqAyM6RcFHQyhGdkKqLPOO/Nc9H
st3twNFzp+uu8Q4HRYWbrR5xTZlPjtEMV4+E/7is6itfUmx2v0Zs5HI0ovcTYU6GfUU6am7hanCo
PE1hGXIYHtLvHPArIXN0pfLvMcNKBdNGF8B3k2e4xaKbX6q9a/QTZkMck+wj/7Sm8JYsbPbyzT/1
YrO3U4ODik9QjXBl8Jt7mXMuEkt8tmfJcEko9Mb6DYuKkJqARb39Ku/Jm/2/57dpmi0AW/8az/Xg
p7kbb2oAkH+UEWnqF9pzRsHWJtGHEkRip9/yHMmYO4XshcIWa94saYojtJSezpQ+Pn6iiBgB+0Rz
D9AduMcaPmwPY3eNNELYQhQN6t1wFlx7PLiBKiRvj4oOSHbl9dkqQYH8k21osood2t+gkyB2g++s
hheI7Xa6beISuB252Kah33rTFmShhw99+dhuysUz0ZvhSbyfCzQ65RCNHMWY6icZb4Lcgi0gimvf
bTApmm+f3cWmX6s/jVFjoyPNfknnTVcKCBttiI4Rx7rdiAPwzE9RM+dwGNGqCsKUjEvjzTEWdYoP
AnHYa3i7xWyhNgD9eoUkYKDGUDxQ4Axv2uTLzJOX7Qt51aW96qCmqsBDW8z/uI++Q22VE/QYA+NN
Xtmnrf1lAMHyNgxxuWLv+2fWkRhPTF9dKrtlBOv2eb3YrrVDnz6BvZYei/iIuXsKxr1hLw5+tUpU
Am8avLMqj+Yrv1jJURPHbxArGBZ5fAv10wvAYI8NgJ6oBjKl3S+az+XcPhlZWmGqdFKb+Nh/FfyW
MiOqQtHkgq4kUJeJHCaDIrH9fKlhg0K2ubPXR6b8zNkCCei6/UfSd7NS6ExzvFaZm9hps1Xll8mv
g0blcuBe4n1v2bRhkJpKn5haCXogghAkJoWYGu1Hp4JWW2BRhSE0Y2LMR7F3j7CWCfhhBvEB37ER
Z3pSKsTXHniCv34NA/XUCeKb4U6lbPEvWcGUldpNxThdbNpUWD6JaNU5BvCLVHEUkWqm1UtldANe
KVoPvArhuhmy6mBfTv0k3NnFwBjFVyChFn/l1VncUupG3l8KWWTkaG53MRn77BjCQjsvMsuIRBR5
SJj6IgM6OaImvjaYnRS+j97Dye/2hTptsI3ztNOs1IcNje07TCBCI+a/fZrFfYdRgTPvcBKbkm3w
amdlmzK3x4CZun1Mwq6pD7X5fQK40IASwuSi917yZGLpV/GMca7aaX1bB9q+OVt2zmZ8iE40KhpV
sNmw5HRC/vCrkHy/2mctr+8vcXHfm7zmxrRUd9q3ViZPPTZVxtyuef39souTW+MYb2K/8himUSAF
QLPDevafEqmD6RLYtp/z0q+cTgH/rpSfTkPMLKJM+jn0V4o/ZV/earOoXduVBcJOhG6dQwXt1AM+
UUatZmo7eW1qWcFJodsuPgyI6MBhvVPk45y6uy+O9RWwCf4mFHWfGXZpXK4waQM7AsRbtgI1/68M
urCUJR/ebLF/IGSwJP6HcB5+WpN2DPvjGyaSjtVIepYaXyqMNBo61sb96Ke1ntpNfOC/1ZGbjbr/
x4SRKD9TLdIXOJgv1BcsjYXx1Mc4nf6c+SUkgPLYCQBhYfX+i7IiUMEMq4IW7sahNZNDpQCPxD1E
32SayFUOWBtVO2I/IIUXu1DDn3uIVhe4MaYkxpWMoy0ZE45wmq2pLDsI9X7FC4fJdyHwFzmvJJH3
TFWmSSJhNc2rPhOjtMpD1mfQbNa4udn+jnx9LEhBZN19WeQCiVst7hf/pvaIPRqddQ5ocJiyti4H
8ZfxQs6LGogYFCfR4pCmE2ZPtuSsc+dwFIPTMLs6meL0QQPD+6GmjIxfP5ZRLI+7h3JdW528jlea
TvMogwcXbb0ulCzt0u7gXVgvOd1yL/virC9osIX0KbxyLpBRrdr2EJseMtL352z6ic6OBXgIDeN7
mn0tfwepfeIrRfP4626jnafaFSBgn4bnWWMZl2jeNjoe1wMdHS2ZANANeeQ54ZouDFkPvN5waGj1
ZPC/KdMshcmOY5kSPTa+JHBkaKt7BS7wbuiiMMx0UHjYqD7UCYcdPbdDoVlAyjASeQL8yc04Et/o
999XgUXFvJLEDR7gs7mYzGa/JmQaqYD4+EVBIKBdoi/jtQFdBNyG9lu6RQcKjVbzkM1Q1yBxxMzP
r5Sjd6kMlWQw65ffqJ3I9Gqe+1+/Wop5Zl+s+EG3XFJdVwZcm4efnuUKgy3cH/w6GPcghsb9CrCM
omxF+OBJgZKQxzoXp0U75YOd3dyr5EaiYSeDWPxJdcEOaPR7aujfASA1tG5eCGc4l+1ghp15oF51
iLLjR89FfdP/6E6qMFgm+jsHVzhYW4WblhBolzGpMF5h0t/l9n8VI3rFzgyFfm/7Chy8oFSHCXFp
klLEA7QNYfZXDpZoxn/aDh1Rnssyc5RvzZNSh3IzsJXkSKFqTg65GF044wWI1UtI2AprgwM5uq4J
WbwV+6HPa5IPb+nXuGD3xo7YxPTCiRNNeyFYITSqvs3rzsh8M8yqohLbnz9KjDP/KwOszuQNZTge
orPnx0+5+Iyo5R97YUcPHfhhYVJAlpsWLqH5N/3jOjiPdofZ4JqTGBO1xHkb7WnkmjqEVzhaghi4
8HJ/rhRIZ5LkKFZ2k4VSx62wpz5MAsYgFFSAWhADgcq8KSgfPqTx0eqfx/NLHfOcr5rGHtWPNqoE
gcpYasCP+RJXG6hzs9keG+hJen8NJ9xeS9uDGRG4HTN3yqiG4Ngqt1bD+mIHlWnF92VLmtzxAkxx
OJ4BloEqMhpIfLr2QZMYKweZI1h5ohKN3VEMc05foaKJtSmEOMkGKpmxnDHh5B+vy/fIDeWxfsWt
F8fzw7Z/HOnJ21OIp/Xm9H0Wj7Xb7OpztuCKOoOqAZqL+EhGuFFrr++nYkHsdYTTwBxGgAL+7CRT
Uv9PQDcqq+9xgujiSBuhjVG40mlepZom6gkCOxox6XsY0qO060/CkZF6c8CYd+gXNF2OVwS/3t4P
y1ta+ZTPvhRB40YygVS+FlTSqXIOqBWh+nNo+Nub/vvga1tqY8Za/08xJe9NeG1zqr4YAhu3XzbC
+5BsgcQh0IS34qChgnFXBPVQw5suN9He2anFqDdf1O9BmwZmqW3x+dBmlhe/gaNwnwnK4aCQv0tx
AycvHknCFHzNEcakGUDqejPqzMKGIadbTBWTUoPkAp5mzgRaaYnnzoHHSRZ1sKJMqJmLzYzeG8rY
QjAaYg2AmTgZ1korhd9SHdz6bfJQuswKcHD4FUq3OUhYwyTwokTOXc45/0ptn3LN/U0mn184DWAd
r+ScNL32D0zSqoWR+a/kHKRlEHuizFiV6sTnCAQWSnnc9/ZdD363hFAReMfrWiD5qcFqb1url5YH
ARMgC/tMHahSTRJKtBrjqbPk1O4p+LPG0Lobqorvv7ydF0Y4TAlXOcEy26W5FWq4o4wAY7b2v62t
dwQAfg53vjSCuIGXTqkWuGnuZ0ecxZmIXxtCvf2qN4zLCqfjjOcRmieX4ysfLU4uOP1K5yjkB5jN
afl3DZB9fgA5beveykOQDnRfmKOd3Q6lppkQq3NlZsW/KqvaLeHW9240CRp1EtlnMzWuVlURcsDO
9uMA33kVKoVBjHTLI8X9WhEBLmvFBCy/X2E/OHhaTAI7U1K3a8kiYY9abzaKCFMLit7hLMuNhoQC
8sufk91HQGOZgFbnryFCI76PiIaxCo/+3q4oYFonoePTZ5xtW0sQ1eUuDaJbPCD4nEXR1ZGxbKOi
I8a0A1F9xVp59mHmyV0U4XVX6JHMRaQtBl8KzQ7bn/Vn0IM54lPqy3EFvaDBmenDX4zeLB5inCeQ
sb/qnInXP+U1kqMjoBbaYAITc3XyqKb66/eCC7qAa5rcZ6P4jneaj0j0pQ9G4p+nhvvOG1+t4eLK
zzPPR1ZfSG8ls88cLjKDcSEGASjUq2iZfQ/X3VN1DljKOVKTJe6rl8rQDAdwaIQe7ly1Vu9AYGPk
VzP6X639uh88bCYPXBWdkiXgoFaZWoZFjucIl6K5+ktZn9ILyBuaCH3YbFl84SlINnsxD7GYyjVh
qsFp7uCkEG8DXvIA4noMm//PufQES1MjEO2b/hOay17F/Nv+g+7VNNbzWJfw8boVwkRnTz7EpsIR
2uA2Wbx7KxntL57BsvsTl2mJtLeivD/ZY877lBbgZksNmVIIYVSBJGF4l3YGqy7//bsIlbOaw9Zo
stlo7+MUuC6ViN/HYOCfmssmDPbSC8Pn5ctjJfEylg0mEjBmDrRPUvTKsc7vpH3o7IlJsZMMVifV
lbZfZMPDVzaPO4JdWJ8HTe5zbdW34OJvgmyRMN0aqBb857mcQSBF0n/fohF0F/8O7y+6E/435O+R
7s5qxgAoNkLJeGjFapNEw337u0a7oj9m4NqMJkY5fnE0PJzfZkXoXCa9/WLPWw6I5sZombBfzfC0
3Zk5ULsMe96rxHwy4UZtTvJwImqOTBF0I27Ylux6gZZyYlzpMYzzzycUu7AmZGEupMLjXfZ2o8a5
OYm0c2mmDtL9i6pBrsZN83JTMNd5UW3yJGpyr7uNMEWQ3uGPwPfErRxLP9Yvo+nTonLO85J+f9OH
LkRvGVf/mI38DAox8l7SUZDtoAunxr0ZS0JrlmCozdm6uW/oMr0e1zXTPlmHalfwgWpfKum9OfeV
faLeCsDbZ14IvcIVH0d+p7EsbgRIxWFTWEBvCzRqbrjE22zwFoUXy5CXBxOrrnbMVP1ho7S+iYau
nHw2hf0vMoRHMFFhJtgP7f+lt04EfYxObY9ERynjCstZxib4zrqMb5m+Ykp1ewz6FvCYKgdCoLa1
Q/QNXcGZ+wgktF1Efm5u/jOcY7h7sqF972jWinULQm5/MFY105rn+V1w5T3k58GrbsnxrqLfmJRE
bQ6oG8lGxPmKk3O9EWebEfOzBAA/qEI6H92xGKZMntK7QpntAEB8eAo5G1uyB3rltx1WFsnPjZRF
EyKevaNGkRP7T+eiXPWkJj985H9ibbQjqVRRf7Rz5vKwUjT4Rs1XC6IBZ65DzM/v2QE/gTE/KwwC
dxG4lABj4XQrOVAtOfr5J8T+mpWdTynlWfNXz2Dx03xZ83yELO+3FLeF+mN0fgCgmTjjlqQ/Sh7a
vDwEapAa26OsnIHrMfrK4YJxTAaTK79g1km9NreMrSXRh4HIBARcN7oYSbXdxmPtyOeNXZR1VoNi
RVly2gbuyMsRfssw/ndDzDbarKHSqJYBdeS+Rooe2Vxlntdy6o0Amt9DgSOKH77AfVT8QPXAMBEz
2UMBT58KQ8jH+q2GyMtjTU/1TXRkYbT4RxOywhV9DJnFkePnG0OliwZeHxbldmL58C4KIW95BFEg
jTsP95nGy77ADlYwI4Hg8kk1PId7Mym30saE43LUjLQ8/JzmGz2iZtvep+PsQD5H26g383oBdE32
RURJuj6NTlSsqCtoh/vwY4E7DCkwCKa1KhDM8k3Z/Nn/+QDUQG6shkTLoSSrwjHDRPa5Qi0n3PZw
cQqhzZ0vCrnvGi5H7rHliSC/19hn2DPkeD+7JiMNBzn2O3BziR8OqOkobx17sW2oKDYYKQ5WR0S1
Nat1cZm1Br8tzXMq3QRsUfKzaQmz877O8knnHc0GRF5O4FE0OjY9GnsyK5zF8ChEn3wrK+ylcN7J
yd4zc3ZW0yiyFxPAQJgQPXngNwxnayw+X/h2DsQgxap4mRq4mGa+I6i1BcO1qiRHq4D4Jpt3tfMf
YzIiLC4YR4keWsy+kGMFu2YNVZ1VXtCjtvWFjhVAta1NEtpC2WH1KOkDEGoVCGVOyvn1Okn92Iup
9DDGgiaTKLV/W+PxA1+qDVp1SOk0IyPvWJ+JvuE58jNZTlwhs+bQeVx4fxvq6B8W/0kFBCHVZiaH
r6HyJ0uRpjRMSURp0YVkJvWulxL7sw1NZIHyfZsPUpRU/32eyL7EYPtu5n3Qf6njNARaGtGMH/bx
MowrfpKcUXvHXHrJDmkAHqukJEVL1gFt1C772xNWVu5ZoGOUqSC96cF48RHPVp1vQw9Rr5/RjCNw
tZlu4FPBA3+cQ3hEY27xGD553TvAXAoQrZEVtrH9YgfQkm/Nq1f/MS1BrivbHIhhmK4KawrC3wZq
D89vKoVyGnADPCRHmKpR37TMNofVU6s1hZyuhCnj6rhRg04TaRtBpIeySRbB4WV4+NexwZ+OlTH/
5H5GZI1lObPD8AVerlhU3VWbC297a/nwq15ZIdCBI5D8KjcARAdE8Z+qXXuQLj9pV7IxXLeuIVQV
mMt+MQ6i1qJBHykIZnFVokYdo3yYgQV6dpnsTBIv9p6b4WH4OZO0+ctbGhsxtVru2lNe0IrAWewF
PFwrakr/RfIQugUMBHJdr5/QuuFhLq+3DjDD7J6FFds0AlOFCbq5xnbvHWFC+/16lvkl5yFdtdHT
3WRWlnqql7E03rlYktQYtjTyayNC4gQB0/Twz7GshezUfwh0qTD5aYC5E1cHwsGclcLJz2y2ncnU
jJ05bbfIrjN8xvQCpvVLZRN10BILbyoM/aT55Sjcz7eEiXi3QgcWyEdu45P90AucgKdH5u3Il3Op
Rt8D6H3zetApNiU3kOuRqNqCtxYiNPF+wExdmsTnEMloCDiM/gq8wrKfFwK/bhdb0ddElpB8TroF
HinFBkmlaSs9hGGijnZ3hWuabFoyfTRqugAHy5u4FB3mTU/yBQIMXcxlVroKsC3kOXgX5IvDOhh0
VQHGZ9IDHQkj91g2trHRTvmMiPTLbf6nIWG4rzJhew8RBOfCCK5jrNHitW4LH60niXyDIgV2AGzU
oeVjeNBhxNbwX9BdZbpz4+s3fGnRsnlqPWGrRC6upwPF0cPail4Oyeow1/DOdE1+fZl5elD5GYgR
I3IoKeOtl7thpYFv4SQByK/edutocZobo8VaUU6p6qheMHSn5+v/IqaHm7AyCz8hkIe/DIm60D7d
+IhTiucuwe+hOetJL6kwXlDhIzwLGCWowOGYDrNHyEtp8HCxXTe7xM2iXr+376lJuLxLFOtBMfw/
MLJWzuj+9Up5hDfCrGUMkz10k456ibOuV8PZoYnb2B+uCH5PollT6KC33n9o5Zc6v9SiocDpRB7A
WzrVWhR9qvk59fL4Xks4euLs6T3B/ARrMVnOW14jgDNcu1ymqyXGb6bGpdZNeF17qN9SBA7USLlX
95Oye0JBTPsnyZNdg1zpw4OEftkbIn+BDuDfZWsABDLxaWgiWSKdZzzk/irUbZA06RRIZTEzWby0
mWtEl6VSDamj4qQgluhiXH04ph1RdTkvHKELI9rRJortJV6s86hgRRO5RHtY35mQ7WRhZ8Wz7oRc
qeXzp1VZQ2abFHYnqT2bzzDyowuRacCIaqhng1jZ2aH/gL5D0duClj+9HLAUP1YDFur9FFurbQAo
CO243eeLwK8050OrnIn9EEOPXnXJ+qJFKnbIIt4ir+xVxNSUm4Hk6VNslBtQMH39nyTBd1F+dRIc
ReJI9SjEbosMrw9kq7mY+dq67jdyC6MqSD9fFQIaJM9WX7MK1/WQjYDFFlAdRiwZz4G7HIShedHj
sfJf0vqKDm+Or+z4bXwi1RfFH4fkGuGTeFc3kdoBxseSllwA44EDz1/gst8CQZjRfaZPvZyCJ+uh
DcPQjYRQf0b6cwKmcdOeWzRT3t2Xe6nIVq1wQvb31RDbUOAbYsEVSZ4bfq1HnJDqrWA7yBxCKcXl
gWdURe8WCo+qmXOIzoolG9zaE5Y1rh8+c9SE0ubDCyGdAnvqJUz4SbJXQxdKloWdgA+fpZ1JxZvQ
2UvH7gZItkyFWK8LAhOWCkWtZQ2KBKvIMQ3nKO59v7gGTyLgE0r9sIf4WIxFYTj683kfjGSQ+cuF
muWPNSPMQ0vtZntoNQ7gbkogntT9Cy7Ptt0w9JgXOswgIdU568DCRUXTo7VuyEgsvH//ciK4Aew3
ceChdK1MztsX6A5mfAAON3BFumjONQgXGWACyBc4nAFH3igxvy3QosK1wm/XKZGVVV5wPbAXAI3W
QQfPgx8rrlMIGMiQbylYRrgQkytVwrMSDbOPGzY6MSaCk8EuZZAKhL2YSsLov2hiULDKGIMyMfJA
keVnrPvetsa+L54XSWj2XWXc97OisYQosPo0JBIVR+Hs+fGDKYsEWPB/0PimCx1DQIZ3ZOSdsy/3
c9zjdtC4aQB1uoa1tj8JClbURFukKqMbrL3sG9+ZpdsIiHsNScLKJE+8Do8AssMzmVP44S+dd6Vt
Lo8Kvg2QLGUBlSb65LVKSO7UCQZckeDnhouRjs+JyM4yVB0Ggo0p5Y5pWt6GkuBA+Lj1nB6BPJtH
1pc9pZJveLou6f3cKjHTJ4pV8PosaqUAByI+Tqcfuu4dbwoWZMQV3Plw34vYOpJYPpMdZ/Wtwmrm
3URFN8uQfIF0iII2ei4SQEE0kKfveSrFRAogAqw2LhdtSnz70D6gzwcChkt1bW1f11GQnjvcy7mm
wHjkjiVUKYm8F8Q56d1fN12IGPJPgr1Hq6UbLfPecbSbcOnA446NxOa2tEf3OScNZSXZo8A56fw7
6Z1n04z+X7DkuuuKn11VKrJHZbLVt52zQjoReGRgehOkrRnJrN+9znq3vnRCx6ZL+cAdRWsxdxI/
Bf2vPSioYWEBJ0BrQ+BaCchcKc7gQqiiKE7DI1FJxuJ3oK6blAehF7s6gYdL1nBLaCJyHDwV5drJ
IWg1n/S78CEhdLDVk+YsiWLxSgAleaahaeek7ZBd/3IVhA2v0QpsY0IaRp6UWy46SzC8PqBn+Xw1
VXGb8vsbU5yTX6oEHgpR8Ah2vtrZ8m0SBzjpF7VYOT/yAroAyChpRyZ8d3qzVNPFiLv/ITXgbMes
f2ynsIvfTpxHoumVNJ+nRnxWwmy/1D86/SbFcj7tSCSfznlr42V2459LudFXjIc0IDrG0vwdE33E
NveEgMQDEF+mzWceaH807h5HajglSEQHKhTL1XePPYXjeVJ1KVg3fN1sMpYuJrsQzn3+gpmMI9B1
T0CqhNy5/tzrNy5NlWVzWvZXGyTg7vQ0OKDvw4c5fnew9T+pSBJmF0N/yPFae4H63Jx5HHVEoFtl
OJoUdcQl+ZjfXdE4umyOYEMNV8wofxjddPiAE5D1rKVvvOE6Xa7UOTfH2hEZ6sl0o+nEEryWAy40
zQhCej4Bz+KKdbPIfbhV9RLpm8Nlz88KU2BfI5Pky9NMhdKkloE9zmlQhBHaMqvs0k7QFxOQg55A
umBrnyGs/v7YdT3mfQtWTk745Vz5smWk4tJfRZRot+i/gGDsNpz2QTXtLbzbwWQghS1hD26WM1UV
pM4r9x5urX7qIDztZcUCzSHTnlZd2M2dGPM25QgMbo8AKwag+8ZbC3QBxGAtS1dtfHna/2ObBAwC
bKNWsutbi4ZZtwUmPlcpzIgl3BNRr75/UNVYcnPg4q0NsC9klRxmM0AVF4RC47JTXLeJmgiZ9sk8
qbcbkf83fvLOsOTKBEuOx5huGTHM8qm7vxEw8fNWDGSEQc9a+pdnE353aQm3lFg9eI46mUwPI0Hs
DFjefcUEYGiUHwauZkx+Bep2hFdx4FnBL5grvOCt2vib0UeOJU8PFqp9zs1De9JauBAJo3xrxHb4
K1ZfgNWHn1MFGHBnxipuB6XEx5XzxYJy1vIfc81NPwgb3sdtQJ8DPHarRiQ0B4mD2WnbX2egpC+Y
Z5l644JaPNXT34d87fHIouYPK7wVa2cS4v4CizfBKaVHhXfXlZAkID7qZ+Q6KUpLWwClI10JKru9
R4sspAqA5BQ0GbzznxSqZ9ogEuITQnZaub4woX3noSnIhNlMHZX/XG2GrcUIihEWbOV7FyOridqG
Ll1ngEh0ODrA28sSoh999PwpSGi6z06k1yk3tGVSDspaxv3czWbLmdnxKwCCSwuszjJ4isfFLUk7
EqRHt4FAr2JMb7Gnxdgs8rAbOsQQi7hwJ3Keb1RqahWLqB3LqtCmzncs6pyTYZufzMs9KOJTX8Sp
gwgT0iK0fzMxgr8Ln3dZ9aKrbrn/eUQbQlpVbySqm7UAMB0HVukcOWhJrhbJD5qWIUjErxiExv4P
Q03Iz/MNxPiYXMYNS6fJ+d7LraO3O3UZgardnCaTHne3Qu0M82NQYbu57PJe154JFi0sDRx5X2Bz
Isc9druF8XECtSGCdUM6tIyqsvWSnjFm5waoXWUhca87M7hIEe8ku3soZGFzbd+LMN4D6+5LWQOv
LAdz78MHu+diMclalGn3Rjz00swR+ItnEEE8Cj4OhINr0p225dbXySz81PQcShAHdbU2cl6fDuRX
FNeet+AbJmgArxLkRBLBwG1wWfurJfsiXfT4LZsXdL7sezszLy644B+JBo+Dl6j0BJN/s7NuuJBi
uMTaXRgYQUoFpAcK5SKlCNmp+uEnsY09HHpdCux4eug5n2+Ma4tKs12aHxgu1mnMCuhl1a5oeHzp
sqYisCxE4u/gHfkr7eaTZEWwS9WAMVz6hh9UEAaeZ2ehdG2KgUqYlgvirPpM/0UKk1xcGhPTRDyM
MC1QOij/KccF7z3F14skUdUQH2gcx5ljyD0BiI2vyutOXVkgFJrBLQ68AaSe0VG+ZO24ko2T6EHl
wS2w5LNr1RG0Lgbo4izKYC+moJJPRy+NudsLixpeKPXzARRjwcO17ROb6hgQomd/O3Ls0wfxkPt/
kkn8U1eHRDHj2c9Ppy2IMZd2I9k++Av5HW3jfxsM8ori9DDFZvQry7XS0RUriodkBV5uUiqC3RzH
ocdJaw7IMIV06J0kJn2HnLvW+cyVbaAUC2gE2Je+i6NWFI9s5sUrasH76ZoItaLOZEQh/a/A1GLw
OjHR/+RJt1nQ/660e2JU6DFpfWXcHEBK2+y9yEDNhkpC7dXWupunnOXR13KFSgy/najvkLGc1l9R
7vs6FkdYBo3hgBeDxRqvjQr0t0k78WnID71KY9uaDTJL+IYnCYtWRucBBsufgTLB1+tUmODaqHUx
O5gCMUb/zafasrRV19IL4xfq0PUh7a8w2fgluEWZxMETvHDKoXNxQGlYi8RAx4DdpEXf6w7JIsSR
LCukfS8AKNpzI99XEA9ID2uEOvKKPDFcAHG0YBtW4D96SCPZK5BZlXjpK50l/Wapnq02Hli16s02
NgEvPK/MCrMOq5qKKhhh4xckGcV1fCs7LnbRY54Z+jOCSy/D93k9LWWfznnJX7ixtB1jxcdPb9K1
ii3UDlECAEhXQWXulu94aAT21mV7NvoS73HX+CildqgYzlaZu8eg7EHSdGbCqeyabYM2duLH//UH
A0NzUXpmjv50LeUqCC+01s5M3SkINwSWXU3GRZle/mQsfNaBGbnmXznmopY2hx7WkRu3MJRKAMrQ
u/lReluiir+kI8AllKa/UeQ8A4xXGu0Qwh3SKM8quLa2139h8Fd+shhrpEF3b3k/Ai2NdErOh97W
pW0Xs5KU2TTuaO7Tfd3Iq5wvdfffwi+0/31EVk+I1Bb9BYsnm/LCtbV2bLW+744QJm2Fvb1nJczk
d1/UgE6NS/13qgUriLN9C4jAS9dwZCxHORccxfedkKVF0WiJN8ioRHDfnx+6vBJR/Nl2sYR5PBTb
qbrX6IZO2ecYO5VgcploWR/EcYO2bjiOHC5SJpRf4Ch64/sh15RzPlKArjshw8ls9LIyovrFqZpB
zdnII/FJfejfpAmGPgmk2Har5pcKBiUYg8KLe2VT3WH4o4PIid4pr/yXvmfICl6KtEr58FiysxC0
U6P+Zw8eVry+/Y1nmQi5tvpwF421CC1sKIFKit/e3IrRqsbbUn3wVTSyw78MDREKXU9lhnCWNj2A
Ly6bc+WS+YavGDBR+5L86MYsDy1DtM1iCDTUEUr6mbObZe8BQiyCrd2Xp1MW6TTX8r6DnS2ALYem
/ZjXGKZFSJo4H1Ii+B40aEe6oHjp1NhNAKz0XR5tRnVt/dcE1+HSzg57Fi7dZVTd78a69KJpUf0z
8X43J+/cIcjbonEvl4jd3+K9iihH1VH+lQ2r34Lv2o1FfNxsQCFnfri1vuQ6MFCOGwhlXY9njYNO
U6FD2LM0DR8d+kLwi4u12Z2Su/bTEiY8XFAj3wEUW4sMPdnXXjG70ACtgJF448Uy+e0MX0Z0J15e
Aa0kKHU/Sz3jhPcah8ZGNxjzahJHY2U0/IvPvOr3vyOJWwmpi3NC4WWru4VVtyb+BE3086rnSF+f
LHGZTmyE1mjxJTsUo7FqBk0KDZ0agJ88U2nECZuotWj2hltYrS5DHODAnQdphiR1r0Ccc0ulInXW
Xmsa0vfbijNt1KsVKzgUp93llZS+sq5fktxfmLJfuRjVYdMm5/EIV/Jk3Q9sWpl13GR6qQUGfPIx
rrJkQtHD2+UO93+qPdoHREU3WX1ytTe6ANM6mhErPkrszQ3FgyfG0s0OMbTZhrgFgb0fIwfrgUO+
yaTmTae9NpAfDuhIgrU0UyNdZo25iaX6O5pT+AwMwI5K4W/2xPOQAPzwFNgJyqzpVPTUsw+Pbba2
rPAhWIKuVewV5HQ1ePtjG/wFn8r89NQpLnufG1KJpGDIzOjz8sJsgpSxSMkTj3TTNmYN0Qj9TGu3
wC/cggIP4ZSPKHCOJsOk9nORSS6gmvVVZW7Zg84ZHK3pZd/5bCdTVFROpeJphBRXi/F2anG0RKOm
+v/RP7eAxCKj7OqDhQyJAsFrypQXOhSTC0cp47OHzF+YreaJMWWVuL2L6b5esJ25m4TDAlwFIl/+
N39Kn6WUjUtcelcvoCXelr2KJ2+ohtyjRxUvT3VSx6QNCww/gTa/a5nivChyd/CYoUJuZwaZor6Z
geBVoHZ+cb3bwzZ4GOWtTJZOB5/x9poMI7tePLl517mmtN4w5FlQcf7abnTn3GmMM7++dR6vwUwy
al9XDHsoNWyj8wd1pnAbi7PBC4wu4ZdMb4XiQl/WLDp9tSFjuSEen9DwKxVh40DanLR3Q1iEZyO+
dPaWb5DI4Jmk8Ecf7RFOoykfwOYWLw0KUA/wn643XAOY/icx+gnCtEUu9iiVs6ON7irqikeS5yiG
OHKWk5suSix0B5sRbxbhOXNqJX5Cd3STZBPqdmGtR/7SFDb5Lx+P2Jx1/qhIaf/WJWRsKND7BmxT
LzpTeeqMPK9YTx9RWYeYovOA5g4zRSmXUmpR/YVXFQXkWcEYYfq/nF5j5OFuEdKVcjpT89IIgfpd
v7V5Hh7211MKX9KNIaoCaL9qe/tDzGGq/DFya3kU/PMMi9CkNNqW4+gSwIHgzvpMdf1I6rtZTqvf
W+sM9V/9x0HaySCaYs1ScE2Pwf7TYzME6Q0i7++cY0SHT3sMtFZ6wVzmeUA7ly521Zeqchx7QRHa
IW7gSMvi6RB7kYMjXohSQROxYkIFyiDD3NosP4PrtjFBkz0tl5U9KoKS4Y8QikLBbOHlebvrgpbB
jV7PxoQUMhKBK0jinzsigttbaKmFHcY/IwpjhkXtwm2lenQUDSd0u2LfLkkVM5YazTZksXe7RZnt
9dGgLHhzYXYkPkem4Eof4U/Am9pJcnW5gaZYq6Dj20fEneDAOrJ/lctnCnYTThFtGtsWu7B4BDZD
If5qvP4JnQRpFDP4C16N5wEjo9dJrFZZ4jCCy6Rq3Z0WFU9XjaXUqxegitFt8nFKrbEtzqo1jFTt
JEoy/VRlp/zx2CkR1ddf0V2leYq2vSK1hVETJ2bFo0x+L11u1WXvsVzEvQgzB8AjBWiKEqAFgzKk
qVMu9czrOnkVWxO4nvevM5Ko5rZp6VBOSLms8FQxcWSahkCVcKwIzbIrC+b3WpaF4kRF4GNrLL+J
zBBWEwTYvMK0EqN3iLra8MRJf+ot4VKZO0lD62bnARqVtQYNFlwksWsaahNS/BDJ+MI7YOwUwOKM
uwEYBjzVwC0stSTEwwroZLstEHEeSQXPP9wKuY5TjLpasFihhffeseokmGTaSmSZD2aCfr+TyMJk
K5vRI/D8gkhHsSBnBcmbGD5D9KTM/qgZbDbSqazhXRTeOgj8cp0rtqy+CAyhhWsa1voViP7GbTIv
+Rl4G2u2Y0YupFT1CE6LPeRDnV4YXWRKaPFBMT9K2F5CTImTrVf5xYcvdVAaasODCRDsqwr5cxgX
FV5o+53fAYhGF3Dx1XZFEUCckZbg946lOY7fa5VSrfR8R14JhHgprp7jHBCIH9vT71jqzXRGBjbr
vyQiUAZ6NyIVl/o0vzU/gjGj/Id2uaaD7oQObGZKqeEblgI/f62JKoaYf6a/bfzMUSBdOfb1tLqE
3oSwViy0BttDdtqbcbeSurJwY/7ZcCvQxYmkQhAc4ZHLUSxBDPe/O0rHcBxUE+LMjCXtVLEvxSEB
NWFUjFu1Eg9CwjhgI0fcDGvoxMBnwqGz0LpHKciafPTCN5mzmh0mpxedL7ozGKvK7MGH5gtKMatS
cGsNAppLR42PaA+fEfBL8IsLMx536nbep4M+PmWiga6zwn7qrrHj8tH3t+RoS+aYw25nwiTRXsni
R4azPwtT/06jGXN//wVrYB23g6QMqJNSjpsycyo1Bg+B/kvKCh2lQxTYQz/HN3cLkfD+jOW1wJEJ
J4dzfT8HrHJg1o189gBAmGnBN4EjDIurOl5iuTMElVHr0Z3pzaHQIkVrqKzqjsXDveptX4UJvRpy
pFS9fidFgSe9NqGeQ6uwwv/oidOt8Gq1hNgdux5SKgOgEmCy3RULjta9NpF0eKhwpUtwxZyOT/+3
RIlGe91dmEl7YG1KeneAyrk52txNApzJz/m/VJ3mipHGlZyqbU/oqxR1Y2R6Vq4BJhjs8lKS4+j6
/Ix4MsXfG0r9NaxC9FkBlrmfzqa5Wy7giQTrj7DNm6JqZmv0KateRjj3V+ghma6uLoZTou9iulQo
0M2P/0DSSsQ8qKrtZbJXJ5q2yOeDWFfcKyPH43WFSC0cPhBTDMlynejFA06Y1bs+5CYX8jM3LvhJ
7euaUK14hdzrmfqpHCGeEeJqmGlBT/y7r1UEkev/FIWbAPokMIStlaB3+miX8Y4TH7l5F/BACP7q
JYY9eOlL+BvVDBPPph/+cfqeJxBzsdCoSsZdmUsO4mzxcq4pZtsX47BaU0Or/XXzbPUWqegCCzsM
TM0QJxjZHBVipfUiU80HVyg4WvDb2b+rUbPgYEu/FpQxUrcz9VDcAxiaFCp0GGmRFhwW116mFr86
oUfkGx3WcYD3v9GG2adKP7LpJJwnxuaSIgzJhZfN/Qvtno5SM7ZAeEWl4fuANsC9r4CfwLp1Pusr
OgTc6i9zVpf0mfee42azuUCD8X8OVNJqcVl9OtWmqgKTcODx7YkfZZlYKp/rIftH3vcSiFcu7hS4
Umb/SMi0C3mSa+bu+qT918ebyrwYFTbakdpJD7kF5yDsMq1BwL7dNfyuD3ichs/NfZn+fk5qRylZ
vK2jlzrszCH42K2sn6IonNP4u9LeMnp5iffMyD2vPSbxaWIY89ihajO5u+R6mRbEJE5e5hEiuoga
fiDL8tDk5fz4OPvTKgurF63cXgoO2LTedWHYUCZqACp6BWq3zb/VIYBd1la18ZJr0jibdyPN/E6R
Ey5RoJeZoGxVZ4czmoxuc2sRHb2F/NjBksu7klKicdwiNZYgRiWKoYdICZ0jea5aCj18j3Ew64OR
RhLWxQOv5aoAW08fjpFQFe/GV29MAOdpGvGgq8uOPfA5xsWoouqG6JG5v8HlJgF752JQPLXIB4F4
cBYdVBKLiOpzOLgg7tk/PZUpiZEWz5mPwbcyY9YW3DAR99aawIuAkaJt1UbY1pcqim+IspgAZ0GE
2w8i47mIElSn8V+5LRhlN14cA342oRiYswFb3f9PSyre+39zY7QIdr0/M416mV5Ubu4C/svwgcUp
NCsJcAJcyakifaqWIDidiXafUfIRe9sJR6wMRFxHFdQisY6c7nlCYKSGWfmYXhASNHR0dL7YSTce
s28aCYVe9/PNv0xgN8iP6xTEIUHoeebcy2+G13hXyKKCWm/NZh5jVqpLS5Q2OEn6ERubHDqLkGeT
Fnt0fLBYa6raIrpKT7k2gypPqnUiBgyEb5u/HPtF6q5Ae18v6zyJTIB6tNFIEYGCS6YCzFHBRnXy
qw8AUkCTGvLkNQjD9Mk9FZ+8H5ViSwtLnRazurGxBJRKH7TswjSJq8DJDLJjE8/WbCM/DhATcZot
lzKBGUAOgQ1idsc/1//RiEKKnfhmARMrAJYRzY6bFYDJP0mau4ihW7DOBIk6P+wsDGaFJYRIpC6j
Mv6zKcURdYKbhs595aRD112CWcBjc9PJX31JrbK/Jkl7ACjAGW75wpXD6ZyDPa9TgfR8HsHZT/XR
Sdf4sMuRlrZcjtA1Oapp23kM3zuSlClGLnoWQ3p2+h3l0vDXlDJ3UTfOJyZDSTAIJ+4vlRIvEE/s
l97DTfjPgCPfAq2DEMIsGRGOMF0cltgO6vfmnbg+uZYTYgNNGAC/OLTmGCTRDbZnOeAeN8rSKNSw
zxd73cO/0FyuAoNkWsD67zjmb2AOSK3qLQy1HByI3l4rMoQPekhkpVRbod2jYXCb0+OhfIEIib3C
DIqt5NTDc269n9qV+hj0i2mBcMwJcbVHThhoe4oq/KZlru5y/1QvDD/c21aslh3ZMiDHUJewItJ/
SqSYynLDVb93jFrZ4fvkCd5qHPxnFSWNpHaaReYFmehRNogXuj02TN2x2bxFDXomk0k7z5JUvYJj
smrFtwa/HWw3T+uuM44H4/q42LykgUtGn/87pBriJJnDyBpjWAvRvCQuK5QRKPDzpGNFDSwPSUwr
jxrFcYRhy+cwfjxj16tzsCLlM5w/3nyHrvn1oeh5ayWVylWKSsHyuHzlIuPAEeaDsUbldR4ZGrSy
KXM9GjKfql92sj5/Hs5pEVCL+DJvQ5c4O+g0+fRJeuO4ypzrdGnhYGBKdQXyVJw+o1m8mQHe8/Ev
CNdVgR/y/MFH+BylJZZVBmYAMnsUVL4YNzrXbJaGCmYmOl7kLzBuRYuJvwsT5yEzsuUn4ekNyZzF
/TkNKkxetWI5B1yo1ECpfpdmJSneE3bjg3dCqEDocsuIulxXxNQc32F6oe/NU/rJ/Zoo2grFBMHo
tD8N0a6Q16F/Y1wOI59KAiCFRtpLMYJaXuT4/vV/d7dQ15SFRmmEbtGI9XO5bDmOcn8NbBS9VlLk
9WxjgFW9kK+Zkyv/n/e7Q6F+wrZQZf/ZVmbVQF6pqHL5xxwScHj7yuCUTFZyT6ZNVWIRB+Wsv8th
kYpk629tNVge8thxpc9SWrMe1eiAfySBXTsYcP7d0ijOl1TN0Tp8o4UwXsy/2zoydjyQ/kEmPnpW
f0yFUKYDfQoU0mQTWYD7g4iRnfrThwosCrCxtrzLTFUi4NbhH0C3xn6le3zCAqEBNknKr2VLBkUO
DJtbpCSn9+6UsTIc3h06ZA6kzmJdUj31fG4q66tw5xODLRauPBHlIx7EzgRRWhzpBeX1ppBqbcUd
n1jEbkdI3pBp+Q3bP++NU2NEDdBjYtsIGdHB1wH2I9MWWOjaWYM6+fd7HkC33wftVvBjC9pZv1n2
o3NP8jS/LnkVDmOrnYbgWDUcRrkv9amnNq94MEqhz99bGQN4dzX3rLXfCFxUmNaqc6L2TO679aHi
lBGCBvMYYDzP16m9NVp75HniPNvW2veXmmDXNqUauCzNIXsiOGtsBZ7IZThCZcQGhditoR07E4pS
8+ZgVDqaf+9kMgUGN6EY909aKlGL/rOEa8hdlGo/SMW4/BEaZ23Fd3nSweZgfucsiY84HifNIqTs
9w58d1gQv7yHZiYzlLFBmgPy9oMq9HOlcPVthdEmOXfu1wg+LURD+whUdNjDbKhyZ1Ho7+lbme5q
mjzLufhF8WaCgvaKS1+ocqiVG/TxS4rCfEcVPbbrqg96xh4ql/SnBri3GaI/mguURt+tcIdtF/1R
c+3N5Q4lsw8+cm8NT47AyS3ZybwfpkDSZGDI+KGtZrVkFTxw/6xNSbQB3RxKo5NqO176A9DMMJlA
rU8DgBL0skEE4AleO0QwGFVtuBGNWVJVrHPlU+Bv1CANEMEc02dByFp36zd3n+S6a0jL/trvwYyE
cESLvHrL647GH6S/XQS0Y+UgJTEIGStVF8XKgxrvHqE1kqZPh4Qds3ssPb1ufVD5p6WLpqR+2kEk
3hkooP5tDVbho2gy+ELgvWkNWqOItavVu0PLRfjbXUktjZZ/HiYODP1XYix2skICsYpzs5H49FHY
AiV/8k48ZXH8sD/pZsbI/JwswgwbmySTI0tcRkvtNM9jlWmMTICmeY+Qs2YMr2Zs0lPBDrJb6/Mf
EylQh7/KxyoYwz710GAnAg7zPe0B5Yti57N+dQQGcRevnKMjlQSluryj2Bcx+soZM1H54UVWKJZa
ogdSLSdtIjARhdjmJXfPNM5+Q+7NOQF2f2eO4b7OpGnohZK5VycjYZFhsWO2RaoKCxBkmmWi/JQ1
M8vaPGKmKZANjxFOophjnL1gh2b0NlnaQwkK7dWUx+XkXyQ9CqcoyepoClh8eNBD5Jl0F5wp3H7t
u7Y2E0gh3zxKq/GwXgTELCxcsk8RSmi7hGLJB/dZoLipBpeKOzKD0ImU/L1Iha7UkYzup8UL10fs
JYesOwWu3dLjjxGVDBaUpS2THuiWowwMlEKMx39CyrKMdQgXPPASsGzCOENIOgFkDUyKL9tMHYN3
gNmFyGp/jJMppVpTu6lyamQ+nF1GU+qjYNoVxhLoBvfW1XW2OMyOv2Myj0Cd1ylLM9T29iwtxMF+
NBqp44TJi269v+9tpZHs6s/SF6AGSLgqtxJu8Umb+Qj2z3sztTSYiFswYkXaLh/p6nNaoWC8ahEe
PAtuYwY1Q+uJY1esPUtfb6mvQKArVBwxYQlVeb8a36O94/1tJZdHaDndTfoqhxOuARVoJpRP5482
dONegxb7PcIGh+Kam2fsaCJ0qWjPv6wNDTYXgweyfoE21qx7/w1sX+7odVkPoaR2vi7k+VB4a/4f
MWi42h1P6VcO66hisNCIqIeuqt4TFL6liqrdXX6+HqmKYIbMP2quwrBx10aM3RWBdVLsmgEouZG/
Ojwer+8ITSYhQnnVMNWxyZY4oS5DoDIkqvef2BttkPwsfgYX8z/xLQ4zrbUCbUycY5pRppgOtbwB
6hbZXdzwx4aDjSJeFY8UEvHT1NrH6wkvqyuc+3kyOur5nu7yqCcx3NggjKEg5d5a+NAa76xeWIgc
J+/YN8vlHaRdR29BTSH8Pi/FpeCYScJRUwlgMB7a+Pq17vdnTVY/G3McfUw0loz9ujwmD7FIhGBW
/S5cn1o1qDHUJsvCmA+kKkmKKKnPomXwckIHYG2V80PUj9ataFIBHZEpsUlZuKUWGdTxQOpljSLU
q4Ob4G9kAknGd3T84dIcu/cktxHYC7aqi2rU7b+vAzciMo9Tf0W7QVZrU6mrUTzmB9aPyPh0S3ZK
psc3zacGUxNnsBpR6iDyje3/t9+dsDIBGBQVzfcFmm7Kdf3NY/rElXRE+SzMJwoQjVfHs4pLcQ9s
1Kb4FWVz2l+mbHtKWTBmTs/NseCpU3eWIhYCzldV7rpUaTuGVBEV0Q+w5Rd+BAi0OZCK6tmcCOZP
FzP4nN+ERbyyGjnTQZ4Du8pMiLr2Q1hMG9uaKb9aEjZ6vLlUI5AtP2pCTUZCvwCC63CsMa+mQJBj
d2LCbNSiZsqleJnIgv9jXhbCYobOvMUqDMzLMaQRg+NvG+4fq3UHY82qWaoUy3YWWHcRUTwUvD4R
Tcm1uikd5W5c6puZzrl38c+OKN+xMW44LDropruasnfZdPW/i//qdGU+2Yg5Vlm1wRppSuE5zduO
WNXQ7lymomO8p9Jv2yrR0Lsfc+lvKQ5Nrltm49s6CjmWols0Ky42UGQ5PPu0hfyVgnyxOjySVfoz
4keb+s7ILjxl+C1MqjE/YgviPvqgVqh0jW1hR7/CwM1umYRNiuGKjVOOQyCIGdqvJB4Z8K7ZITId
Av8v8vA7AxX/4J4up+GEVLrg8CWs77rHH5m60NjZkXx3o9T3HpMY4DjxI/EROg8251Ht/kyuNOpP
3CWghox9r89gP8gU18ASdalolYIxkC2i3oD2NPXYFd0AleC/XX3IdtKMccMj3YBKJ/xcABhtLZA+
Abql/ccDShvfvE8yY/lXsnJ0xvb1JXhpMqm5uA7Z1i32G/mOIEebiCMZe/Dou42u5QCxLNMPCvUd
gF3xMtyHiyHWihOtvz1XLwBX4LtCDsHCNJ0CwN42NcKG35RyHqu540Tg84ObA+u1RDUte+pYwF4L
klK7HQCTWG5t7iOgHnX6rp24pabZVgweVTSbqrQgh5QmdC8/c7hTZ1Kxa5zDf1M1oY8wJ0xafTR0
lmyjHRPd1PotgnzgMi7+Brd3be91SvuyLZFYWU3kBSCFNNik5HxSYCbbG2i/A0oIR6Q/ZB8nU4Mu
xC0xV4IogJXd4zT3K0USg83EaftpfuBTSQVo5DwaC1jJsh9GOIrIvO/qt5XwmLyx2oB8ydygshAu
n6ytjeM13u0WUjnT7w/vdAz6yHnUOl/Nx6+gAnBBnXcymGjpqIxxV3CtjUYeMDXtDc2CzJW2uEDu
inOSzviCgQb7bDzdo89hjBxiI8V/6EN5+04Vz4Y0wDWfxmQLV5S2EY4OOSxHYVbkwRvrB3ZGe0DJ
0KZGJYZuLDUmhJHfZe4Kuh+HVoSzIt32NxlfqTD4geVR22XQTMA0qByIndXD685oFFN4REOKB0ZJ
A5kEsAjdadm4qFBSI/GB0lJUSvxMIp2riCWnIYtgZH0wLn2Q8QRe2dNZGV9IIKZrvBVzYNzzjO2k
0e5yZV9/ZqeC8zFi+WeBT/pLnqQOYveHjrJObEk8n/LOLsd7o8CooaFNXWj7DDoicai8A8GzOAao
BKMwLqlvGScBmtQETIWZdqkuxlXs/bNZiNxWEybYDSVbj6QU5wPP0l0xresXT7zbSoo/5wlxBEu9
utMkz30cpCyEXtUJDV1fFWjAA8bd8fkVaW44sUC1SifG8BL4mtR2ayWV6DOvG6rUj339c/nokoo/
0vF6rzYDX0kBASXcGPRbTaEFzrN7fSuiVOM+3VgQRcFsliR4dnhDEndezf8UJ1WCc3PxqcSV0/j5
r7+oBKx7hnWQqfzKLr+JwLqKCEMCQm9RUI6t008E/kkYzz3TPAAz2MLzLnMcCzZnuANPx73G5opn
/CvB5RMTnl6/SiSo8G0FzMTkZKlZjn7ZwJV73KqmBLigFpoVo+olXE71XFA6+RZwBftf53HEB6Vh
OUCVTXNZk+qxs7YnbriyzveQNW28Dv/e5EtsTP1eDtJur0408nlrLIAu6goyhk7ymlHOz07QS5b/
pzdZ+B9Y62YZDrk+vWM+ab5pSnGru7LSdynrZm0Vg/EETiAN3WouSHourNZWEj+QjZLuyDcS48SY
ZKR5pv5DyzG5g8GxONvZwwqSqOFo55JGmkJZQkRZjIC8BgtcaQE76zlc+JBYM2WITyophWsEG+Gu
8tQzGBuLvgVHTwYXA2KMQV8YXoqp7eXcUXgcdaI9siqlYHdTI7V/FapmwSpTOx0HGfg4UbyTVKhA
Lf9Xrt68zQ9H0JGx61yibZDFATCM0dyqludwUQ9pZ0SD0CFus8nJs6RVPLeaPyKpDDmpdk+gW3Zm
U0oR4KEN1zeaXB6d/yib/RVihzR09og7gvgRGDhyNEIEv2IP/sEHwxwqvmGwIHj1voCk7tIdpY1b
PVZYl/rP4zUVicZI6RWFo1nF4jTAYxm5NerM35DBW/Le3XOvYCpX26t/kOKzrmZYzKqFF8ewdaKo
gpLVTFrO1pOxwIus8JAX5XCF02tfa3exDgleseT9XJ7zU/2j5wz3yWDQP/yH7I28W+9w9Bv29OuN
D2FuI5QtXANtbvvaqF+4wX8X/ncN0Z3jstViYU8KsTPMsdbfn458SLzoqx/yIia5YqJOv0alOFJu
U5l6KB3nto4sNZetCOSG+aMjQMXkUzp/oxE/GWSXe6bH58Cl6TiTpkPOCxT5696Sw2pavIcpZJbh
VVza2PH4ImOf03jC0LtszJ/Jsj0iCJp8+6HnUSGI29FWoFqqExKI0hvW2bQnzGdECaW5ckOH1dRs
u9p2kisl3MK6yBmGR2R6Ik9ccOoTnYQBivvimyGfwLCK8DuRCgNMjDsxSgZEG+SyMKrZQ9tjYphj
sZKY1hOS3wMWZvNnJx8TGcGi39Ki1eYz3AvocVbTPdyKjgPnkazIzEBNcJdUoOGioxXtJjlGjwE6
oeWorBssJjTfcNNKmosLrYTmBLCaAgL7Hb4aFSBtIXevJLV7bWSs1s7H1/xYhTxeuXZ536I6YRjS
xEzQAILJCh4MivvjAJVmpL5Y6zxL8e+karPHcEyBaaSPDpOxBte46QIa5vL73uy+Onl+8MU+EPLJ
+bGLWnKomwBYfS5OuOKlqyYtue7OyFXrOphBCjfwm3POoBk72EPSroK5BIJLdNvXmM12BpHOm7Ri
6nGPD2sqv0ArmIRFiE30YC50BN5k/0he/ZGoR2nuHO/yRD3O1Qpqr/Sa8nPNaWwqvkTQ6sBTdgTz
c1gg8xVJ5OJKXypKCAqEwfPp3/my4Ac8FZvE6GNcUVqANmpLGShMkZl4z+FsGrGhSm5Z0TfuHZe/
g1XHGW/hV8k8AD8RI2ywrjqTV1odKZkfF3PKBvAvbLXM5ltDXLnpVBAk8WEe2EHXGDk3RVJnt/aY
QP9nj4tkgQk9BSYTDz4USF4iq9ahBIZe7soeGLDvOf9ejM+GpR3OQA2Iezmuf7L7r2THIQkjquPO
cjBMwyLmqe4pxdh0/9TUP5GaEiueOQjCzer+rnwVQ3IFupNEDB72OfIyvP6oTqnJTfqulsFX3xIq
284GKnN745j+GAdO1GIAYmkJkaEMoOqkO6sjM/bGXfhC7F8ozrvkSy96zEyfp8lOpcl//mpaJf1b
hW/M5NKnde131oT3HDRhYLv/XxlzzvzYu7ww3Ntopj1GGkUnWYwWSs/WEEtsPbAlR4ceBdqIT5NS
/PvosKzEdakcjYUt1buSIfqsvaObPioMTk068hmqHpRCkx4G9cscG2AWTFGpT1ygdxdaqOgSNGSn
RhOykVpIe/3QlpyNIPByKr0Y3nBnwiqZ4975GssFnrEwEqlBHSURnbBCdx5XsEetKa57uetJVXku
FptGqUjZ6SCcLdlEPHSUFuwPYcT13aAeE3Abrd5UvFeD///H3pIEU5QXl21/+f2CprWsiXwXIPKd
YVm/7v9VRZH6Ab48wtxCVRn9Zg0h2SwVhnoeZojniseDfZDrwHb9unSWt8ULqsAjkOlOKo9MrXA2
50TvyvRoCx5NjRrxKUTvRfQMdXnIzc6L7VF9RPbAud5CESdsPoMY3Ew0tYAZVBtz7lhjA3C2ZXlV
JNVWM53Kz6lrKveP/ve7kOZv0nyM9P9wLYke6+yRmcXJ44bH/6eo+qqv0O51KnZmHbiYnv851Y/1
FzZz8ozCHFLLNDFYJiinUwvu2P1aCPglBlhXFf5HyfPLUOG+iwm+nLxJEayYG10Lf1QnyovBAIjb
PFuCxmmRiBAu5Q+tn3u4QUr7iUCtMlB6J7eAcWjwiC3l8odlrErDgdXt0NPyT9o59lCh5Be8ZCgy
q1nwN23Ycqvz0v+53LMDBfTvt9UKZZrL+9uqs7qZCT6TF3IWKfCU7E2b2UUm54X3g4vWaeJvMSXy
KgtwPYhw9DWSTqSqjj/sCtmn0OSWMrXfDCxf/FkKfAOitPwUSMgHcTjrFwYYnlvSCN5e8VJzZgBf
6bQ49KSRynpw6NESrf6LF7CLozF28IQdcPzBJfyttT2g+SrbH2xcy2lKadmAZlQyon+9vtgvwu89
0hQkUj8Tc/bng2yFE7KfnY0wjzjZSJCautB91SPAubpjsmWXDAS0HOeDhnKgB0UKE+Xd2Ir1rA/8
Pl9S760bHdPBrlC46zE024vftzXxz9QujzxmQsqz/+6XR8OT1M3snOCd3bymD4Fu7Gx2xT8lngng
gxJNT4q1JVZT9kqEP6Vd5RULBkgqZKVR2qEarTFCXQF2sKBata3ZGGzG5c7df8gtMGUvl6Ew9SWV
XWZQUxXI7c6GjPgXvMaRzAczsp3REE4poSnTeplM1WJ3AnU9xSn+tdPM6FEibKO3/kFTTXhNKAOn
oo7NhCxk80A2rcbQXXjH/VQXi041fXK1pepLamZJK8CVnII/P6BUclv6mTEdHcJu9Uqag1BQYbMY
wE8oGMP+ooEdtPJmAN+zxK8hy1za/Hf6RvLmt44mm2Bcu7XyzaBs9RyjVQQo/H7BSMVOy6WK0Ijv
qnxl0rMMVMpN7r47gDPL5K8Qs2Vs+gkkfCOhhekO4PGcb3SBF7NROJklxfnwCWrYl3VbvGMB4EnW
kQ45bjVJlXnryjeuFZr1319SKFWt06jYQMI4zJFgwG7D0/D/wB2vOHxwgpG+ZSsEHz69dIWCXdPc
g0lgN5/ZEjd+F6UqHjyqzI+qzEvLrqTDd+wbUy+b20jnk4FRv1J4neOSrlbFX8wYvcQC1XtWILIV
aejFHtz8Ax6We1MbrzkqCCPqpcHXjFCdke5xnToF2ZbjRazTcg65DG14f14JR2FvMfEwtUdHM4zV
DOfh6KAZqU/Ess3Ss6djgz5MmRQTaSWdMu1dMuPICVf1gayWOKAd1/uAhgNvPGyeufx8AB0KcMdw
hdDW4w0K0kTb1k2JnhZXjOlCLsupEPlDrBzL0zZfLyspyfgzp+Q1TMSjCxzj1QMGIbLZH3mMZ3rn
/n1x2B3JSmVtMXBUiiCrc4oIKyf2ziW5lDq+hLqS7po41iDg5FWMPed1LwQbExmBcUkJG6rT7AOM
zYP9Tj1fEZLUqOkxlDuiTnKFPBsx/yRoKjpYVSEwbljYQSa7AgSMdYqUUBvMYwxCb7Ehbv/sUr/H
08emb4AlLZPFmDWhyDd8ETqdGrvI+T5hmHjFC02GFyLly7GIB53Xhu4d0zoFIzYLeBB4kIlvDxB4
biLiXN5KoIdT0Yh9BAKSRwuai6nu7Dw2MsWu98UDVKu3aN28Uzcmxe6wr0D6074NduaJPJqKtR0o
30rxqeBGjFz3ZV6iQAh+i37Vo2FJz+okEkyQsFBjixRIfwZQIo7TIfaoV9yBFdA5Ta6erTokXpye
8GiuELZ+1Y4HzFdL/QDYbCBk0yHE1wSAzq7aif8j30IWGFFtUGSBpLIbV1tSZ+vAJ0hQ1uAbCsRt
Jn035jZ4xTDrXdXPXJEmY5qYRdnZgwilkBlMdohrDy7qOx1NPUuhlf78Kh0Zpfx8MwwkUegWXCRj
iLhP1fGF43qDqSaUZ7Z5DL9oGkIiZTXtbhtrwj6ZmvLTXeoPyoMd+FiEHlqfBkSy+TnSHiIRId2Z
nwVJ0fkv5W7Ip8fkyYsF5utEXdJGWduYxv/6XN/nXOA90KkB/hZcIRNYH1SDEfdtiI+owB9N02Pa
L0fm2TJicTxFmF3zA/fhAG70HadPWmCYFe/vXrspdtxue7tkZzfT5dMLKZTYnOTaAHJokgSLBuGl
IjIytuhP9GSkX/BEueOKa4RLZZVs1uyzFOQyBj4KI/RR+NpZu3CfJwitAJ+X4K8wvY/hnF3lJuBm
Vn8AIt7see+9ScGUuNDNnVAN0wTi3BTY/wbcvZCbSoGd28EAoUiQz2XYo9Zjb1ut6XkxXQX0Xof9
+LeKYEoR2578Zws4ypBtYaOp4sCDOCOfRk3Ad9DMRjdAX+iwSS+kwxI979todA7NfNIa4No9/UOz
6dq8L9Yx6+a7ORu5FY3TQUnq1AzvZFEPf+4vEaB9WHO7sXbQiqxhWq7QTBARym+Is7JAxmHQ/tm3
QQd3yWo80UKkd6nCDpCIqScGpWEcnCvddCVLcjrw7wuB5QfpRUeKzNhaeebVmFYCT2V1B3w55hYW
/XFKbNWJfRls1/WAJLq96Ot0/LQ/0jpfBY6/WF5x9TfbsW4CSP//Hf9CO6yQzhWwNo+ePOQQYbhs
28r4Kwy2eqmtzXaxsePbvv5cOd7ZVJc8UoIxdNN9auovyGPCBBXCxDl/08H+3wcVcnjkcvqXFS1i
EypXHPnsguiAsx9HtpfTw0H/KBuDeSAoT65hlXdaRUL80lk3nFx8C/ttj0+C9zTHnoCa08WqNFFF
RO7ZtEwKHXeF+fJDabHvupKoVD0PKn4FMdsAIS0UApX6ig6n3umzL+GlTUZfQIxjl22CRlpCtiq8
pV32ty1/08h3NyeGET6EG4AP8cegM+qpov2CoquUdLS47GRAxmk+1BK+Z5/VZs8ad5KUhd/cIOE2
kxwHSPTNv2vnqzUOQ0JneNNQy1G3UHD+oaKo7W+ZsWSiajT6rpQg2HI/Aw6owpJ7hRfl48d5XwcS
w8je7ip6dWFDQpmKuic+6XIlzQMla0Agogi6wVn15HEiNVzYNkzZcbQq/I95ISDHKCrZWp1vOuup
KwBHSMLEnMd+rxYp3/KJHTYkyzyODO6dqOxMHsY7IydQbhV02jCfnjeFu2Yn/MZDmnZM7njsLG+t
jCDr+sJd0EBRU/uGumuR8BaCFZjk8IYxxi5HJqB7h+2G6q23cMMSc5IcK28IX15Pzcf2QeZ/7GsS
6/SoR2AxOVGB5+dMi3lumn4spUXba3F92o4j9n3fRX03NI66/rZAGppTLG1F8VsaJjGhsbx+vZi5
2AJx3mbcDMCUoKlV6HHrPXrI9ZcVFFBboYeUYcA+7hVO7N238Y34X1c9D6FJwd9fra1EAEM4GNh7
Q18A2rdgQB5cWRdDcY30FOmFZgykmNRmt+Is51ShB6b8myX9aJYQvYszzmTWNMaEYyit6baU40KJ
tYxZdGqr7oGqcyyDp2fxAZO1b36vXYYNiR1asrsjVxK0aVRK5ZmWy+2ygEnYWN829HsFvF6DackX
xQrNjkIydsu+zg85YR+ewR8Y2torxjE+QJJJ6h7a2CflR46uHdqtWEv3tyziqkd4zkBuCjIhVUW3
c2tl8H05r1RMuL8WUoW+rel/TPqzj86cj9mmKrKGNig0q2aa8fYNSFT8lzWXa2AZh5XA8eupLIST
eBXTm1HWM13UdkvxrbDjJNVAQ1Utbc/dHMeqIeNGQY7VXzPTkgYjK6iJKLTmhLbt4RGcnBSeVUI/
QLb5kZREgGjI7frIqpUZZWsCBNCenj7ClO5lhuxug9mfzH4XC3PT0l48Zw3PZGIoT049dqTsSTqP
MnqYKG0RrTdOU8pLwjrcwWn4p4U5WXYnfRqg2en2mHj3KHwZTm6RpWQyu7vYh0b92sgHhsI/UVZ4
VsWqHVAqhAHUq9sfnhOz2hj9qVsKfZsNKgIFH2q8u4jesIaMJe55cU6G01KE6f78X/bPQD7HXYD8
PsUiw3Ud0E9yEQu1mHDj9UdQZWxatsXMWi7//bjzTKtaO7LFaBMYpK32UuTHYl5PgW45R6vR1/Vb
i2U3qICWfkjgI8pn0EjJB7vobVoN+0Y5mPeX0IoZfaU1Hx6bnDgTth/puf6JX/YDpQWHnOnqKdeT
X1Mx5AsNDQbg19+4oyAC6TjHPdamV0Ok5UXfazDWg0oWrQNCld0j9pvf3+DP8WPOb5whuQXuT9gR
5Im35Cwrqqrc/i6Z8izAQkNVepvGLs8xsQZucd3yPI319jU2LTp0x4//C9Oqp2H8HYPaboa6bz4p
0fKxIec6qbC18bHPWkpnqxebe9NkihT09IQs0mBJF5GJ4i5mtm9WwReRjZCYQgRM9MbTAAeZCZK5
AFHctgw+joWSMX8ngHBxp7pAyRMeO0GyRngA0Ow3jmf2unbL/aAigqRz8aHaPG9GEsaHuemuS72o
QwcHMQ4SX18nsVhgFMd21CrXgA3d+pYA7yX7r8o5OAB1y+Bvn9ZecADV681m2tiLARM12r1pZhom
TCO04SoUVGyS1Fl7UlQemIBSafdRyhRoY9MBY9879MRm4ubNMelOsHQ+LP2/wFOvU6g1rsaa1DwS
GkGKJFdRJtZUjESzRgqRR/KDepESxKLMrfXQnDlpOeN9HIuhvdAx6jFkyTfY3bJrP+w4MuT4KdzJ
fpolbmRQnT+uzNGNjNoTsvrvEeexxG8BagBVTGAIq4pFz5C5DF3MD5KoL3aDWuBg4OiDbuXRVqi1
YmaivFiD6852kxDGC+WCi8F+vdNL+FKIwqpR3Y4Kfpo4l8+cZpJZW7l0WymISLGqM9m8I/xpFBp1
6KgKAlBN3SFeQQPYNx5t5jIxySBqoUsicEMh8R3gm+ZVOVm6THeKHmOGftcjPgx5P2PvuwoNz4rx
WBbhOSR3LS1qfwPm2LFpB4uqMgsOKwgYgVhETAJmkwOTAmQqFYRYqSAyglLsm+CApgwPSDAkc86D
oFfJn3E30K6SbBWSau37KWCTR79EOcUGeDgJYl3Z4H+Kk02PuDbZb1Xs372TEpdW4AIu5eQu+SGp
1nbePmOH4FQdEX0hLIEO+X3UkVg+3u6Kx2opbtUHcDkv/2r3QK4oRpxZzmIQTtCbI6OT2y80reWw
qNYAghylWMiZvgSP5dojHTltW2VVoZ3ZHmrD+s8ogMFQkJ1Wg41JWq2ZcGrVfvA828DO9AUSdqux
5T3uTNKe54DeGbdhVesSj5Tbowv02A35v6ckwpGAAMVYbO+sbdOkgOw7AIsAZJPmjTqpEKsi4H99
UAnN0g4EYh4MVXBpkO6XcKEiwYWlT+iuC7hBuZJR+TU6EdaqNDfYOSfkWetEirA9VXNZXosawD1w
uop0JBjwseJ6Qqmkkcx8s/rKDSu/CdTopfQKRxo4IslRCsYjWKREMD26HwV/Ux5umsK8Ft+t8HUK
q56ukkfz5TrCfo1siTcUyAly3jRsZq4nhh2L9U3tZk2LF96PtYdJRWAANXex5keqU9+DQnwYwgis
8KrsH8fbAHUMOkeM3fCOk+LMIAHc4wDTjqjD+wj1cEKPipd+wymNtsSYMd35T2WqcXkWQDY6lb0Q
mXCIdCnrCgmro/wk+GRmAzBIpHq/ff2FM/ckr2fgX15tQcDrlMpVTHj5h2pBgSAqUJLsMtYxN9fU
MjtOuidOU+TsTZABeCNTpLuG9EAcNTDu1FubiPDk1qf8NTkgW70n1zxy6aVDsoU856f77/sZe7Xm
AaziLAu/aHsOMYdiOV9HcU/9BoFFqzeL1J11NqiIszJ8Am1brit6ep18jlFJkd8zQEpnCIhfPNXc
C7RqfaaGItG3SsRYrUJdrboTiqZgu5qxmVqa2ZXhcbdVT61ZTX25F6PIzfoW3uyR+G+daoFlxAEn
Z0oqnRht7YBoB4nErykaMraF/hyx+XDQR9s0rMxtNl6hCQPzxUo+8PZA2eeW5cfR8h+p9MyCYeCc
sDzoAokWSCaJfzMgG8bEQLJ5OsJl42gxAtLqb3XFPZBZ267jhQ7Kj2/8wz55nw0vX0EsczCzt0Jd
6I4GFTJoC63s2ab/l95CEZwgBDTO14UeE78pE0ljk4I1aOZdfzJlGsoCHaB96XemNHBxlJVldKgu
7LSQzW8juD34iT9KIxqMaX9R1aU9LYTp5SXZ4d9LFvBX1WQ4rDIzNroHSf1lWiSCAFOi6qFek+G1
j1zRdXlzMKoOVQZ3S9FClOHhf9JBM+C/ZBH7Ni6529LAheTHxFLseYZUYanWFSndGBjYtyC3fjQ8
N+E0ojsTYxey16t3afB2UoNQFH4sNY4wURBrJr2tiOfkrhwdUJqPZCQczI9Mj1qOVssECptc8MOu
K2bVrmRgvXsRTXd3QlDCzOrizjRdebGalgyKCZHHya5l+Q/IAyn3w3C6lxsDfFvfxVTc5M23GjQ3
oZqaFysqAM28Sosl3VGiIaSlnXwvXM2yhpgMwe9ZHZ1j9uxVdtMa95b6mmq6nOajJuc3uuiDIoq7
7i2flL8eh9XVlsxQVlvngH3trZup9mi1ZCd/a0jjYslq8jYnkCDsG2ozwhWGxz9QKd6AdLsKvwOd
EnwKnogljFt4JwMLYRUxiWQI04s52M30TUZr8e5DS1j1bFbMkmySZP5DtA6ldF5ehbu2T9dT5YhP
r0XW6WoVFv/TRVX+86OGD+JdiVtzQXwrv4CtUZB19v8ovQyzAlRaU9hkdsn9goYR2heodZW7sPPF
Ae2taWw+fTgrYhVisWVfPmwNQQ7D2nSEQQWIYuBubqGwNliUQpT9TKaKRrhUG2tuTJaxe/CpVpfQ
Mzjhf0j/8+piuFcfNscb/EX+kqPlYgwh8S8bxzvPMa4fyC36jICsfbjtWTMET8eJYGS2vh6RiklH
jVVSwChqmv4ve77VekWi3wcwhYFyZrbshN8RO1WZEJXuGElOszFl/RLqfHK7656x/KxRHYy0Wz6I
KcH3xF5BynnNFu/KZ7cYsC6pT5BcDbO1yKvOamPw18fCjdqzEVnFPp0ahWeDILYeda+oUzZDzJ3y
8qZ6SW7x8Cp9uCl63IHCDe5a1MokFGldOVAczzwWJiZe8QkMjKrWa4dURZhF3vk+jvaZWSXbYT/D
kvYnF0ChJs7uxxrAUjmFl/QPHUrSna+90eB/gEgdDOJJ3VGJwjG7mI+SPMCLjNVOVPryHqxV+ZPz
zFlud6TBnQl5BWLOEI2YsC0it/fNfWsUd41zqM7+8nKk/bHYRBmzdTKd4J4Z0fNaG9d9lLQrIsJV
6WbOwI92Wt4BHpdjweHBAQTqTNEnmv6JpgnZwzl6eS6uLAQKQYWR0XNerkECNNbZBdZeVZ+NdO3V
/LkYkAsoZA46utj6+0ndfvoN/DwIioz0hFZXIiaZiJqcZOjtz7gV603FoDt1HFzzfzpyHmfK8pKQ
1pSB1OA9IUgBfIeEEVifyQSi90+RWPXqAmCfUDuqWLE3MYm65jzKxL3H0BB/A+hiWRtj96DfEAsN
OIMK41ZtZONSuNz2NAhTys4b9QSgMBmS7lzIFV3XhE68C+FQ+dhAQANRV4e95n/myaZdWsxop7P8
CigzqjUK9QVTlpqr/xudXCwQ+CatwB4QdBQn6OzGhRFgKRU9IEu9v+1im1lFjudwKkOHRGe/bg7M
tvwyb0nGvmS4Ijd6wCRiPOQ/epyQegfba1nf/R+XIwNrRsBwFXgBewj8BGQ06EivxC3kri3OiQoo
2Yxyu27EmujajroCZ7zDerncp1L43bYIVP7pKiAhMSm6jBLrpmEz4qqD4O54aECys/bKtVr+GsH6
ot8GIaGwLvepUlyEBquRahyppDfApj34hhXo7FIWCYn7c82EIUrrNWl4AOYaR4uBXNoG8QVsVGcv
wbgrevXV0cNRVg1gRJrydEm4kO09ZHrzHSCTNhFYHX4/Rs7/3Fx2oFPCMxmEGRkmdgtWkk1zdQ6L
vw59/oJpJSnHqfC+gcM0KzT7qWpuHLbUkBsVmYDXnZ0FLA0tiFxg0gt7PrIIQ7QkGib6RyhF/8Z8
6zpyQB7hlcGkkBDafZDjFqvQR+KgbmCVGZxBEaJAcoKeqivMe5fF+vNKNWDivJtwt4esS1yLFcLp
spbH92VR036QMVeL4J6CZzDArfcg60hiCdxyfaHXf7pGhdozf7QYZC1kqjczx7QLDTFL5kwFTJzB
XTNQhcKnjFN4YrJrkKRgsxCFNEQcqAoqBZlOqjHypLe4dIpqtp2JEqQzylKtT8wIRinARNMS7Thp
DJGjobHyIi+LR0c+eDuERNStHr/qS9vCmka5FrYxcL5t1z5o+ipzrr6JtMN/eFpPyXWdFf2L1+70
AOFoMhjQvVcLT1NdDcFJOighsY2sgS0Y6GLrn1cgBAcddPI3eoBiH2glXJumEg7yjqsIPEp4txX5
XZd3udxfUv8G+MgBZ2subjwK0dHkQ7kSS8hvdx1jktx/lETb8sIn8ZW7tVYsQbmQdXIIpFne4xV/
SWnzfFHJ2qEa6PuL8jlfZQ78PsURDISe6WwNWuh7e0//uGuSNQk2zChOqpTP/Wrtl0LKG3hb5DSr
7I4QjZFvvUVUWjsqxLF7gnTzRanlGnNLvbmjjHTaul1dHM5DfzgXrccW7WjZJ/OkVR0avFZESWTl
MHWo+QR/K6+9Hs/PFm2QHarEjeRcC/Tq5Fhw+IBHFMiFms6d5cc5v6FqGM9c/z0iXwcOolNezjtY
dkmYQgetUbXmZeo/SqKip7MX+FSNymzTHjJpkxEjoT+XHJflrUMsPrSNssEbLcz6eCC9Zugv16ET
Yz9lbxKN5NFw5NX3M58iyav6gu12iEUv7l8vjjCM7NwLvHUQsM1J+vwg7WSgTSbxdJsLIXXVHCVs
U/ORgDFIz5wri0ixqi9unEX0y+xmM67w+zQ4M5ippQ4/J4fNJwM3r7TJPIuLG0rW7zIxhC1iniGA
UAsGfhO/3c+ZKQp21jDR5syGg+AwfTC8J9o0W4OSRoCWMK4tM8CDRE6aSIF8Ua+ZbVRj1EBBgZam
8a6TDcF/o80Pu2PuOIBcv+pa1SVJAO3fjWcrjaB77a4c+bqYBYfCN0pIPMQWtisSU4oeejWWr3mM
zzEfFWAAQO3PgAntYYQ4diMCSNMZeoU1bYM7VhLoTOhwSGgJgTptSeZBhIa+8kY13zJ1w87RHfov
5ko9iU8e8hRkLiAJJmbFDAWAt42bU5B7QqTWzDqZC57VP6x3/N7gwp7pu2e8Ljb6b5Qeuth4EqiG
a6/JD+EhNNo22qr67dpZodbQrh+8PH4ct/u0IytVDiiFWoD62xXJJoFiXKXXGkNQQ85OBZMHMe69
tBo1VRjucIj9uPRdNIT3emaepZbQgtYVPGBYUtD3VvBtIehxTEw6XNMJbW2VxzNmOePJXKKCepVo
WfVsVqt0EZK8wfXZdbW4zfwiF0gpDiKw8ravE0JHZ5/KO+K86sk6vKgP1NFDJ3PcLl2tce/DaLT+
owkwueXQxzqjxCWnSOXzGNiZddDARq2Cl4VdNjmPNXKjtBoYeVmo76nKvWca4iK/HHjK0gKlZdi9
AQGUhYydSXg7RhdAkNM6OOMxgXefdnBZejHue815kln3ArNr31WbHmJ5dcpDereWtAYUDLLbDQPH
Jn5AlBrhZ2pRWKFgQK4leJVNAuw5iG83qWZH3+xPfu+a3QQ7QWHPaVRQG7GpnA6pmbNMCYZRDJtz
R00CdZBu4apq96YvhvyN/A459dP+qsUnUFTq15qUgVRmVtNvjHgJQoTqmMDK4Sm9D9RASmtRp8P8
xjOFMcQ+R64vvuOk9BTmegCA6idRUb90pMoibobWtD2C3sq/koVFB/oJX21yLTKeDjV8iOwdq1q9
v1Mx/cXMabAuLkmvKABIrVHPTymBZLE34UGoQ1Qj38fw+UikP/tBUKTTBnDYP3oBCvECoGDdzZed
pjB3c75tAQUW3NbPpZfMBoA1H5u+dpsxo7GXk/flH6LBnji4K4ucx79pHdOoh3h8/f+OG3ZC5n0U
6v/KgbDDAA/HA7rYFv/GEnHo233xXCORYKbHihHmBPIBPRxjmMXJ0jU8mFU1aqHy5Tc6ZJxgTsX2
JO1t9SnGXBnIQikQPySaP8PZ8WJ4XDJXAjQ0I7g+h5Xs1+bLCVfwUz0So2LZMlqnsdbx+93jh1e/
1tXmMqAjBmepU57KcMn2ZtDOtaeeeU94tvtpZqR9tOmHoFO4RSxzuCdMxdbyWLOvYf5OzG0G84fs
/whCWJzMdi2gJJFI1buotnhZzM9z+FlAt9tbfNJBghiqto23moKPCen1ZwoY8oGVZqvw9lzEsJSa
BFAMBDkE96UcOhD8Y2abBkWQCL9n97Z0dcB8kK65/AeZyH7coSRWCdVTo9nyQhZh0dTjInhuuHy5
bHemLZqFD1rCCYpA0FkCaAQRKt/H4DbAvyiDYzwsiNMSF8GG+A6jeHLl2BGPaJXAn7q0Is1UxMw4
jHJbDRId3JNEyNmGAW2zlRdDLiJGXGQoEdsRaJTJ9LBHjvmqJyCvqdBHFJPHtbK1oAmPAC7He4Kk
tUrtarH1dzZo63XbuT2AAq9bmkUrV5z1TXac1qUUFwiMXuuaSL+rZTLfiCgFdujhSFS4zMSOrsyI
J9s7JfYl/5+JSfaZAuV0KGcjrxtsD+Fx8hbhImmtitsAJcBKzkBP/6BoqiGHYuDuR5oqxglE9BCL
hmdaxWQAKcJl0BLMknR5Gxegf70arKkZzqwqDf9VfamwbVLaq8Vuodj1RzO0w1l1V7rN3dHljcsX
MVupghxAU4kTFqG7LMmloztrZCDJYULxEz0VRKE18pYVEYYWx6G61S9o6Q+OF8KkSigfGSi+YvY1
JZt4e6tLTJdDLlAXLuyDh3xLZ1hce3KWzk6dQGeppCo1ewz4ysXYB+VcdPBgDj8jxN7exkpio/EZ
MwCI3Blwdehymeazu2aK7cCNdT3ECfDCi4Mwod8NbDyOjXK9nWfI0BsI+AK0ggjnf8xrE8qKykL9
JxLANZS7xbhut2MN0/8uTqecAy5qYlaKdg0jPNE4JI5ttPGT4Q23MerKYuruJxw4idt7qOO3XVun
PiFenUh+DkDviiqqqPbSKlUQOtyV2Mk+d/2ddDCDUn5tWP28xH6H10m0P2LYFxtjU8xfRKJL8Pjc
yRNg254wJwLRYzBqCoAAK9h+O8rL7PYcsCPeZg28YCI0WvYpr9xIMKDKDdlux6dn2d7AdSFJ+MUE
7XpTnFXSM3aky5o3pfRiiGLXbmXC9/unTCI0MaZd/RqNM90wc67/UXqZ2YlHbhpuExshJfa8NtAL
KamEN5ygJkUXBGBz4G0LHxdqFqlDlOLzbHjdNYHg8I10l7RmuZIyReqGaNO0z6hsyMRUgb3WA1l5
s0KFuPIl21MGlTFkv7tJPtRqG/XqIWGyLUSYgwfl8QyrIbkRrcfJBbkJk0i0iP02ihVUqoAaFWZD
a0GoZGwVDIaeAICAjlLX76frSyNmpx/ogjbzeb67JTgItHWStMgpv4RML3qnkdz2pN0lSDBeZVXO
2ATtNdglCHiVGnON+r4n/7CR7MsYbjqdgQk6qEorLtFfflSWQLJKx7c9vMFR9toISk4NObGqVIkB
9uqjvKcKCaRlNHlTdoFPs5kuXwQgyAHyGwIk/M/N7kzF6nOraIWJ0DU+sesHK7Sa9lYIYa0ZwZrK
VXKkQnN1JuCToA8C+6ras4UE73k7vSAGO0/HFt3KLEN0umAzxIP92vuCgFNYOxXGyqShjmWquqM3
NeSyDegBaYDQGXuL8rmKKuuQkmxV2ODKGY29BxIgFF8KDEm13PDX3gqQUlcHMLb+H7ca4PM5ANAB
Z2bvM3Z2FDIxdn4aOp+P3eZxtdnhHEhM8e7eW/EvjTRzCee07obcQDaxzESPYIRwbXPITNpVit9W
UWy8FdB+sFwg7JnJ8ydlD90kScJ8F0B3CMCNDMVVt9N/sJ1OctDf0WriwcjDc9GOffr/mAQ1o9/+
1v+tPN41fHkiVIS9Q/8/ezKq4zu6Ya7tVQabic3YKJLKtlnqUO2iMlcB6lFZJYi8YIyzqArJx/+I
UuAQNQLdtea9GgP2sNHbRKqR9zod7Xi1Er9A+UBJu9ufjCsrm7lJdAGslrGPjVMPgYYOGp+ujIPq
guzVLfQZ459JfOJjXSUzmK7+sm9xAQBZgAjdVOVMIR0P/B4CPABJZkFrfNvylbJd+Zss1kRkzBG9
TVv2KQKtQqg/e0mCAaHffMzSqDNpuUsoip2lT+8Its7rO/oHkITs5WQyiDkqSTUp83nt+TDN55xg
UcqWP82FkKdQp6KW5SP/k7mid/bEnGkmwjKIk66wmEbTUyd5TbftUvNxEHZ6EaSTS7mnO17ZSUhA
vExmzLwEKT8mFiVdTwZTns/0AWh+1AnSCw/Xmf+CHtmruAugIQn2/rDXh5MTCbutMNDtZUGKYpN6
lQubEcCrKbega4ogcd99HYzsJ8E5DGd3i5/zTly6LPJ54WMniPo96wOssplgfoChiGR5cY1Gatna
y6NMim6fNlQtKsq1Ak77PKtQ0c3lYYRSirfSj4WukvskQIKhT8oSaUd4VBoMBTspSwVPRFBJLpB5
BFA98d8t229Ml5eM48fBD6cZQHZHF3eU8lAGUIt+PMrVoP6CrH/s2rHoEhdEy2uKHyFjoXRSCxt4
dDXzp3rHPQb2VlC1nk9IrcQCJC6zaqHN4LtPPaLJXxS2FvTL4KedNTFdEBnvimbaDXC6dgWrq+cu
7DI+qEN+RERAgFaH8NYmhe+pOnWHgB1tnADgrKWmTLt3ISuX8i5hgHuOOEOLUbEby6Rp98p7NJmM
+ICDBNsLwFGLG3lJr95V+XFlMAkEHIwKeIGyLLsnYPdBXE5GXcQA9+qOm7S2p801Nxvset++IzcI
zwUwreW+xSUNID2Nyon7yiXKagUSYrvGXEenlm0EDvhveQhi9rvBil00n+bxlxZdPxMMKsDAn1Er
gm72JIkOwLKdP8tJBibN6vTPej52bTSWGD5FGgnj6zba42zGFydGk8zjdcZnXUPbpite2MhjrUh8
/4zTsxMgGDyQDyOf2YQYcOcQ9oZQ9ug6HXHvvkIWOJzB2IuEaKA2te6oOu31rZUSmUbMmg0nitOp
bw0AiZmHEYiUUIZkO5tTElUQAlfhbqZGGjFlESfWg7fSvhSqP/yXMC4Xynrd0hBPGTIzVX+K1k4b
yP6bYBoVo6pSzTHfKuxdGjnOqaidiArSfZeRVuUNt9yrfRVffuYY/KBcqzyaJotTkOZTT4T3m6/m
Bk9kN/8ONOO8J/fyJ1bbaDTiDwB4mYYMEmJ7CIyP7jGvLmSMImuFefUTk1cS/zDn/75zpkigh+t7
qUGmNCvnoHD6KjYmNeikQwN6DAryZKGOa2Dk4YF/8rDJHlOH1lk0+7WsWFQ83UUjPptuxhCd50Mz
nMYlLtCTQwozeG8mjOngMO3SWnNBiRs1vieV5dCerregp5fAVNUSGliQF6b5xlOpDxyH8OzSEW5v
Ozkp4dxtqc4Uh7dLZA/lhS0kWliLEfS+qa/7E/A7MfoSoquXEnQivAYKPak8mDuiZRewbaRMpH92
NfN4h5V5WDKjQS1IF7/i+Ya0B32vc7iBeWi21dEMplli1+e9xj07zBtC7DvU7oef9L3iKwNdyURl
AOtG57SgyNL5WwptWaEjY4B9YZJTyOvBgEVf7OjOZLc/Dz64li1Uy6E5SwryaDqgc17aptzzPxyR
3FE+XamrIBR71N6hUhaf78LeUmJhXC1ux6pnkkfi+oMvgzXxH/6Tm0TH8r4PLOLZL/xlfBxdtAb7
7uEB1SvxBG7uvcwRF0jz+67Urh95pi0E8Cw5xiQ0Fxq8SCcCctmrnKnPLZKlSLMec4gLg5yCaQzR
dApgtcW/fiAzaDqpdiAVaTiJk1KL2eGeIoK2cgAmHtF2x6RjckDM2YKnHi+k0qEXzb8WJ5Pv/W1B
l2xfJN9X8is0NIaJOnMXCSRkO9lVyiawdZ2A/wk683isfmK4ySc9T/8z3XYayARWDCv9zsFcgvui
sszsRDZlJblEOqncRlf3B+Q03h4hH9ikYf6RFpgRaJlAxOKjhsGHOUB23h1jxQXTAXu+kbdJnlKS
iIsJ2kDvk+i+UCIIu5ZL5tGngmt7gKfHb2Typr8P1toziGUWRz5usBw3t8GV4jP7B1Uux/wHN76k
+DRI6KigJixi2vlMzxemkozPpnfKaulDgaB+Iyy6qA68Uqo6TYEnW+46+wISEWx6G2P1f3UjjADr
Om3QcrG9nrzoThYMnBB0ozOYlESuj/8lLrtsOGGN7TlQHkeNbpY9gxJgqY9onMs1031/1Vw3mFSu
NeJgYWGaFaFu3r0fYLf26OfgJ7eioFy3SHNp6bpUi9DM7JppV32znf1heNSEzd3WNV4liG3rNB/t
NazJfoqed02JWqrKjrcssyUj+EPQCqUiNagSUT0mfUbxlhOcSnsjXJXSXXG7a4h1jCPRxH7WO8Kk
9K2FDi59CmMks45qadT1EjY9VArT/anuAKEQcY7JLLtmDZio0iTg03tNCbd4QgXNIPjzIkslC33e
vhrEtIJawqWFXjkx9M9nEDciqE3YpviJTrIyutaCeFe48gUjKIrNMepSLH1Pt9cAcjLAUCs6I45i
48kGQTMhPv5jxaXtgQcJoOjmPSevJcL5FA8WIr1jakLsvlKZFZi31ZtsdmERqiGTtBoCwlzfBopS
rx/Xl4PvUlD64YcwUYURBK08LmoovygJdbkIenLLbBqL0w/F7c8//LAe+X2xczKfV5JKDdHA/7/d
1jIyhkhmbbqHFrOB7uQgA7En32jaBzi45/cAzuADJLVAMjE7g1eijjiOiPIflFa2NDSS7oX+Dh3X
bp7N8OzvGgexCBnOPhyiPW/R8ZVIza6o+yeq7hNdAoCIB+n0rKwx862A5mtmq5w0qgIms4Y5eabE
HfnUXENJHvu+++TxSfTaFBJNaW0a3t11ljLCbBys4ioDZw1te0G1TWDSBVezC9y8GC/FeZgwqLY+
OkZyScVkD1w4l6UcbEMC2UxJf9vNT/81IXjUX4MeaJSk5EYn7soSSB0/kCooITJ2gNM993EQfpyp
BEUy6lEydz0nPfQ8fCD/zpPvMwAnrWVYy1e3H7O7UGlSssjW0bFWnLvEXJBeu+ELbk1Q7dsx2KKc
A6ojRYRhmGRFSacsGnAhN5sEfzgYAiKp9Y457/GZo5gEYmjQZgs/JQx/LaekS0JxaHDXhLXg78WB
2St0a8Y+NCig6M/YgAgjeNUdZ4vj2T0a2/ji2Eq2SoxPFnCZUK9NmyLRhUMX5BGUH3O1u3n1n2IM
+wGxG4RbWC0Vkx/YEiO7SC33pgomLz9Lgdlhj6syMDY/2L6eJbzu/O7MgPn623hKYUjTobACaonZ
W6IUGKaX2b0IkeuSoqQneZa54K+Nl/JaHuJAWyXSKI+RqrUla0/HwhjfH5gFMjZyJEostuDftov6
vfm6vEFRV1Q5dRpDmsWewT8HNdHJCK/4POAi/hkJZoSTxMdQ2Zlwc2mBqex3TDnJ4eJZXSMctMrI
uIHIbv7s4kf6yrZSvf7kV2w7leMu6+9vZJ+fKDt0DgdvQeLKoLnn8lCB4atg7p3AnC3i+9JyXGpJ
CO9Ck1aRiUoWFbxTEQbSeb+i8ySyhBvfL2rD9zwAon4q9okUn78VAWsEy4n9B/fYhF+Vlt/97chQ
IuYa0I4nWIwpnt67u81VkYE7kKbEP1kwY7d5SO/lh3+dJW5FbFrD0fae3ik8WcKnqHUI06gSfTJm
p6GayxgVr/Zo2LWh7vLrLmeLp78plIGE+BXIbf00gAyaxnI0X6S0mIdCVqO3lsNPGiSzCdyzTk+u
mteT6J94TalnByEOF+nHtAem2oP2KHo45XwyUB40phyfqVR52NmcRvwPI2rGm6kEoMOm6pa2CYZb
3zo9I3SmxSXIDygk3ct83Q0rL9DDfmOnrhpUeVOIrkTFXG3F91ImQFtKGc8FnJmMmR4cFbELmi+J
8IBL5e/OMfTkIPqi2M/L0dabChmXxP3Y8xrbV5YYaXSEvLdfCySl1Je8ofCjdsNdPYa48t+N28vL
J+eCpbshM7ttav9JONpCTcOcRG6/Y287U2i1uOssBEwmzZ3F+SG/EShY1I6OgaPuzagSzaV7LTEZ
CUF1g7h6wKXTd/dO9019SdFVDDUzxDGLNfuljwAf5pgBKosz4UJMPRFHnWv6I585qpB7qW2QcBHi
zDv5oS3pzl+iUvGlso70xSLasqCNZuTxQB2KF01YNuU9DDLZX5or9ixlvNrwtZXoueijmC4a2Kyn
gHf7PVZXeKaPujxmi3pjZq8a6wrgkPZp4nh2IuLo4t/oXfGe6j9LeZmM8NhqnbMyAWACDPttiYCu
2I8r5j3nYPBQdCpyPOq+AFpT7P+vhuEGc3qA0m1oeIb/EOyb44jatOTrKbLp/4nHf1EaF7LYxPq7
JGZkGXfGmVHWFAiEB6/EGvD0U1LsgEbqgWz0RVqvsQH8R1bz5ewA/sdE/HF30cstRN/sZikCONlm
rRzlfH2VS3GfBR2Q8XfpEic5Hb8rFqhBzgv/L7MtRoD1IsyswBu3Sbi8tE18q/pnlV1NXnB/dSSY
Jk3fUC7jw6cl+ITxag8869mL1bMQ4ObD1kHs3sMy6D+PKaTARa40NaGMmCrP3slzo/7mNE5AvjcJ
fk76cvgZinjagGl/47SYbKjDlQ2yKDMcndwIGo+eH2tPj5wteuQ8t6l664fFf3dYiEg1NRyPrIMa
PGYuf5dsJR8TsBjJQvL7ueG/Dow1Pe8zG1AxTSsIP0ksOOHtgFBwCqRL7tei38tyrBx3hr/gBGwP
t1IWHy4wYK8TWSha4nfYD4rSAexkKMG66eBc9pNJNDHzICIj+F7kgBmdpUkvcMITtSQFWJzMW2hg
P9gwPS6se8d/fe+uJpk5KZcAQsWaEXoGtp4HCjwt/eA7wejIEwNEWpApbeTEAxJBFfKFVccbL+ql
KcUbEztB1zJuhCJEA9I+0JVxnxnjWlLB4WEWKyePuDp6OTCJ+MegM/PW8SWjjS2bK771QiJE69k6
COmtd+m6E3whB4crCARXvPra5TxKR19GwYhTbCm0Lm3dFsJO8OefAqG8SmMTcXYqFhLAlxUdyBFr
TK+Nzm++hBDQFd5GLbXQUgQcAirG8kL0w/mJ4F+RKX9ehoOVrkdqv3xibJ/aIcpvoVm97P23HT4M
6rhc174yZBMZLxpIIQrWLFL81ZFbSuWFwN/thwaisjpNJ9d70UhZcNs+1Gp6feUSNJUyYtaM9L6b
3pG64gWriRK4xGQySU7JQ+UdKoAeBIooCs/tq1ATATqw6lDWIJydBApjvM8K+CVQjdJ88deA1t9i
m7aaAl7DlkYGy+1bECm2GzzrT6XSzFKEl7ljNBy5rMEIhFMqs25eP4pxIgKg1BtjqKlB5rPWAhGX
vtbku54S8tI05YMDb+hl7UD04C6HjyyMK+oMufzx6kytn+4lyoSwje+ig9V/RCKLd3t5ydUHBPG2
bRaYgQEZvgZNFdve8rXKVpOU5anLCPYKoCMxdMBkNPXhomdxGB76vQ8tKlDStF0An7nQmo+UszRJ
f0vpurjzJfUnGlqkN5SS8LhTWn5L50J1S6QlCvSWJ1BG2M6LhXs3W/vq1IFNOycugmePWnSPrZRJ
1fiTSFkZfMb9IcWcCOvRIFz6iXCrf+kv4AAlwNk4msCUZlhbTd1mRe9uXSiGQCfR0QWiHB/M+kVj
MJeGYTiKfy/ibHZGlt7MukSytZxNvGL2epuydlgBuGa25Oh6G2tFELLlm1wHtAN7eg6JPqyRd49z
I9kiKhdk7lxbSVWVlnuuqavQFgCcXfjQ4F3HgeT0OTQ1cENzyPCWUi5AyQiwcb/KS0Vk7c+RIn6P
QvYUCG0fDanvA5f/z1ggaCba6vyCIHno5n8SHjZZkcDZgSXK+7ZBxwAJ8ZrmAeQxv5J0wsP5ZYuu
aAqb9cnKpPO6YgFE5S9MEDb7bTu3ftDNrRNKg41eUgO1wFl4V31Zz+VVnPIzCJUB2WxdOkqWBhh0
sjXCQTOI4ah7fppxfSonUuVdigE8FrN7Wz3SUj3agsQHH+J3QWwSW03HeHuPE7Hi0d2plsS4NO4B
cobNZIJXQzCClzHTrwD7Q7nM99BCz+fn5tN82n2dlLMz5j76clXefL9ikwLKoKAJcxprAcldv99C
s8ZaKMdAxwpZrRdUE5ovyuF4j6CobJ3szmzeIZEWSUuvlKGZhU3jUVrb/4fAp3RILeyNUuxOkZBv
zTwGz/2GsTufzhDHIoXZhnDT3gc8GqcOHfzerHGoTYa7wDcQHnYVhe1n/U9Lq7ymZXRyxYASgpFs
QvxWCv0EEqrVUKNTY2i7uROUdtYMhWSdEki0freH5xffquqfut/ccSz/+xRckfWDXlMjdnFIWoew
fYothT9UoEgY35j5tZqRerGJx81J+5XXMgwOB1RbedO3HBXvab5Sb6gFN2gtvjKr+ikW/yICj0NK
JIYzIXTuQD2tQHQQgEWZQP0isMOpkUB9QXROe0FlwflXv5aiw32tDNpb0H2hj7qHKIGLX2/B9DWJ
1yr7v+r76pyyivQDzO4gMc5Zx0wZgNGIxSm0zZcOLQWnsIolY8jJO0zWiKcP8C4eE5banHne9OMk
5b4NkxQj+f/SFuFou4Cudi7IrXvYuEH4npk1P0bp+lbK59g84drCUyUaUUio28qyFj4s8hwjAyxb
IOF5LhGEgATPmr+588lMUja6nSOBzyCpwB7hQBAyNWSwlOpom2Jfp5Ozdx3IbnITY3YeWKrXJM/Q
61YNFLrFwti8hTuxJU0fpS+wfcGWyJelj/pqzV/oyTs1KceR43KXl9x6D28k+Mr5D2hdfeshVPDr
TKGTJdKdxajKPZQpGU4blQVlRrLD4CVat7aOmJ4syCVkHZhk5hcL0Fwf7NuAkjr+4hGbC7rH0lxW
uyGGFniHylRL72Z/CxPinapgtij72c+qyLgvLibbRGxiX7FB56P40pXTVsyIHJsaIyjLpSK2vgeH
MA4wlhf7SG8C254WE+e0lrP91cWz+3KEOAV5sGtL2N5w60uwiTs1w2cxcNygV+3tq3HVTOc5z7dB
qElG59wPoWwbfwbjgURPNlJJRIm+rXmA7gnxmkIALQKnjd34gECMQlpDdU6NSAuFgz+rJWvCPhe6
2X5QbKjjgeBqVeZCqNoszG1+xl4gSQ9K2pHtjDNWtpvE4f+WO0VrzP+ftI2XivF64y3a+Qg/U7lb
d7e1m9uaTzLTGPaQBpEYZpme8J2kGZgZDERO51g5HOv0CY4tqQE7M+aNdaTN+bpE1hOXJunyceMz
J7eBScO+UMPDD7kCrxQm5kQN8j6oU4MK4sKH525juLgqsXZUJs/Z+h6tc85XYY0pcHxUOb12XUGr
Cf0KpqG1jqUXmkEJtpdmuctnDqBuMI9EvG9aDw9ZnhnV93DJdou5wju/osf8JruZcSllRa6xH6Ke
QphzobJlcwjDMSjgFezRxNWcLVECuuUXW2zD7twflWUVv4QvUYBSzHIAsf1LxdD0CAJpD9rwmXzy
mZzJWeiM5dlD2RPW1egTGNb1iCzg9BKPTliiFuxaGs3+MW0wL3yAYXYBjwaUXq97odZybqFy5J6C
Jlm1JFdVDgQ1fbxWtU9A0OVNVIXUS62rqlttff7JVpy6wHeWxZiwKx7ddyDPwVVraBdQbmGdee2w
uUvu1YPb9OeGllsA6npbnMMh53x0lvQRxn7pKLPO4iv3dEb42iTMqvksP4EGtztJe6IVLW7Tukvv
GCt/37Mu2dIWCU4lspQNtHAzb7DyLEPS949qFSu8K/gVuijaoMSbHYyFsrj9yo5f8Vm8FHygqQMV
agWzkDtYQ9EK/XURuhi7qTHNjtNjL0W+thtus7FeeG8T4z9huT/e4zPaeTTpK3OQPYXeKamrniNH
t1U4snJKhoNzSIX0Xk/fE1X8FugBiuu4zZsEYe7r/KNcX04iJJx4oeSeL9C6GnVPftUL3vUgOd61
ChRgCxU7alV7sn3czocTO4r2a49c+9RDT+KLt1k9M1Xiet3ZKsw6M3fFpsz7jHGjR0l26gbxX5js
PN7w4hYtJtfxo8y0q3Hg0tq2xATkCEAyL+lr8vqErnGMaSvdMdS0AfDWaCbpDS3l6KMKKuu6uaqn
FiS8gHFlYOY07B4Gs0ljmrTH2zD1EMOcY0UyYnT52FYaiuIFHu7yJmNxW3xvIVtG4unl85s1fk/A
dciLC2gCTsAjrCBlDdElqU72zlSK3Yno2jDJlbhKxi/Hhr9WcKCIK7yGZNMsD//5vJDKK6EQll/b
QdXr3KpVs+TvBHTNanUWLKnFCgs3o2mYYYiVNB7gLZBn0t+MNeNxS9GrF5Y8qU5GqrK2yP0Ykwkg
UzAqeaUOIMKRZYKPUnrl6CXSCL7b+Gp0Kh96w7aUzka1i/jx5rxbyNbkiEqA7RwnLupojJSPtNBX
WWesWVStj1K1pb9+tXAUPQXk46G8Ub0tPOFIJw8AtT0UflwoPNZG8jLAO5H0qdK++2vKiJggsdlh
wut/xFh/XuITQQleFUDJhDw7gyQ1yFK2a2LSE16XSz9NuFPXtwV9NOtW0Tcy0OPw7YoVDXD9uz/Z
Zc++ynVhrDLyyB/uvFGYin4NVRCLI9bsHDgZGxhzNQAbu8LjvJb8yqKEn31kZiesYhZI2B5//T17
ZiyfDSrjZavFAs0JhpcFXWd3suxpZ0XRonwWajXKXoJTBR9S+dv02Jydw0X8kdk10KzNPPHH/NES
W9oC46GQ7waBoru1bZJ7vh/QMCedBdsDGQ4mAzBq+/Y0sICZQzdrEhc238zuzAoB/wldM1tX6P9Q
AA4aoVJalI54p7/4UMccZZyEwAK96wke62nmhnjVNPdSmAkoZon+pHrbVU4sB+Asfbnf1iXZhxON
Vwyg7pjXEPa83RGjrPkICA784secqLJepHem2PhhPAraJJggbWjcoWlVxfUXqD6UYs1iskuv5ZTm
U450LJhjlMJ4oy+b40i7vupkTu3D6ev/0+3SmUgpOAV8YAYU/9RZv9zYGfBx67GLpM8voyOAur5Z
Wu1KYYXLQYkJjZfm26DVVGim0vtsX7B0BwM9l/xrg3twJVAVYq2/qX3zwTdK8oKPvuS4uE+Yj7+s
hDzBP7SW5GSbAFdAUEQ2RBSZ78xrPkrh7vv/BIOMupjF7WwQbgKKgkOdAmeFYpofsY6Bbsx/8aen
my4EdNmc7O5AUGs5Zv7i1aggR8gbKGnkc8CPVXabl1NYQug4Q7kvzn6lMan1ktJIfPeiYFcDyFSn
+wIsvEfidRy4OCtjZwVfJ7jzGfZbnUAUYZYTIeaB8IyueCXLz/qWZxk3PW5GXZWLfnkfX9WLm2nd
tX9hR8trvWGv1i5Bf9G5lidNLdWPuus4G++XPNmMOJJGLahpNMbytT8QDjM4LwWoFuEKnMazxKUy
dzHcxKaBcWUAPP2JFmMbnLtbIK5RXp/l7OZQxRJomTBfBACTdbHJ1xTeZ6ESFgzjfME3S67HIpR6
ylwM9ykl+y+ub1yPIZx+AomcribMI5ijOq8WF/HuhX4SwHgbLUIVk1+lShKdnB+eZ2JtHWg/c48l
gu4MwQdTdSp57IhSHHTHGjsu4TZtLmV4TfjjTmo8TzkzWdy2zMH30kOpfLIG2/YhR4+u4p+vTXC2
O4TLd9g0uuBP2g4y6FwlxR3n/DeY2XIAAgTHJ2m1lVslB6ApHewpfr6yH4Y7qRckmU500K4GFZGd
KurMZc2kmCqsfRMQAxTWvARJnczkpM1g4rk6cnF9t/Hy/caN6xz7GAFuS+129koMwL+hUTEa73EI
XV/cXvaOZJMNxU2itW30lzXKonkcnZxC4t5a99/4sA6Yo+TFCcNPff5HAYwwICzzXUIVJLzfupnI
kLZyXDjoJjCgBwykx9ose2yK81GKtVpCLfAe6WZhw1fPX1ZOvUHmmGvGo3oLBWfpCQ5EZZz0yrr2
r5mRHqfJlbq2RWjRTh0WoQeBU10G67xdiL11+0xyAaY9qNPnKu9rrSW9Vz9Ip98ixks5F+exUZmP
4A9c86aF9z9e7b6rosI8MZxShzSKc+xZAeqn9Y7FRsq10XDinRjrAr8+PtmQe19H6SPaTV4NUwop
kL9C9yXlW/a6ZTLkdi/MHJcvmVPt2NjXBbeh/2+XK1aWsRRyohAFPwXXD3ilgWLL6BzkkQr8DR8h
kGk6ErZ5CARXxxrEfNdvwDFi8ISs6OdmXtOygvH0Mal9dPWKm8U+fyL5VZn+PwGuXhoH/muRR+J7
y/NKrTU7oEW1xSLgxhdILq0S2iJVFQ4KbscUZ+XQxWKktZsM38zYMQB7hpi8F1IFQu48SMVXGyH5
eZCdCnyOYRdI4O4+LrH4hWLfLiAnv4K7PeOhr5lH/vUUFxIB2ZFx4MjIlKRmx+qwcaDXON8e+QeV
l6/N1iRzRyUHq+d3fcAD6pGr+d58Tk+7CdVqeQ/Ks//PP5tIxyvcdp0aAkeWvePgiJ2N17q9z/K5
agx08jHJxslH4AVT03op23i6V32YYQCLd6JuPEB0O5cG9DfBmHIvaQuSeS77EYZbV5k/qpC8vTQq
vESmNE0cRwvLhlUa9OCOAS5xLHa+Jyq24AW1D5NIBNCDBoTK7GDut4oMWOCHzRQu+pSn0cGmBfB+
LBqGGarRIsK8CTdzF+7QMnTQCNsui7j2G2Z0AGm6aDjnHg/EicsrvL3UhmKCSH7m1Cxy4qP5uAV+
sv4hhD2s0BMavkH59pVrPZH1ODsLGRIr8ul3w7UuLu9U5ksANUuL54JrXXqhXPL5bOAa/7l11xmp
8j4DQ4HfIFz2Oqy3K7RrY26zsrR3IxLulsr4rECNATCrsXCm4LBzDHSX236l4QNn68LkG2eMUIU5
xENP0yyQDIpwrGShqL61z1/C2irgdUgLvrh9i9G1TMhZ5RDaBRHhlE0NJCCkDkj4gbo5xoO6sLTk
cyzwb5PCwm2rJChQyQJmtdC7mzEbgJZ/F3bgFSQgyKLbqqIQE1BASlxv3urab9bneJiA2WRKb4NJ
RancVdzIC9ewpSKO65DjC9eGyyQnORRMW0Cq+XecpHw15hwfiQDASyo6phUQn77trcXZ9NUd1hKD
MRtJhc2uP28SsB7aoSN6eivlHsrYEvLTcIG3beDunhUy0STbUrVOHPzIstlRb81voeexgbvturRZ
Y1KqsVBrwIbr5bhemPVIgO+o18cfogc3yvnCGCfvcHj+kUsuab6YxqepkblF9xxwx9L5a6FYKrwj
UakYNuPi5ypVnFVXyXQNQvRL+cVTXqDfv/+P3XQ/y8qU5+w0eCCPQ7s0bTO68EsbQwY/P7H0damG
yR9DuUGcZf2J7yK4f8mbKiPyq3WyjfbI26vio7tDVTY5aVhjOQnVnRyEexCzLdjqo5p+QpLtV2Gx
1VvwaWua+FkfHRlAy2ttPz3yjREdHXmOtAGDlpA1OL2Xk8sy6NHHzSXnfPwfXMvH19im/gpz/wMr
a2W2DZNYVqmYgZQX99uQGupe8wrxiDoDM72Y76Eszc64lvErMylRRcwRN0pvcH6j11Wu1MlspXYU
w+2GGVtqsW4ayXR96Z7EFNli7TdDRfFBRsdFlRc13rV58QFXs3t39IsKi8o3Y71O00lx5aLNbrwF
nqyffL7F4u028S+zPReWbdqLg40IVs8ES/whOX10EQCTh2IiCXYklqKWQLDZCwDO0o7DJAQP5z+r
JPoCg81VXi9M3GG6KnXfI39j2ddo3bAYVdKh9Qty8C32RzDZhYD++ZuE6Zp+vtM2e3yXMEWipIma
nsQNC6LLMQ/YtZLpkX0OZYoMvlp0ZjdOmfe0ozKOs+7pusjW/GBDw0eTQ4CD4o/rM5+Xmjrpkxxk
NBgRBZkvghH+dgXmgloGSwfXLpVGNrF81McJJy2p6O/sNdaY5kHDg8wuV3bVbo+zWuBDE6L+04Da
qfjz8mbbNvitLc0XH2CfJaIX39HF3EisHaOuKX91OC3W+sbpI+MSf0pdKO3VhlYQCj6sC352y4eJ
OHDZuUsGmVySMnVesPXKQyejaKlAK+glBZxm5b9LsQQKcGe8mgCjsj3TzWpUzUBYnERW+F0rszK6
DuSvAkU4bnpZceLOnRoi5k4GWUo/Z4qIYr5XE1uV6O0JTg3504BuXmiti6QyO9b/C7XZx0LpGvv1
ogaSqHHXSkIeQa5drfp7y2fD2UQhNFldKPbh1/sGi1VV/+LM+ENDg6HKm81mHQJQ/RpnnAN8jPO+
Qn462at4bluRceZoWYYJQOtYwtBVOPEyJvjA9gJo/JJTzHnpOYUm4MWyb62RNwRpTyHD/KzC48/C
ovLVo3w3Q26R30TnOaWEdXJokPXij4Q2hA7IpAKwA4pnrMacJCrGsnuFo4wuydRuRPDO+DD2slhL
/u5bpZUU8mDvgFrANiaLVSUIIp37S0JvIiS7xW6uCPx8XWTfAxqDF9BotRRbJu35ZDTOXZ/V1d0J
m4udak747ucK93djWZaZWyaeISErC3Zc9DkLeIHG/c51IxY2YY8gaM9LTjJcAzLL93d087dQAYpz
t6LMCzj5SZuUdVVYYuCgrJht2LK2xVA2JQ6R5BLfPNmp/6TsyzA1grP1hNYdedZ4g5GJBVinwKDS
APtN9aKN1pEPnesYrz7l02NFjGhCeRN34fYIbREOcQ97P3gHuNAD/8scYJ7oNiYvr0kaajzkixRj
LAlTb4YohhZRqOw97ZmHPW3Mc92pi6lBnTe2lm+L1kbaBBcHuXLLzMx3LjxQTkqsye4c19KJw3m8
6Y/I5o2o19EzY7jdoX8V/IC7t7eF5hAxJ/d4tkeXKMDuT4qvXpDdH7zQ5UTxUlzgkqpU1dkg4r8B
X8SKkzYOzLxyQVFXjHFx4Xbb1Byix+sW85cnrItuAmYfpmCBCDUPWeUckqdpwUZMIPp3JKUfm1t3
PtIryMob2OUaWMF1pN9cMRMvNVubNJ95+Tc0KZzCh/XPB6gZfYkiXYRjAO8c9BGrzrpexDMEn4qo
77IJ7EZrAtf21zusw3EhWotZz8NadKBVVrFJVSYwBXBOgXhUFhv/NKaH1x85CTsaNjLnD41dmHnX
NHtMons8LHPD3tHaFaFvh7JrzjZGJcwB/MSL9s23RqeNwNLa4m+y4C1uDxJOm61VbgfYXNVHACSu
Jvj6cnxtVBcq0/3L3Hl2PwqsQ5vw4V0aD9Bpt/Q6/J1dWL9u+aiz7qGcX8kwmyIVTQaZxI7BhbK3
3m4OF/d2dGtdteacnfLJErB6ggxd6OdAshM1NCI6MOCnvms/6duPOYgx9pqbjuEqQNmAstZIFoxM
QL/kHaZo5vZvPFCpjs+GfaZdYk6jY837Nt75QGCECfKJ3WKN+NDx7pbOtjZ+syDgC3xJUmOJPa8s
yHdWZVDKp3TsGBNqNDA/XW67mlyERjFkHMH1Pz0r01RvtS2buRfSorL3bjAAaeMXJjiPZw6NMjuN
6ByYG6eCNLXgJ54lFIGzeQNCR/p48xWuovQUQvKeWO6AS8/GAPCasgHJ1AcuZqXndM9J8H3uRaKG
zCzAZWYjqtz+K4ZUB4GjK2er2eSBNg8BTxeaJYbBCjfT19ixxxWnNfYSZ5e4CUiDx+wlJLer3P9m
eqf08+FtkJwk4I6K2G2deCc5GdagaeuSbhWTEaba7hNjYVfZv2gG+moVAfmc7dVZBdeiJfVFRadQ
FmCHsterlLfN8Gv8SBILS/irX+CaG+KLbZ7it+VGftYQgbmZWJXIrbm9ZzvuNJHsvd9tumUBDscr
NXVcGUukF3vP2ow0fYwp5OP2SBkq35pxDRAGGkajg40WwPJ5VKTtzEiaZTLYfvE7+hO1szqUTSTK
t4S8iBex2/RLzaTJoOnp4J2XU1WE/N9aqjPpBkwu6pFSvrXKwaZd/JkzeyUqjkuUlGsLZVYQ5TOY
EGoKilNZEQpbUatbkCVObrQBGw8whGNOsPBW3R21S8TRH+uoO2vuQmCxexc0Fv3I7CDiGP6mdS7+
3H05P3EWKzTGR0H7LCGTc740xrabEVpEU8ZaSPcS0p31xyL4YBD1/sqZBJmQmdkbMMgBiU6V1kJS
pZL7gb94DFd2t6sHfZPLrB7ECarZZpSDmEQvndwh5GA5ayXR92ifbS2CTtGYd0a9HOk4W1Eyr4+R
t7LlUhPMHp/MZTT8WzBBFXQ2JdE83k5WqW/XLeFadGoY2LXzU9YF/tVRMNRmN/FqQkBz1LfiajCl
xEFcNixu5J1c1bn/AfLDs2dE9+n0k9eBkkKZEN7h6O5OlIR4hALS/28Xz6Xbj+yaWWwq9d1umoPR
fzFnpvRu294BrZmRJtmkmKLZ2Z6Ir4c72WMv/jfFKrydT+rtGHmcnV9NZCSqfyl6Lrte1zbp5y4t
UFjXDXADoiVJW8xWZbxXTb1eU/zq+Uwqb45biuO/O/yfLfAZqV9Geyeu4Hum3cmY6QxhE+o477CB
ovsU1lJDk3M/g4vZyJDnxVtpu1gpippny7EPI6FCGR079R5600tNz+k/TU3NQ2zjAspTjFZu/Anz
sWwbgnz1y+q/XR1U8mxbmqwZ9e9c+IHp94wyOVCPW26wJtDHwuT49Z7IcD6PVpuXrJUl6VucG9Py
hob8hi5b+UObj7AOcSOfqHi2211XeuUowWUcAAbdDRiwAZULynuRWIpIXSgra0b9zCxPrjrFP59O
EdRdIzC/sEiZj2+J/wQczLv56ZURU6HuOHVrNC49h1iP1QFATeebdiEsrpnUXS2nIB4maCjhtllF
bBNP6+QsOgNy1Q4eGe/rUE/L44HPwRxUKcSMC5d3ZPSU3dfyaQ3dgKzm7ULVfY+zsg5bYLfQMg8f
vjcs/0wzFEALHrHMOxn9V34GQVeXJOlc9czPrEMevgPbpkrTjnmkC4LkyBNiIEg1786CF9Nw/z6A
to4rBR2QmisdombdRqnbtS8L6ArXPVL4HEB9B782Keyg+9KXrLZeZgmyG61MEvrUGoyiCm0UcxsK
QDwIEW5/6Qgu4D/46CAHrUU7pKtbt40Mz5Ju9JbzW4ltEDfNduCQADs+BPGU6FfYfwLlqKjywWX1
ChnHrhhhm+4qC+IitI4e56gg7ZCHPb84lAJT/sutbPVbV5+9sUB12zlC8+/p4RqNDgaMqQ5liLrn
mB0sZlBr4Mm5YZxmEbYpE8rJqV920nrkh3BUWN4g47IqSpZ9ba8Ddc91KzQ9BOte8Me8tsHcP10K
Z1ZX9rgOaDhjrRQbN5JJHMMooSB5jztTplRPHNAj8LcFA3dLcWKvk3RgorY5b7ygBTFECYnXY5KH
gTCjPuCiJ3nfR+PkUFaY6klM3dQalE2MmrUYIxwlyi8tL2NeyliTSbOx02PzGMf50oqIOt/35Ba8
MGqyTMFYW3SyFE5BQ6JZPEiO27HYhdOdYLZD6dvHogsUAQZmJvP1fQlfYQjnPmw5qEqST7NtOtVF
QcvdPJsK3TzFkAAZbJJcQIWjwNl7QQ122UfPQorfml9gJHsSIDc9JJsHMeaCjIFaq46pwDts4x//
hTNGnbgH9SVjc0cLbQMUGGpOeszLptjuiHrzIyN+DiBxD5i7bVoyXHQeyc/C2ODKAHdLUeVE8Q5i
orsAZJTZdSsL/QURyZRdebD3gmK/Pd343tUzMrRUAXoX0GnoaCCRE6VXQU/8bNKPFgOBnqX/iOLf
x2UlUPmf022uza6lfrnaOFlOw4pfCXU6F745QnoT3sK3A9+QARrjr9xdY1l8lxXy3cOygRgbj18t
qvu2pv79xn/yEJVzsGqWgb+yzZH0zG0ntJPjXRzW4o0CyMmo5aA2uwFl7jlP3UnX2Pq380hf38AF
lQBDhf9JH63YxRbHkudOPMcuiSNFh9WmXS4U0CsvTKZhMQZgNywiEIKvrCvoTzmXwVMi/vFKsQWe
fVyNUa8Wqa/u+BQrLpTwNIRzPsdPSmJaDlP+POY9QWHRkgLBF8DHgD1sxfQptxNjWZu5Ht2ASDrw
Mrs0V8efE0izwKkUT2IyOTe2zqSZjYX8eNHXNwGyBUlNpye7fkkPzH/U2rL9FutcR1V6LZ3h/9G+
G8QSOgFHX9dVSQxMx08/8bdAG5dRpf465K9txpv28K19MF6Fq06bJIsbx+5/m1GVUp77tf5eS4fU
/xR/6u3/b4sVmt5YGyFvw5cq8EYCWD47rgcSI289/nj2vZXxS2EQush/nboePTHtQyXnDvvQ0Kcn
VgBJxI5TwXR79HLYv0Xmb9gYIFwPbN+DVOTRjECULM9LRvN94PdSG76npEWg9fckn/cj/Yhl+n2b
TPv5wd9SZtogkvHa59FW82qp881ftAWjpdF+CybJF8waOgGhveTQxgStjSrmVBZhg9uz47XYqM0A
2LNCrF3wWq3FxZbAUlJtpW4BdiQQNDWBTwrhJyptWCeqF6BmKfusst9L0FKpNlBxvayjUcLlLavl
5yfJ8bmF9TidoIDGzmliIIx1OMQstqgnrtUYtC65+MQOvBV/JNzZH1vJ4matmF8YIiVYVb5fIwuA
A4vvoLFb1y647GO7/qeL0Xx68x1+PIymkYnB5F7wKRVi5vjHjTdIFIXT3jW8YLh4X2++DikdjGz/
GoPDhgH6WSOyCW83EqQ3O8MRc1fw5ZlHqTxtiGdRAG5ETCdKD+SaLkt1noCfs/vuzsoVqTi4SQaK
G3YLl6KeI74lk0WMBscfk7VH4xEHkrysMucn2WFgbGA0YdIkgV5/wO3j50Bg8Aa0QE60sUs0P1KE
W/yWURUaSFjJpu++RTB1lxVbvH89UrWJyGmaYgWHkyTAH7h59HZ73PNbMzL6L08juC+rW0rzXu2Z
Z3Il1u3aY2EfJuGJ/rrnFye5XusE4Z6m7pSlmyzaOoFT+EUGouQUgbTJCvJpdg2I63kdQKoo1Htb
qVB2YFw7wEEVg8htbg8044NNNyNr/0gr133CaZHnZl/UM1J78+ccd23f7Nix/604YnNZF2THSNfi
WD0Oxu1VYyWVxytnmHs/OA0pp8jA8dKhTUGA2pO4XYW93W/jZ//RYWR4cThWs/cHKaKMx+M8FwI9
/5DxBERZyg2oNaP0asF0VUv/wbOt15bS5CGH+CYIr+MEN60cHLrSWsykZUt+pmpypf8jbcQFZuMI
Wx2AwrPuWbr/BBdW6n1VBXBDgfgFvig1s7+SEcTQK4G9075PgyH+xzbbu5BlbPeU/NpwqvSO1B6m
wcRK3MBOZi4iWzKewXozK/whScby1hljGujHG2miI7RyPwa/1Ql6suqF9Qyhfhggs/shZYCQEULC
U7K+1dfG1Rnrc1FaSegVuZLxvKMyTDHKiKsUNpow3gGmP6F/WvN6Iku5It3DbS4C+4cZEkBPPRM4
5YSqmAmxM7ecfYarDqkPBbXK1H0pa+yCp1FOr39d2YL/UWHFpeBBpC7XBYARtcsCtLhaNnedDQ6/
qqHoIVFLLJZ/ZAsmzClOfogUbVXQxmSSyNpsst5qAbSQnZKV53nAzJl7UWrX9KvR3PFCv/4Mg2RT
eCbi4l/nQknvSUSTBYrUnKW9nZ05Mgvw9CAjoizSlolqzz+YTDiVKNnDA4ufQ82aYRt2bDRR9AZ0
3mGpXvGoBomqbk5fpHvmnB/+RgHB3r3QTqvQ8CIMio89h0ejpBkubJ3qY81qclF0albpkfH6y90Q
aBeLz6N83LEjBbDA0FoCpXsyemdKTD5/AYdyk8znGIfWBdKUCYJjQ5cyGkK/PcWUP7dOSx1FHOV/
fm+T9GTv38AGWXL9SkDynVfMyV3UKUjMGoqkD3D5jgYqLGm+LCy8LNANpFJLex6aijsqhB0Hb8fw
e6TDForzS15DoMhrHk1SzhyOUL0W8ipkdWo7Q58w1qDofbz7c+ZqzXx54MssnqkU/0QVwdxgP019
ljkytoAQMOKM/BaNvk56XOgZDxY4gAOJL9xVEVAMa68spfsEdj/bOsutIhJspqRHRHK0KcLJpbE/
zod4xPzE1TAsYedYMI5308rZQA5Q5n2qvsv0eyI3OD4fxvRYwOeh1kZuneEn3LVYbA8hne+igY9X
Tr8Dz93+6iPv5rEQAH4cjDax5o17a/r9s0is0sWvnbYehSSmrdjE+sVNlAnGhciAONQ1h3g5xcKW
E8eHq3NORBPngs229Wj3R3i89Wt3In5TWeScKb/vGCYlLv1xed+OBgHPqPZfVaq8Mp3l3RqhXuRC
xwaU1bwLQwldiQB/8UfX2p7fMkt0qZ4lhaK6oKVjmzRoPXR0wXPbWlyEH+SorMUInSYPKXU6wxIP
WlJBJqdeeJQo+0Eyw3eGmudvfu4os1Ary3PbqGpWkeGRnlue21vFi8jVEXS7effSEhqhOGMFFM8x
UIOKctAPXlI6BUiTFygwx2ILrSdRDKRF82UUdPcs2JFyBt+w75gHuqdHzWinxL+iFd4J1EGmKp6a
P1C0J7LmT6Hw6/gG5BnNvR+NWYJ+/LCAR2dYak/V9wrYQEEIkfg/pifY+O+gKwxaGVDi2Rz57q++
56l4Mt/nTiMb4XdcT+qyQbm43uFNck64YkAgvHhHgMMm/s6SREkZENy00KTOGMYrm/bdj/MR8yUz
lVsPS+Dcpy5iK+bAE16sYlBcWt/VhImmf/KyMNxngdA2+G6wlup4msf/312lQJz21DtpiQZpLE+V
Tm2aNe0KaDh1ozgLtcfYHe/k/gjp1Fn3hFMw4ElhI8aXMrOvggcGdKNYQivfsbuozTjI9a36JRal
pe2PAKh6/qJs04vsCNYTYi+kni1w5ZrkoqkXUENMMxUssMK+pUxwQQOsdhnJpIETqWj3iXPv36cw
qMGelO2tvGTbhtNEl9KrKZ5MLoflxnWX+DdcnwO/YiNHUqLVuMmcCgS2x8Zxxps/JqERpwC1W0C2
XVyIr7JG0dFZznscfkpPjQ1sTZn7qhDoXs7j0VkohmtsyGQYqgodxkxMHJ9TxuTxSRw5A4u57fv4
ZV0j8Rqyt1EQB7QCZ2hvKFq7EwTH2VeYp9REPDqUcLXBUpFuAnzRVrsEopktkPm8iRrU8IM/dETI
bwDRM9pHLFHXAdrSYqdxSjU6D1dPsoMjY14cBsCQucE1c/PJMd3pAzwzLgftjjSRWnysvHcrszmw
9ugv+knB9MaWdWf5yFifzM3MOupXfc2Z97iP9DVKj4SmaIVYWK7cOR9J1zaH6Tzdl7Boog6tX0pu
VHNTBuyIGBCyrgXLThdl0qCIv7T4GouBiql1E4NYO6OGgMsDaoi3lsgAYQZ1nOPk0IUlWRuytzL/
dT0PjS24dAS6R2/2qG4lz8G2Wv6oCeB1ifzf10BJKSBgHPTQSqYvThwKpidtWAEItIjbYZ5NuthY
0NpKbiJuG6ECgfTFq1n5HdJoS+PIKDPPyEjapV3mfNzajBI6+jCAInyQUrzyvi7oS98MW7gVYriV
7SEH1Gd6CLek/fHK7nZCJevL+qkiC3zSFOL6j8S+zsivHYp/N9EVk3/+s/ZjxiGDFuWu9hNRaiIA
TY0UCso1WtKuX3eH41KU0WlcHaGpx0QFACYQS3NfwbRAy3sCPBAroZgeqY+jJOo7uicVoiX1oo1i
RWyGUWjzt968x7UAmYecCJb9h61XFErURpVV72sUv1ZcTDWjBsZS/d9+Xa1b7Z46vVMcq3OWvjVR
itidDrkili2prlkmWhop5k7Ppe7QFYiJzcYQjvTV6/znpEw2one2m9g6uXLDuzHmf47BcCXG8hWb
LoHg1DgJ6o3cMlvdHN+a4HlTcDT1Hy4o9bofUIvNvwWfdUqCT3aDH0J3tFxicw5Ekdo0+i/wXSXE
UTSeSSlUBSyDv+JkJk4Wr0+bi4CEdKx3qjssfp43dGkJ3dv6z/CCSBua0vxBThvByGfK0BjUZx0A
AM1v3zJ+y6KmEKpi6E2Vw5V8XtrGjOueEy48P+qiUFKcp5ef+JqnukBlrOIbWD2s+rn4G2Aiyx7i
VKHT63AVEfaOyI/sTfbpPrrFtauBWCH9muYNKC32A25ajTbhQmhMkNgQ4Luwf1FHDRo0gvKIDWhM
hsnixyIvTX2lWwKujbnOUpwT6TH2xb7/U884BvlQn8b1ppzg3JTrBK9Igk+G7OjAa+x90lbfr8Qd
B8Yxr+jwAef+xVERUzmaL4SF+ISBgVVRqRwdDKL7LiCkqt8wC+vg/v3/MDh2cJeZmxE1NbPucMbk
+qZ7aVC3Rjxl4S+eKiRMB4aihM69Whw0Eoa8L0WUvFqfiU66wRfIx1ykNplgnwO8CJfMtZUK72Pl
B3ufd82dUXDnD5sp/mnQC7ZA6sl+1fvxwhJnYpm3bRTzSHt7jtSWE0ytrew328ajScHi4R/9+hyC
8rIBYpNCWPWuR6Fr8LR+bcQd3042RmL1aE/6yfP64l3H++BIQBCyoowLRYldFcHT05APjtg2TB2X
f4j8b5E4PbLu2Cq89NVLx7fUdsCegMLSHMyGhNiH8OI9qrBQ4yiw0sU3Uxyll6Yr69SeO/n9naMN
PzM1XIxkNmiTKTXdOro5s8ExfsdV/FPiWF39auexI2kF+W9o7Iss2ji/7u6kArBi3cXm4xuE8jMP
SWPxxqvwV8EU/BJFPZtoIqtAgiS8ql2yFtQQkNMYxwEunrXitDK/MM2bjc+Fiha150+/Xh9l/kOp
AQUBzxby1mzuohyffRBpeGDkWZRjlXe8PkaLFz1YLqww43k20Ey5IruipMSmSIXoV0OoNmMjBqco
kA1Y+/3nKlZwFMVkfDQR5pg5iJBPfxDaLK578dz8OW+yM8oKvXJnqfFh2fbIqTbz5OgXt4SWTCWs
P8PkyoJjLP1qsYOIaDsANdkoEbmGwxfprIc4vRTN0NlNaApqZCjffGDdjzlWXQ5xv3u80mIEIDvY
91ShQE8YJuiOnV0mCmXvyk4SUAHAvTEED75k4b/dhldFk2hsOy2120VIcEqywl1q0MIhN9GX/7ro
HRns2CliN6cbHE2d888n5goyu0TwhEr7dWrhdMV79NptKctwreWdlXU7ft7ZP0S7Z9PG2/KiC+px
6TZvnHT8rrXNL4e+D9t7mFzuhp3v8wJISa/SxyRGX3qBIWd7+qKHz/6dVgEyfzAVy8p9Y/nPZmza
oeCZ2vVZ0PjuITr5y1hLTRZ5yby+oN9tvYZLMyMjlwmfiK11TjEXZbqScxK4hN5w116AZpKm3Sae
/ag/Iw2VS8r8XtVEIgt3aYDLpUel97Vg4Boq/mYE7odZVKuxLNEJ7ajuxFgSRgXB90dj/zayDWgl
MpCSIyXHGuMar1vjL1iod09pQAi+Y/N44xD6K4LHlioMw5n//IjOTNrwHK39zMCJRcMOe4E5s8jM
1yP0MUQLbdEb57ZbGn4tZetCVng/ZuJJLd6vNQcNPRknhOclcQO12OKwPK9tVK3cpEPMqF9gzrOB
GEkijBmUVZaLc7In+S6Jk3T3G2AFQJagO2nJQqOjIMmGxJCgIoCxIJbsN57xudM2NjuD0bGdhfAk
L8hEHgiROAK1E00bs5ZaeViVEND5e+ffLZnL3/8SIhrJgO4NYgjeqcodczMjLrXK5la856bjcbXP
qvzfBK4GfQhXmbSSwk73Wmf7Cl1Dvit8yEhJHYqFnaHOYjZlMlzxF2EQdlbaIKMoxZxjmyeOCEpl
VJytmLVi542m8MjoOjj9SiOyC3T/nDYiXbkV4tPQIl0MNnNQvKtENzziQOyZmgpPeWXsiqQrnSkJ
vuR2k99Yv8AAqVKm69bIJ11wxh2za/O2pANSTYC0TGS94t1lvtidjexx83WuURWlgnRxuoSS+UjA
lvJhOGJEsukq1xy2vTKkfFP5GMSymZMxp45B0V/sLQMji4P625ueEM3VSukPqqGOYU5Mn3Po2Gbd
vuPqlO8+pMOEotTzC/7PPW3qb78/RZ9BLdGkVUBHyCMPs30KxDqn5WgyZMBOqA/Jms7+iy/Mvvmi
7HEoy0ZZ1XEurqSKqKMBv7fneKEuMF4FGJW6KF6EfgwfAi61+kjMRM7FGWsmTtYx05d6agimd6dC
kU8063mkrEvpUpJWOj4cIXQ6a6NZW9ipnLRnSPhdK6yoKNWHHIOUUWBdlPTMFbAujURLkv9HnFpn
KFmUopQdwZbij25uRDC2b2W/0njSZGbFSu8JV1Y5vCgB/K3El/kZeJS6tRg4SPcJL3biwUGxDVZR
9QUbE79A6kfARpm71SjJ1Pl3IfDJM5l9EgBEvgu5zcjJXsMPf6FaawK1rDZ4Xqq7XF9NxUu3JuOU
mDfBrOIafsZyYyDf4JHBqczqhyznDiToh8SLzs/5kS8zeqIrROPb+mpJTPwjYonk09tLG7p7xL7+
fmO62i6p3ljBkqkB95n76lUuH3ercXaB5TaxejxVtJaqEnp/7iTFd96nM5jsV/poPizfTeE0lJ0k
PO8uPAD1V9iEL5k1dn/K23EOplCW0qYLsj6Oasi3XpvIv5uxN5to30z3fal+/C/8QKyI8V4hw5jP
0bdFjnkXfB7Nx29ZUK/XFeJjraOJpSSZ8QMHTowAgg/jSVVvdaDLk79KEwZne6a3kmoXEDFLmyDH
CusdmNWWNmoKbO4MiDnNUqciS1kuqAzydjKsH+M6MMuo0uM4JLT/97q/CIOEPsxW/rel6RKW0KeC
/6Kc/TGPp02+pgm48ZsmQhLCTukiuqT7UP2qc4UQb8NbilHEkI2sSd16A9BqQZePf4Ww9hdLBdWl
+7uUOwLG//xHuKhamZCD/bVFq/n3Q5ZCTYBgP34s6Xic5CxEJBDDz5ESsepcrdDbKPPDT5wXLD5U
A7Y22GFhJp4EYuT8HX10Lh5m94N3+dH2ygimLg3tZ1T/MdZbJoNzXOYde+5eFj/8AUdbROUWY9dQ
FoQ15bSxQ/91TZCrB0YVZDCX3E6kDAWyQHVmjGFDhPTgP1Kher85kpQmsVEc1covIXX6jGE0B/qp
iowzXIPsP2WSPP8LG+gLq1+5zD6yo0yJ8DPN4gEFwFALQJ34SMMEhRP1qqIrw5Wp9AjeDY4xDV9Y
ZX6X0OcmUONESRcqtiwqBY6RsjQwAKNenHivoDppnsrU0Kp8Qq940ZwsjF3qWfDdZ59ovxiBDiY7
1gi3KpYRH05UfOlSrWslXDulrf4rrB5SgbsbC3hK/JwmGFeRBiMz4BqPCN4lPPPdvc/HEtWUjNpD
xtNrMgIJCNuMfPkBnXsIiY+QuXz8AOkbFdnMWkcrw30Cb1iFlORDGM98Jm9m5MRshveKmOymH19G
DDvpoP0G/ZajZJ35ljMCvShsLIXtkhKeZqii2nBdQBv8e71CI0Dx2rb7DauErp+8XzwITsG7yKsn
Dzhxrzl3oq0AWsLnSGYIH3XgPdMN4/tP7zr6e9QhX41RZdOPOvjosIQ3i2nwfCKJTqAMckGJ+YhI
A2QTVZQGYYFJfPzwOgTevEH53czDNVZXS459GTp6Be21oE6kDkDmkISORfBuwoPqXity5k+RPmOK
6QguWkw/Ae77/0zbdfFeazf/Nasg2DUMhS3egn26wmH4oT993WtGGgTruJhaRoDgKURhHyvgtCLT
xhqeQ38u7huxHUeUFcncYNx8o0kESzfgtM9aHRNt6rKb5y6DDhQMGKremqkoOT8MEetk7VMb4GDV
wbO8MeG0sw5xVOUDVqBQZ1eOCdQBEbe5WBM2JZIyK0pJSp2d+MPxLc7h3mBiieJULLMxAu3H7J+x
EF1sjsw1DRVzgMq6H9IqiIetyCfv+NncjvFODPfvcRprQF9y7nt5kyQaZ9pKunMy5nAuCo41BKTB
3O/aWxpezaUyDszYlET5TeiWG8lOQr9MwGOzRJ8L4+fTAeAL+rAOmpkI/kaSGcrjteoGu/5hz3+g
LazUk+zktTYwRrkL6uDV+K1PJwqtEYREPECEEWBlzN3WRHU5Veijx3Ewqq1Qz1DaR9/SGYh4I/hJ
PoLKypmYGs3wixSvbFp3lq558WEzi+rVwQW+ocWio5GrtkgQ42dED0PsX6ASB5L/ZQ8ce7Uc4nDA
/bUf4bKc3N7RbnrT8aA4WnyxB3AVrqDrGsGKnHglb1MHxLw0STbChpa/kHkq1FNekDfh1RHu2Ud2
LP4mq5eLCbzz/PHAW4PVnbc8mbpAj3+PUbZRhZpskfcc0oge12k8ydOb2sdY/U6vbv8Rf8Tob2Yu
kdRgrkRLE8RvW4hS1tgKC/lXihfgFkd12lMdpwQJLRQ0QDNpuCx4MLdD2Wbd1hOLdl4D0BfPwede
ZGXzgHVV3NcE/zOIOCi8yLAYZoVn6Ymm+5bl7UEp//ulHl30yqb3f92YTINqC0IjUmo0qSY68BHV
qF/a6Ql91GTyoXFRr7FFDcUHSLm34frjECYLIeGmBX0FpDyk3f9OFpTST3zWxfYfCDknn8+M9ZmU
Hz8dDVSGerIBC21TY4qp0rGifeYhxemC6bPkwj1H3ociNJ0dibEobpQV/apfigs6gBSTTAYK5hwR
+Uo6qdWT1CmVjmq1UABUaLoRdmO76P7lMSLh6LZzc+4ZQjzScTa9pik/MSUk6ViGQTNXhdI0UclR
tSYiplss6U9CNvg7wEf5Rhu2P9P3LVMUKZVKAdMMavABoqTL5EZ0FksjadBZKQC+QNuS1KnMW2aE
4hj0eJ2DHLGEJ6+nEJahgyygzlv2eCyZqgrRSJcSO9XTTslsGHbHaHcL411qkFl//rPdeWdfTPtU
brcjUsHop19518jWwfLJbpRg3LHKcpK0MNdeorIJHR1N2FnG/TKgyJ7Wt+CQ6WVNY34BxIfSsT1b
FI/jlN7y/5JVHXtXUS0vv3ziX07PINJpjPCI23K7ZslhEsCoIclHDNcTaeyhNMZ0os8P6GxO4lqq
1XpsMxiRy8w+mtdVUAtLZTPHFuAdOAgaHZSXKcj9P+LzA9x5ACraKb+lncFlDheTpmwsaFX/hWHY
D3lgqpg9cLKQ4HS9GiuzcN2A97KA2ebIxcyKbxUlvmwpPanMVt8I+BsA6TDcQBnsV7LVeO+xl3cr
TyeqrDhG18Imbj5QrhTQibwTf3QTkGRT1yVNrBDoWzyGLGhl5psy6hXocUJTM9fTGuDGFbkJwOCU
k0FnIUxvKQCLEINXZHTLhwu2ItsbnHKY4ImBau8ZqkPWxf8t67NPlI/3pPpr7xoCVEIaDP9kT0gb
AJK9tdnjJ9tvccGjGd8vZy8gsRsS97y5eEaZLxWaT2R8CXZ/fN0C4gfdfiD4InCv7F4hVFAocply
U98ZA09b8D7afQ5Ty6SYPAHCA6K+GaV11TBr0Lt/kWw60kcpHbXnQO6COuf/94zsHvMgVysbASj4
jfa/LlKaJG6C/bb1tr2NjckQw51l25L7A7MvjCejhZUIja36RkLIbL7xFghAeP9v+ETS6l3tyoMt
URuhp+iKc+Nv3QwBiIxj8aiCKOJRZgucFrneMsmkXGAaUdYR9uHyrZs04BeQWMbflte73qLOyo4X
UVjsudshdJYWE5C3IMH38Ubl3g7bgYI/j/epJW6xjYBIHNEp2JKVmDUfHikixndAsGMZJm7D7BVE
TZSgKcYrmREXR1HgyEJizOCJ5U2IdRxqflECXPr6/N451lPjbBMBjfxHpWqq9UuwIJXMbBF0B2M6
TY8CBrGf1OiC44Duc6ZGYJCEj7jpMPGP6hoG1cmM7Zjku1MSUQzOiWtWLB6zDURm6oNyk3r+IXOW
EWemXqM2iVdU7S9QCw8GonFp/NrYYSYPV9bsnnnCH6ddKYbaNRDBD3FFryKl/xlk1GNnvc57NPXO
jVUtZ40n43RrnxLoIkW2V89/+7gSivvqoFLiRhuHiYhnwbMuFSXkj7aJeo048gp9aCzqi5hEFEjR
oYuiQ0YhtWPDdArDY76tkJj7axzK476wRtLM/P0Vxm7iNIjXk4Ejro06Fe/rWr/dtYpeUzb1ltlq
oo73i1/iGbFNDET1c/Uxw4lOpuq3F4bDg4EsRftbftOGzS9YoTZnNxTwsy8bo3cGqVryvXcgJGJ0
xZxC7l674yYlJ/W1jkumh4lumrqvqz0h4HRQRI4T5Cn4OeeIyVxwEK/HcQXx3GXyo4BrhKnqprU2
tvNk/MWfwkVO1VyDLkFGpQMy3nwrHi34Rrm4KBZyqFKQXUIc/0IcDi6X29eLGVHMtmqZF+jmz4Y2
sC9sjt0xMuz62xd+Q15H6Bttn4rqojt82BChdh4GuN5+r1PdVJ/iQf/7W6OezNXMQOWQB3tTsQZG
qcnng6LFWI9SGm5/rWe6JzzuencdQJPamPadOa5NT4A3EFClPZcm+8Rsjqd98lB79KCU5uKjwReZ
jDlYFSP68MEI0XSONcGIYpl9JTPqK23Gw6clcO+xBh7NQgcaB23g8aYTV3+dlwR7VuwpiU+SLFH0
KOhV84Nw2/DsELQkbk2sPHc/IeRSzz9G8S+3ITUACmPb4QR1lEhjtlZrhZUHxwXxbv3Ma6d5HCvQ
kQTzaZfaE5mbprli/sjAEryTMEf/au8qqmPdmlFU3IkQeEO+uNY3Oulom9MuUaJGbLj1cnI196f0
QND4ndbX4PdJaSyXCwsvHeKUR+VpVvG+DbunfZoOd+er1DI1kr+PfC08c8F3KtP6EHXGNB/Zj0UY
9NoinNqcFjx4rbxZL6IOFKk5KsAcSD+UZ05rtUDVeAzdpgFm1qfVu5IeKJagM02t7oVGAwWc7Tx+
imdUEcUcLTlsdQAA0ztYu7+bx0X11oIT8Et8ynnDCHivZT+KpeJErTOXJm2+MRAX/EtNaCPFWR9r
H+/zwegJW7vPtBWgyXNIza/6VIirIdkbgiIOW9gGu7dt+cwEmf27OtEoeWXhHxSFQ3vtK9IxIt/n
f3ADsz9a8OnKuNdPtuMmiGGbLi/KpZUrVbadJdeh5F65oGGPBgBMirKleg6PIijjSfa08Q4X4Nvy
XY6uNHtWzNfjiASYDboTldyaOx9bg8hTulZoHe7OjihCHLvUBmh3Gi/JZkU46alyAO01j4arsKME
TAVVfkvZpcC7PscwpK7KRq/dMiLyATZru+WY2hZWIcBHi78HKr5GGEQN+JS5eYAJSlI0l8eBOus7
DfWMP6Hb0sGm7IB7GJTtFOp6cXj80oxtqoYo8zMpZDysTPRHt/MX6+mT3QoIhTNgtmzBq0OHQ6GM
MJ00xjliUqM8Y27fDprC+b4SRrOwWQPFUFS0FysADJmFLj24jER7T5LJQgknj7uCD9CZOKgGeJct
fIMQdxzaWZhHvvfvZJIAGuhik3rWG1g+wLGbSt/FKF1raUMM+Z3xBCCUthzjj0rV6uFE7dkCOCBE
a6oM1Rm0GlplYre3k4qCqHafD5ILawoY0XWJYLUNw77ENgqt25vd4unUqzL8Q3lBq166nlkXhTO3
jxvs/XQtVsPV0XNhB3KCN38RSy2Mj2bQL4zG0bhyW48UAz+N+93SKmyNTW/YPpdMmpzAfpVVNJMX
VKA44hkWIhEfhLnc3g/xgx/fVHFW8zsmF8eIbTiaQtvYRRISvn7CVmimENEhhH85zph+jl5kpWUf
m6gcOKgeNrRNgIAAZP+N+W0s9TxXLskcLEC2ikQ1r7hoXYpicPGHzoC9YamaEHQsn2pqTmbcqg0X
HyDn0LPPDshysO58LHEz4pglwmW8nf9q8IMgTfhWbE71IBaSli5if7KgUDt6xKqq06rFE7z8aEjI
YnVrSRdLwklQitBDgPa4pwRHfOVSGUfon9Kmny/5kwYaPBQ7QLO8DjqK67UDtzuJxd+FODuzkb5H
hl8CeRHwly16RFu9Vdy0wCBtEUHVEhoinRoaHDn4yhw5bHkkmyFxegrNXNuCQ/WvtbvTnPxrt5/G
Pa8oR4wwlwo//NFikDNXr7CVml6EAIA5kZtQDZvI2kiX7LlkHF9MyNHIWhu8JvX94U0pad5YNAQi
7acR4Gt8hVp5bD5Q/9E1JoNkiSPmnSLceowE6KQD7QgegO0/Ykwb5vBvj5ZkC0S4lbtiDZBXwT2F
iWuX7JdTZg1g2KSqvJFuTdPQMnQiMIH20wzZ2TuJqxU41H8QD8K405g95aBfyML0SwkrE2m/CQgV
vIUQPK1C++5h3O9blyTYWnmnt5rhxgkgiKAKeZmu3pt2vddBgnKVXSggYklEk7Zz9tc3YihCYlft
ZjMo7YwkwCHu9aidISkdUYsxNcwqDhgfqKP5ybmEu9+492qHsZilIS+uRmTR6tpSIApXn5UrIa/N
Sex2bHoW9lwd4+S6lc7iEdnWE26+/rSnN7asxCDTrfO+3h951FMbKuaSv3+x3kAc3dPt0JjRuQ4n
fs81I19118KbQVpF8dg4f7X3mELBjbyiFMMwLW9jVblx1Tn6HYp3Ubomq6OqyNfR6bbSDCSA74al
n4qq3I64W5vPfrnmwVkHZYSgr0ZKsP/3lBCfma8LHGcW/UkPQ+HhBRINzhn7YLtVNtHJTokjY89H
BL+gnoRPKVomzvsjKVSScxKy+moqFJWAqHB8tJ+i3WNRS+ZdLv00w5YBb56wV72V2WCs0HCZURaj
y8leO1hM7uQF9PWl+Zyx8JXhHAJPPTdBI6l9Tk8ANhG75S+vT1NOCHYtam5ht3cM944ObLaa5CY+
e9IjInrHyIRx9+l7VqgY5EmFJEtovQ7+pyHZRG6j8kWMg7jHD4vz7d6hKBX+SE2ykrPSjmgHhHs3
nFNOt7EV9CIAaxy0x/uEI2TFoLw4gfjFK718Q6An12E78UDp4e+SyJRln15Q5p9KdgLzd+KVgXuN
6UtgBm0/uKKSp+MCgGcRkokQBomP71UWwJFxBmme1ZiyWn4dTGpFhKUDu76pfOzUXO/xSlWBRHOg
Tv6fGuIXcSKrBe9q9BmIgGMX71Urqva4JZF+Vknb80BlQFsvsCNJhz/3eGvw97M+O2tJRtfxoIGk
ajPz3Z/PUAnO273vKwXAUw+G/oTF9we12AOds04jr2CjzMadezKzW0903CfMsbiIqo4QutYi3+i6
M2Rv1w6bblC9/Gfc8cggwZ178nsvXc83fu43Kap0hRvXBlmd2J6JilXQ61/OIUb0v7b/355uAciP
h7XHx0lP1AXVue83fvSiRgBjFukuf1mWS49g1fbtMKz7j+UrtfpxchLW7uMdhP+bfO9ZLwUTMYOF
Tk3zTFhpyoZCpbU/D0MnSKP1Mx9ZrtZyWqXHSzbMhgUmJwHmzV5JIEbzfh58iqPcXaTucpIzUzlP
oM6PZ8mk4AInyv7cIrXtHXx9EEk1AECNF+YELAPe/RyFkFvL+TLKh4Bf1mRAhk2rcb7w6U5U27gc
b+UCQolgWpV8PnjhJxjpbj59olBU6QUosUlPtCNjLcmwbDEPp5a4aE4BJOJM/14viW/5iZ1rQKMm
xBYy71iENID++ZnnL06qRe40/zsNXgeQ1ir9VT0jFxCgmQMV/KY/nh2Nnk8SCR4EyrCVhbK1L1wT
4SzJE8iPKQ3eSGmdk8e4epRwaOXXg0Jw0Es8PH0fBEbM0VmzDfEzV/aAobajEJYIqPclhnjN/IW4
JoCwwsr2+tkQKd07BTQZjZ+eG9fdxGkksTSLf4S/Bg6gMsjQch/MWaeKaNx05UHFS1F6N5kOYyn0
EMKwBVoTRLKOUfnQKm8TYf6KzNgETSf+DIOHnUHRDeZk6lAkz2NBU60klsUUZdv3CXSblPlzVESx
4WeF29ZLBvpEuvi6dFPFeA/j/cGUJJj9lmTkP5k/Iu9bPZ2HDm3dsTEFlfCvI4tVre6ru+XQeiN1
di5rDbs2WKtr4v/2yCHqos+9Hi5et4ebSEH5Il6srcCfWJ8QDL8sqwsPYDrVZrsTIiQbylIXPEbI
18fEYl6dOq/7a97Dq0dRUlq+GV5IGR/TWD8i3J3hCObabnTISnVKL/tUCPsxaUSSNJfSm6+2UYh8
xatEsdVAq2MeSKAXElge+7bF4LFggJR47xi0XBywvSk8ZnaObkNnEZHrPsAzyTbCaR3lYwVVbID0
gm1nyNuGp5FtUuIrqbftiT7xjEjvvXAKzdZTkrlWuj/xDLUJhwrnEnnbND16DWbSmzgMCLaPj8EH
tF1JeRhp69JQ0Q3pMgeHSHJ/dNdkKwK7Mm4WaXnJ+u0PgbEUjg+UbZImH+cWw+RwZ4CfrbjNPQIV
vgxkfwX5152JjOlp0oPTFYZ/xin8BYx0NrQqoDRRQrphsdnFvbboResGBwy7GLrdGRSt5r8Um0El
dDqJKzlTsSYi8TP7tknzOEiXgV3mIL10/scxbkGwJYyUoeXowtFgdjhgNSHS9c/PVaKukJ+RBlcZ
yIEwDfRoZNcw7z5vV4aIhqZx9EPSY0ebSDIimyYaqqbxeWKjhat8EiDnaMglghsify9MPAn7cm5V
f6Y0PFgaTP54XACKHghauoaVhe4vp0C5XWLlq4agohhzebbihFSPSwl/T6k/iVf38GiBF7GjCtBy
JPP+IQk7IiHz2wr8S55NgEZvBTHMwwpXCJn2xzYKqgAR1JwwoWKLNCHvuneFXq2a8CAOm5asm/iC
F3Qv5njoOi/0QjFaRLfKPJeIK/m10XagrKZhzpMxfs/Hns1ghzjCtJgQlq20WWWSOd3BpZYwvqXf
Me+UNS6jGJSIC7NJvrceztLHeGLNWrx7r1ovkFk9jAg0AEdvRPn2Eko273Iwa3934nHlg9Pr/n8G
gNrmabdkNPLpV1H+9fiqoyWyQUiT2VAVfgwCPRGqq5nW7x5ZiIA6QV1VH8WMRFJrwZbQGr1fe/ly
FMERYgACpP4RWlv+4ev7m36rPxOACicafkPgsyYLSM5OYQaA/Q4MQpDlN8S3QUj2QNFbLp5RTnFh
pNxvGBvZHhGUPV39WUto8myay8F25/SPOXB0hWUacW/wfVd7t0BSTA/gCtAU5Are1nhwEQJP+rx5
Kr0/Zy4Q0MSTb1ZlpyDas7c1Ye5tdDFz1plSPJXlH2uoGFpyp6AuC2dc0t6JszUs7zWpPTqL2uXN
JAOQBxo6LATdH9eLPydAOY0o9y1ZURW3oArgdjxoXeombbIa70k4N3gevVZPQTIrlsT/5cfNT01x
Kjh5rKZF4UV2qgbSthuTGyLuMK5MHGRzbzfYb3uYlZ8kT8Xbob55DHC60ZvU05S4YRK6sq9o/rAA
oDwQGJgqWA6kxo8Fe6rb1iwHaePON/Y9IfVam37WZjTU8GBRaH0Nd2HzH2P4I7EUJc9b+qzoyHx5
Gfq7+sw0SIjuWOJe/b4GSZsdpp6qJg6jmzUiWH4YqxAHzYW8d+ZkxEx8rWWYosAaY5ai4x9rL3Cg
9bDPJd+q4nvPZHeu7Nrw8Gi1rPI/PalvHU3WOtV8ysBr/djWSC0r4B0DKyumgt5oLoV/VTaDznkD
NhsgUYWxRUmffdXkjKSaBnlJkFsPcCzn0lC5HqioA2OH/rpl3VDL0zQk6A9n+DeeL5iNp3Q9yEB5
Qd5TCX14JuHZANV0VZHDItuadrVLt92H9ETODYZFSxQmkB74RDDQeNHn6c/546O2h/Ad47OAthvQ
xh4OAkZYHq8OVdslvIO3Y62K+kSNsq+WJEXH6TCpJecVziASU4hGcFZeWEo4Vv0VDLXBz0vgoCEp
P9a2bysY1b9e7szGg6YlZVM/JEfUeri2MbbwZUR65kHLCndkubszu7bgTV2dQywHb/mLeFexmI+G
9BBzemO3iJW1kSyQ6Qi85sNjzy0miVnU1wqs0/D6cPvsM3cbN6W9r1u53LvGx6gMwKwiiWyDaccP
MSshBzhLD46q2d/BKFYfwaQvU1SNvnj1C9K9ozCFNh1vlqtgaO8DU1kapLbhgx4L/7PuD3kwSobA
id1I83DaVxgNiZDkF73l3IWspN37SEiIrUfZdK9P6lqvDXZ3ZlMg8Z4E4kWsgIkgDTUzb5znJVNF
4c0kukeDuogj64K4LN4gPFzns4pBUk16pZADf2jakBKDuW++MpYpHB1Px4/VD+XbJ5U3rmLgmqpk
nldaqJGtbbLZwmbeI2mUk80ysqif3RrT2yALq3itMo2WFdlNpnXqU42DLm/sE/+slfBGzr30/3tg
FU+De5p4JjUivhsIErIf6d8kLsNNI48XL4RE9S2VjqOfVKLxzAh/qukocF/mQLvVaXmIixiKuYVT
4MHM7onBecFYb6J99YwDiyWk3PF+WHAAG8mN6CxcBEZLtcr2edhdvoCAAJrTJwWesVynKmAHdYou
rDuP53ky5Twd0kInwSr5xOGYGrzsW/wi1ZoXIreBGRIXBXWXV9RU7eGapxa4g4R34AWJq9N6ND9y
o2opt281G7guLxJP0+/ICCKK0Vm+TH+0F/6mqTjrasVp45oeIYysRAV5F9gvdWMU0UzTd+o6cUXo
B4+GUhg7Bj4fXL41N7mzBgdps8hiETjjBAwBVIk0mZzO1sbcDRhD80R4CkT64c8Pr1hZMbt6Vcnt
/kq1nT6CS1gP1uOsHPknyE/IOb2++XEc4uUPHjp6yyik5pXDUcQCU7p7nVjBVXhzJluJGJwJFE4N
/R+D6saecv3dUBm4Q6LtX4dW1uCsDoKfM526IfPa6m0XLO+DjGE0MEwOhUMynpHvdJFsG7TUfTO9
UXZQH9+rXeeMtf++zgXMGIhtyw46OS4o2qqf3GqGD8vvPR6BDOMfJIC3rHr2nzNQhiHjbBj8cMHP
xBOOhN1TltWtL7uEmUPeQ7ICUqu7iYjSdNFwE7ywEQ3cJSuUjsCd+wx5eMvPxcZbDzlYOaTnvuN/
akRkgfRLjrwjslL+nca4RuSHSO58DJa2yI05K3rmqyqz+/JyX8e7js0z7SrCLQx9HAjOHI9mbVJ7
hrtRA9JJPHYGLgpZ5oDiyg5gjNsLckNnUoqi1VFH88eOSt41fSSkOcje0qKQTDUt8YujpiQlUmZ2
SKiKjzNza8K/5p4HcU00iz1jsp7q7sOfOJkU1FEP0OI0kkuDfEgGJ4XRUWaoeB+S8t9VG5u76aHV
RSMxv0mibawU3jdpw2J9qvR3fvj5+asR6veK/yZtBfGUm0oBI1gLleegQmOfYZbL+qbOpwMmFKbS
JKdR8TCILrmNwtzJWeYmezPU3waW7YHriW53pvvyN7BcHpmf0kPDSdAMEAjfY3VHWIqyQBDr3OU7
k91SUFOAloUD7+aZOCHO16Dpv2hlonETakaQ7yH1tJL85fkH0aIjlIfPtQ6YvJTPQ9Q1QB3mRPaz
XgcOwmNXBLq34Q/99crgky2PsjLzJtZlFl3c7y7/le4eqxexIxoWrexhVRS0RJhJkbZRJwPYApbz
R0yCAlFJh0uBKWlq7ThD2EsbnZ52a0vyCahMBSvzUMljQ7TSoYyJIkbY5t7CxmpwmZ6uES3HC/mS
X/pIC94jw47IDilyGrnZBhxYggbCPvpukymxzQiiIxuM13xTRVzrMTtwEg34h6ZefjsYBfvBNaii
ZuYn6CyAtUFY6PdhJqSNCA1RaPn9LJD87wGSX3MmhELNrSPUMJkDydCTW2k32C2PsCR4o5k81WYU
8nrYbchwj+Aw05xrKqQAaaAcKVuZRUpnwFmqP1uE3AoSc61b+u/DkN7cg5H6ofq9AB5KFxYPhz0h
+N93/9fOl1iJ0XlZhEc+MNVmSFAh61DtVjctIQc9moBr3Ff5MqCHsvqEnPch7forQv663D4mEif7
oW4yLApw/CTSeqmjmSnOIdf4+S8jt6M3/t57xJxmZAOkkF4Zih/U5iNFjgYojxfNGQ4KLIGMtp/b
9urLH4f0DhViAE6MiGKgZ+o4XvsQO4z+813+VWR9VsjLFEuh+wBi0TIVCB21b7fHcz93Sa4QQdr+
5r1jFN1/hS6VRB3dl/nR43x07bQP3op2yuhgn72E3ml+GuoTumJe/AGCSAHIkbWCctyNgaken2g+
V8gJJBD85lXEw3I71Jss1lJVSNFKHHeAjPhJWd5uqgPhwTF+62c5G6bDDDUOmwfnGrIjdZyljP2K
bFkRHWoPv+WU8GCLeLlLaK4g+GK3pxlOJlW7Hqeyxf7CRlavnKLt1OhoHl42RP9L5ZBnP5reLsEZ
MrH9PV68j91HWXwff168HxYWxm0FM6CqVHUPBxs0iPIZ5bbDZ/Z6Mr+6gzTAIOf7H3DRWk5pRz3S
ucJnMgMyqpaxONT4tZyD7CxeSoMg4/wM4sXhVVoqZBJofbMcmkxuVO0Yp5g9ha4PNVqNqho6O+xc
/rc6BoQsLhlJcQmow9a6QELlLG6DQ1PFXLuje2vGAkE/Ek5T1HPqsLcmhjjqABypeCCte6AR5QYk
W5b/GGoaOfXHIZNUWubRBiQqudaHpl/MRT06BGCCiuQOtUyBp4rEOSX8AfAIIS7juOY1g61AEOv2
WjUzDiFfGUnOPw9NHOERvv+RwMOvjx5ial0RdBO9U3+IjzS0L7M7bJsKb+aL6vEu+ma8sR5kxmhb
fGI8whSrucZam2lLRbpLvtlb69qNVzEaP99/bxEvm8ucLjNCy8Sg43gvHoNjbWIZLl/WzBKWJarW
6RKYw8AQXhUAWTQsRi5bwcR974tNwKly88TneyMXpr3ufjSZtuptY48nrys4zx997cSyLCxUuHLG
CYSiVFXja1r3erapoNSNfqJX4+SGOqBK8A9GDagII4Jvgox0suxNqH5ZSzhB/lysMZJtpIczMFlL
kZCJ8gImYMdKlXXTw7bXLRPqLcE3EU2Svt8VF84VfDSYo+qd+FS0aMZvYcnGaOL6uEyRuuWRJIs/
WaQZcbPb/nnOIhQpSUyyY2f9NRTAFpUeCZ3XAfsXtphGAb65jqjCaZurgsFQj9gGlytQ/UMMPP/y
AfqHPc2ImdhS6P+SFE4M46fxmmENIbGfYATFLrnibHiyl+JhyDCDcPKjas/jk5qmjYt707lc8sU+
0r+vm/w3hc6KM7eNdCTv3chdUvp5+i14c61fpBxdWyhDYr7m9wRzs6sxzprZHkwFNqdL6DjYh21h
OTDtiQQGp5Z4Sx7tsMD00K16mUxe7ejALjtYi1a2hl0ldlLtgBtnk9gPryPbQhCIiTV8S0dr7fa3
8Iytzc6U24bdKTwKKOcDe87wwV1YTytQENjryRlrIJ3BTa53avkfOSQHwD/zbve1dpkX8w+Zja+I
23k9c3oFLpgp27JZiCErU4Jifu0gCiJhjls9FFc8/N30qveQxqG6ftfxDRx/hnwF3A/hwVseHCGf
uNyJf3kLzNTRWX207Rd/Mezde7g/vyecHXv5BHaGUtKllQrDJnVktlX/H7tXCSy+R2FrkLhA/mOl
+Jf3ToM5U5aOZNspogfhq4ssKQdd5ok2MlW1H8c8qdO/9tU2Tpc9lgkDqejU8vzHLnHavrBlygb5
yWvmmc8YreY/0QsUfhUwihHrvaUHglfuJ21PwJnd3FbUECoaYfaq2YmoGQkN3WGPnzs1nYvDq5R7
YuQF4MuFLVtAzQTljIwmyx5fwHfwLU2JLq7KAqmNKN0VX2+FCHJK3jJRqEvktQ8zPJJIX7S6gGXF
1FiM07XrDDFsS+MhIgMpc217KajZ3vpkE/GoQyG3qr4FTpT7Yrp/cJ939d5teZPJa1j1GADz6YgX
AVpBMpinYnFPDeFr08tLr+06ryGsfW4LB2b2urW7DWVrUetEoUvPIvapCgePS3rzEdN8GpvJ/cYD
U5XECSmaxk4z+I+6VVJmjEl6/79jhKwxKFCdV1rT7I98QxuJGKKXT+V35JVx1jMAL14/JugslOhU
blcfLNA+FIwScVbavQrcwGgV71tT0tKo5BdjKm5QkH+TQ7KevlY6UelFLB9Zrv39ZmppCAvPXY5Q
xzkc+d30SDMDSzZVB/fUQshNSaZTtmMw8vUR1M8opRdRm+mpmKVnqUSO0ok20QKkPie7Q8EaeCww
eAgqxuQWOxrrMnMYnKrKZmtijyGmypmmU7ihLnyuJtlk9Pq/2Qb1Bct9iT5UoixlAS7L72nrZAnK
/qcfsJu5AjNCaFxaTZjgwHsX1GoSPKDlglyCJHfqh7wmZBk9k7XMwr+gypmBtT+YoFSZhvMPcmfa
ZBi5ndRqCmdIpna/gQN3k97UoFdtLKYWXq6nxgZT5JxzUQWMnTCo2jrg1FK6OjTqqHYsxcwbtH21
QdOSDdO+5D4L5HqwVdqLQv5S9Pm/2kpuYTBrTvOp9PUsxbROLxn+h0iMtWiK3flv7TOoRFidG+of
to+qYIx3eTx0UBQdC0kVqYIht2BET5oGvvwS7vO0gW3ZywNDvVU9VAHra0SY7MKM/fGJ/6tICXVM
dp8JVPuhp3xDQZQA/7G8rdXFo6tHVjgxasoAek754D5VNjEXA2eDEyXlDdAVQmsp8GeDFwMtuQNo
V/yNFE9cF+0fv4QZ3R9E2NRlzefwmXYsrE1NlyciGIk1nVzK1MDAjRIxTUtQEtKSizpxwTctU6Rd
PwmF7kuUm3zpF9bkKP/p33LKfLYx2ZPzeXSCOGw4FnhEtxZi6leTXmicsnHW+2m5C/+9S56f+pVS
TZzMyVtJhgAh0T6j/VgBG4PIWKRa4MzUNuCdPM8iBv1587qos+hgjfdO5cHiVlAEcoe0Ccb+2RRK
kwASLzVwhtBG3twttGIWnZ8Q5dRaZ//XhjIZwdGt24QGDGeXGoslcrb+B4zFxhQhRVolWzWBI1cS
Oc8IZvJcWgBs9tHSsEbr23GCKYMNYTZAvu78Uoj2DgOUPQ2I3po4XirbflNm0nkCfGRDZZ+Tl8Ue
XXJlUeOBE5bH/pPFmqUYGGtDmaCXgK/v+0qiwu03jJlvH9PWpwGxfqgKvZf6kjDMPCW0CgFiqwFI
I7M+EDFiMgGlQsbgthAPdr8Do7S+xHzLpRzIs6cof224q4KDBDZ8USLD1Id2Sd2Aoh252mcQKovw
4MOTH38VhT+skIzeEEn19mIJsZfHU9Z53RXpdjNzAnY8J+7oR2CogEoPj4GVTJqE4o32qJ9FvO3k
T+gShCpvZm5b4mG6s027gOht8zEQ+ax+4EO5vOuk6RLIPDDyQSLKpJQGSy/rODcqzgmyRj4BpaIz
1cik5C/zO/jEzCOsd0IOw1k52g9MywhfAXlVYE+f7iRJNuV/kYKkC69Sk2VmQFalDBKoA4JJYBe5
KuesmWxiknGo2TQirfakqUOP+uyKFahz3daOH2VHDN+zXmdXqZqnET3nngga+LF9JGshdEFmnB1i
PH61UJWYumOlWmvVw1JszffWjTQrC+6afGws50KeWtBMhVJ42nv5PXPHGf7fg6d0BRIysym2I28g
D/rdseESpwB05c4+LC46IohimEqjn1yZONtfbkZrddyePh7Ki+ZPvy/aXnLYf1puYNb8kg8owhf6
k0UxDNvK8/SiaJ3avm1CbixWTrShnWYufGMk+GGESWejadQ8PrSLZd6OE6jXDhhCCmVOQxSvbEAl
/UeHNjS9WR/big4S5nA8jbXqcjY7PAYbUKtWAHqUFS8lfozkDGg21Q3/hurBM/pKVXxNuJaMUUuv
U2GPAxUj9itzrQxRMdSqzDKScra6IBcUA7hNuXSKPLP4eBc8qFoWPbL6GddurKl7A7oXWNQ2dX+7
wNFe8iUPL2FcsDfa5XH1hvMlczS9KSCnB3nNCyyLXvt7cuB66EhUSzGK+M62tkOKrSD5X+eQnQJA
vy50YdxFGy9vNEhFveWkhtm1MWpzc75pqb+gggv3H++BeRDpR75r8B6ZtP1wYqX+6sRpgaut0Otr
LWvKLVq1Rj6bcP779Sm4dwitjf/Gzr62vcqfy10vG5EvfhLfSdI1avowU7jdhLH8HHGT2qmch4j5
du68+//Q5z4W4Lh/J8d/QegGNuw9ej0xDAEBy/qP/QIW1cfGLekGA5hOo9WbmMphEZUvzA/iWYQZ
gzM6vi/S+ot9kJhsZDgAZ1nBL7O3tpTrnsnNEuZ1g5WJeQVvJNAUukFrGr2zK16VtHMivH4QvvD3
I7stUggAVU0mjbcDyupprxW3+Q6l3b4H9/b3vhvtdrVg2hFtRRfdV0Z90nIbMb0/6YFwyg58QGzQ
GnddZn0lbFW7p//PVVhyKDc0a2K0noxPjDpEMeHmIdJf3PqZWB7oYPrxdqmZuUBFYhxWOCuk5qeU
elKijw5GQCcl+Om5HEgfHO0+XY1tSQCRDKR/YygSOU4hwLvjKVd5P+SI/npAkcBk50s8EmbtOCfa
6uXtaAQyzICbGNjWWXZ+YMOqIRtzBAmMehsp6fXuIbZI6tscJgt/T2sI/izmvMbZhGEd9EfuJSv3
EBLfcTdNyRA0BrkxP+Ntk2XJc6dmI34Fk11TnO4fBqje5Meb7Nit/ruz5NzftNq8GHzmFeomJkS0
pydiPaMBlcSecXs5ILOkyYzl7TXa8ZjICY50FjhX+iCCqsWmxL6rI0P0mTIK7fA+bvCRcrEUSP2Y
vEd1XX9YS+72s44/zzsvoO0z1lKFyYU9UhjtlbwtXCx4Hris/LKCEXcM8nyXi0WMt5hsvKpeYA2S
1ft1yBg3+JvLAlAfllz12YdHeCl8M0eMpzRTcDtIrEtSNiKev/+zGCtomQ1o6ctE3u/zOS+17igb
Wm3gj2cAMNaINbAEAW61BOqMW6gY6h9EoyKj4mIkktI/9TLPOxQrTls1rzCdpcZ6k8nE3s6BCAFx
RzGb5KmscETuQWKuLHKPn6m9fdtp/4j8HJVfq4DobuznsBJGWMOxJN5OwqA3w2FUmaMQfZUBVmR6
2mqXI8FKJnyHKklW6UlODT7O4Kiq40MI4GRxD3AxbCwSWggWcqBTZlDcxD0136RNp6uVCKKPPP7u
Fwh61Zawzd0gO8dT8mHs8q3L12Hc/QPZlr17EvwDvYwbS3Ugz8fvi7+Yd3mLdBH+YDstk5ACiQog
DZiIDjjyRX3JvFUtYZh7ACa1/25+6TA3fndP1O2Ro+MQGJfcV96GRccLj6839KO57XjJtBqeeOY0
VKU1Rg3lT09eUe50EFDf8/ykLTTlOe/pBPdn3vq4OVDwFCIVXuxxeGiKMZJKgRFG5UXr3lxg4Tyo
+yoqc2Ckk/Rp3yL9iwKyrKQ+t6R8oGKoR3RxevF9CkkL+yT8jkNSIfjKgDfVkV9kXlBYHzuut9r1
oeHLV2lUufz5SAOWd+oL1bqu0qiEAHrqqNXF0dyn7s3+xs2Q9gIcZr/AbCdJEINqbQCoqRJNV4Kc
Kjvj3xN51FUAkKsu42jEh3gmDXvXZ//yXsCxhevx4pKujhTatE5nqEd/02JTm7HhE5ZRFA8f6Wvc
AQ/glBrUZ14tdZfw2+Fzvvw1GB/DD825Psc4se8N9vPfsOh/rtXTdf/0syfFlky259EA2aWeci5E
jAi4QSm/ASuW91P49WOYADwOfO8l/6/adra4l2QzHG2FvrImZ68AUgjwdqjfxjc6nuA4A6K9/sbJ
6RGihDclmxw+LRo/S3+uiCkuPvBFqyPCy03MB2o9Qtt2lCU5/Vq92pRp3QoFHTQu4WweJ6HcpbIU
QqTBnxXL4GXKE5VD05Xo70jQHVdwnQ7wfDN3raP36UWiSsLvtuu1+Oz7txuTbxrebzjgeG+c6s8b
AkG1jx4ymyxct4nH1j33t6x0KYabRevuOWa8TrDwwtwLP9gXNrrZMHjDT9MbgDrd+3/1XQY6rd7y
fTLD7Zbk3DBU9OR4R7Qlg5q7VJeH8BxOMNuHi8jZ0Oz0itLYw1ihb43m2gO50s1oFGxhDbPuVaUk
9t4Ah32Gkq5SdSteIOsl4FLaY4XVAQe4NOYFEeo1mEXIKQrcxu6X6c5dmfRKZOx9jUrybz14oL3f
7bwpWlo8cONXJoCuCTBR5TqlX1FSKKwhFleEB1QQfW218FMB6jXGW6tUvK/dPtGHiJziv/QTl4eC
YdEtP61dQnseL0tz6/n0GXs1KovsKNVMomwhLvGoDcy5Er71Gss7Qo6gt6deqaU4NkwHkZ5p8pqB
38jVnmIKGJSCONpZJYoIvaFhIxBqEWZqs31kUK0fZUG8wEqox3jOmmKE4oy/zuks1YBSFrlEFXqJ
RzEiKdh8ZK3TyTC1paAHFysSSk5PKDfM/dUcGgv4tkVfcr1d3GLhAr8kjqYlYY1TqHDNlFuf1hj3
THitJ5V2oLQHqkAuuDEgYqSLdPVk2QeWdp/KsZlEVdxYP+ntoq0s8OH801aDWIkZxbxJWTrTagP3
GI2OGqgoO1nFPxbQb1bnJIpWV4W4nGBFsfztKGObOSuo7fqUB3HR+usgwuxmh1KGUwcSnhTgy9y9
aQNvPAFUV6NuSi/FxSasN8gpyjxWIYyG6s12FpER8ckRSzqfhuCrgFTuH6cRNfBJ64z0ypJJkhw+
mKlNezoGPy1H8XHXmNmxL3uo0kBJ+rlKlkzkftwVZoLtVqHyGt4BYBXf2BSluokdNbikdKFr8EaM
pFqwZDTVziMTUI8Qj8/NgQ2C4iYg87kCZIgOq4Hcu5sgaNT2dZYw8qSqH3gjSIioQJx1/cBo6rXF
rYkTce2+KQ4aeo6Xs3jZGAviknnlO0Kkl0np/cCfqoJfk0mCPqWhPCEXoQeQLr4aPvr1LtmTlLU7
S9QN9oBZb62jlgv9fL7m/pmCl55F0YWKQKsIvWTjW3IWpEYD/cZJGmqhVhNN+hnqEQB+XzFWcneS
NStwhJdc5njAUO7YsG4BTxSFz8T3B9vdRz568JMG+yTU3oQw1dUdMKB9ZqbphyWz0XRSVzIE2iKt
dki+GuPNMYHMM01jF9oM/YLG/vQrvbGbxPX7twTxen21+jYEsGxco8+a77Jr0nWM9Dampuf8MXKN
0omk+AsjF4tY6xJZsrK+OrTCWcgdcF7RPMTee5VU3cB7sQiDLJSGgHlhGKp9PPCBrQhnxu3DCREP
9gfN0aqccVCLnzV29Va4vlsB3kwwbSaPPY1/zYuItMy2Jy9UKKlbuV5APZRlbBZAzVU3BrBvZ+wo
17YVjAvcvMyzwLJnESsSgEg/ShVBlYzaiRfmjNmm+omHbnt/woKCOE9j2Ws/PHsywWrR+xCoAs/x
py1wzC0Ukqziph42gb/z2yapCOeirjcBjkvzvBJ9ANDQ4+9TkRrh63hJxZaAN618D0AFyZA/2zXK
B50k7w3xQqhABx53W4HeJZA8zoMa+jNcvfXgoulAkrCLRr6lNisk/+T55CkKwZlp09eEuKjPSeBm
g/bVRIV2cFlMK171RKNk0C0ZY5vEHMWG+yaHx63ypFLVBB/GK+6qmWi7rI6Sy9QJd9LkO4JYhrRk
XSe5tY8XRdd2xCWH/bbx3RXWG+W3ERaH9WSxSFy7fr4weKhSgpPIuVxH0Os48b+XZ3foHnWLCtav
z3npxPKPQPklN0ENl/68BgOQclU2ABKUgCS+7hJa53+zTFr5SbKm8rtncrn1IBJham2oK4iN5afR
y/h18j+vy9M6Y6cc55fd8mWe1p75MtKFXCx1veEfDBUAEdEXU9vuoSLdKD65gAWiFqf6k3+PlmiZ
OkVSPyxYW4PMjhdmF+MFx50jgaD2J8YXfY+1X16Khq6pUlSh9pEDVHWH0/Evpdc1A3eNFIzNrNnZ
f/3KR4Xuc3SY1hnknM86mZzsdmc0E57G3gnqoll0DZYS+qZCo1dm/0zT4cdzFxPcTShUY2NONh+W
q13z43VGo0EcsLcl87/cxZjWDb6fjBWLbdvV8IxdkPTCQ2kIzyVYKgMubSOhjl3oVfVIPZHjfXrR
IWOXZeoC8f8zsmffbAv9OCWY2WjgE64jXXO4EWOO+HC5d3GFY9Pa3jIxgCRS/gJZVVzfBnOns16m
UA2sd+7w6FYnpP27pl/wdfpmC/dgDuO/QMStFb45E8P5yax3C46MOVQXbfsn7KEe/9gzwzFtRiDF
K3offNTwFh36iwU7Rndah+olwyewpj5F5dMQpZBnWVq1e0InRW2aHXcMmZHc0PTWzp2X7m3wjLwl
MHE9Q5Ft1gprQhMlxFjGoIP4TVG9sISe/TRD3aSmb+BO0msU7JkdIjDwOvSp6QKz4z7BY0FTjEpJ
gl8iB6p/ZJvxmyZw+vyMvAJmr27MNdWCJQ8KUhPzgc0UdsBFX6E8opwQSuDdNOLw1YexA3byKKrA
HmRxm+cDGI6+sMNktbi77zq6n8Z7D/EMdxip28VqewlIiE9tni7LXudPfa8NAk+B9DN6qt5NfPJT
g/7JDe4OXvbTx33kvH+m3gntK2lBOvrzPXXIp2SgrlMXVWmIFSY0qf98J7soHSbEkunmM4urKhO6
TWEjg/buGc7MthVUNksbGxjgkC+kTBne9bzlAiNPwTtpFbjcuhYhhJWfNzngEkJ/jKf574DcHZ3M
dCr0OLMLLElcylAckzVFgJajVQ4XXiQfhpO+6eKWpnkHk8mhKymx0O7cnKpxdWaNk1dVK9U9O4GF
fIrzCVGgFmVkZEFVYyV8y9gJDikeAe7QZtFA9FrHHECic9A3VdbWSChR/jvurCoZDqAS34XR+MPq
Fpp+1eXkvUToaWR/KK6GMNUbpya0LW0svJJhfVDO7e9c+YvdgLRCTSeIdoU1raWXrXNB26IpN+Qx
4g52IMZuwsb8QP8DuK4rPh1pH1TVtqJqFOjwICNBcvnA/mMawE4NdSDw0gS1RtpztgRSoC2xcVfd
MDb+EX0tAbFGEP6K+JSJjNRbaAk1TRyH9ofgs06njRh7N1nwoX1GJ6T3OYa0EuuUKagpjJlFyUc0
DLh3ygZpWa+8qxZqnDsKo7aImugRNTIVzQxxWdBzK2hQDsqlKyfj9tQlPZpCOltEugNp4AQo/Bn/
xib13qM+Xx2JZmg94Rqsima03jij1kYVGrmAVAKRAkyr/SaslyshQAtuvqsMPLzVuINC6sNfYMFH
1Zo1+V5bNe+njWx/RXp+Kh3GwFwd4VWha7EDUrSYbgIICGrUYmTmjZszLaNVdTXIG/yYiTHKK2w2
Wn2jiG+HdRblAUbEdg0DNEMggE18UL7l3npeVGLtXVxjO1j1CUgV9q7K5iy9WoutEnzFdPGEqur9
V5GuBoXwn6u03ydkNoBI+ZEf3c1+hC84T82MFvvLwVj8KOYsHZH8lgk/44CWbuIejoP85C5Nuwvx
h7RnnplmSsOKheRn6kJaDSeb2jOnIEr6yogWlcOj+Izjx6eglpzlcruS1SC4hh1IR0aVinQUzL2H
zCU60URiGem9x9sJgfBHhKZQsMQBYHObGn7MWFQrluiM12/c4TH+WpaRdpMhcjzRBC1iUehPixj3
aSyay2tLgohUJuGm1R7MSyWq8nbZRyv1eSTAWXpmui9BPeO8lcHmtoHq2snTRkWO4G1FHLQwjTGZ
inn8Yh3ZspLL9zQXUJ/tdvk9c5V0hF0IkoGHc1YDPVXaTHkzDq8CPL0hCFxdPzmdDaiBBFzlDL63
wAKSIj6pT4HfSBLnzctpvywCy0JzQ2ldAfC2pPFnDUi+S9ldcr4YFn+VwIkAec4WGAZNJlHNH0oR
94IgwuU+0omgzRS7u3e5tx8Nt4KpdoacrYqYo3t6IDt+rKX19m+rt9edAjAxy4OpXZwSZrxFanGW
C17XZWOoYItDCJpyIjn5r67y4yamTSTBCHHSTVjy4jDBDbKFBIABG3oCdBOUkPtRmkQoTDRvd219
FfXFlCj4qUAEQr2p0TR6YtrIV/3KGk2Bb0YPWhHMNQvMApdubOSZM7dvoCKfI1Bl+UUqNpRGXmxF
pTUhIc7H2jngQPkcmYU9QP2hw8s9NYZgGjb+8WiK5qONO9nOqreH6akvHRJKlEX6dCS/UxW5+fjQ
ykGH4w0FJI/W+sYgOexPSnxiFvXKjyNQwuhst5XHFMoz5ISFEKBuYd4vz6zilbFOTcXolF3kHgbM
IitN02anwY+EuEeW9qyak6gsPdT4RyHS7hwhL3G/21aZgyzyV6EZaXlEH4fPWmqbc4RaAATUxjBb
kPDcpgYeDp+ocqqR8UW5LMI1vGMS5XUT1vEq2MIzE2nue7LS0TLI1DKK0gKhh9y4IRQiYa67j3eG
VbOV+gyfH2RE33KVuJEnkHjLbH7r+O5CcwDnhU7fTVo/ZnXq7EBfHqgf/d/GDcIxV+7f6Ptn1/5n
0iMOcXg92ocFWw0pJAVe/6EjR1YGDFdDPI1EP93JPHgKlV1luXvny7MbmK7zjO+zFjdmQv4EkF2k
upBvFsvP0JZSrimCpD8Bui4ETi380k7bJO41+5UlmSF8TH4/2L+6v/iUUoVv1FKEROrQFsAYrNkN
4riDCypZO2xrO6ek+2jBkXhI22Fs+GpdTdCYDFHEBuT0OZYh/6772iNxbDlKOokTPuRUyKdkYnMO
eywUivmc8jbvBaOaIIEzqYWeaItByFC06bzrRDgzX/MHWZMKIWN+9+6hXU7JZqArVBww7sS7UFoz
8r0X5HAtcXhp8pZR306a3lL2NT+hQhrL5djHyh00oPNEz5g463P9qpkMUHMaSbvhO5FrhBkY88KJ
H0BfJ9lblG6JM7l8ML2noDInfbElkpyHq+mO7L/RoBZjgFJsiO0Gw/Z0uTjNz6LrwCJSIE90wNBn
p2yj803g6Sch713O/Iuc/lHRUKMrTjfrnz13/C5vrQH6imY2PMH3CbqoQ9dflC0ay7tQZWwemqND
xmb/1PvVKgoV1X+y5ZNS7pQ7OIUZEmJKNam8vd4ecaBbqWkN9UzlaSsy8CwXblCiEXzjz0YxmWzY
//LBHpwAa7nZRv79NWfConYV58BCrU9byjMsXn0Vi0Z4LIStdNkEsFB+eQzaOoEYdly3RasBdSui
xsRzi6Xg1p7xAvH2e+MNZ2FvZPpRNu38k001dRjExJ1BZyue7o+Gz7YQNm3G262NbxQ3qgBltkBk
0KgjnvE+mnXYkOtDr6OBe8krvi1AgL7rsbthdLvQNcngxPD756g4dzYUy1oQ0VvbZDHpATbGyhfP
OKPc4krYIs67DnDaM4mqLqrqd5Zvt/FsMqvH2rjMSCftLtS/cacde09GKYgMHqhtvVBtywyvC0XT
GrUHf5BkVuUkbsVDCYvOnCjf/sFzyGf/mqcq1WL0GMQeDTVm8dylaU5ICnB1OpOijfHUB/PMU1Uz
JRV/8fvcgDO6MzabKYQFE9U12sBnd/joC3OjEosDoz+TZChKc9ZUmv3S5Fhw9Z6hp1QHBT6jL0lD
nEckxZpg2LR2X1XuoAqO64wihqCXyzU+fyYbeqdpyvTPuNLMZWaagRqC/0E28e4DLNSBHJMGIfZ3
ecaONRqMRyMM2gOytPbWjWKWrVEfoHDJgQP8caagvix1936fK3F83BmSOHCTHs/iHtWLE8maK+5e
LuCLl7L3uWFfmUTjFIT4ACR0nk7fql4x6tKeeH8YdRH5XAc5BBUs/ahmSWpZw1Rs3xQckKax7CMS
6NTmNYZcQK99xnLc7LzYmqsxmz32JKCZnF06rdzdWtGIioq78buttpoBk1+eoZrx21wPz0Wzf+tj
MEDqAJc6XWiqD7G+FYH64mHk+tpnFpZynERJEneSwdPJ82polaLjiItz6bk5AH3OSIemCKOhSTQF
92hDgd/GOlSH605BWd8K/LVGOAgkdzBT+fruyo15WcqCYB5pMxr6PSAdQ7OxX+O7a1YTVCcHd0rH
hUISooFbUMQ0a+SP15l0I+cUBW9CEvj8LPoWCLTtI5O67o0ShUlr4qdazbSiU4dNvRbuW9EW5vKZ
wHrGG/xoZxXcbxgbv/a5pV0UqtbXHF44D+sGVO3N6n28Ng/VtS9BT+5cmkGTLG3Y4RjeXjAH4Xja
8YemXTBxc5goNHPTrPUNFxAArYOlBrJ0z0heMDFkw1k4+mFo6yv4OA53uysepqbJrAUtuAhKeeCV
IQGHSISEaAJ8mk83SRcjysSYBcWIIHN16qcd7mkzyQ9qj37ssmcxccOkdX0vhlErAb8pYQPZKSyw
FAhN4EZXkqoIp0QJ9YAq1YtuzcfB5j/rJcfAIVyTtvaBawakASvqXpx9/w1ett3FF+csI5XT4KNz
Xqij4bMNcXYOC6HUHaWN69kN7twSII2u7289Ea+PY/EoreEcoEJixX3Fr6SdHD9pjKQ25weoBACJ
5pNAstJr8UeM7M5gGopWxjmyhT1aEikK5d7Ur04aCnh4g4ENTLY5Zq7AYzfVznDruWzsK5kEGUBT
NzVeNpIHAKN9N956aZE3oEdm2J2nNDksYSWBms+wn2A/9jk0K+2r6Z4LKgfqzG9yA945iN22t++t
Jo3f2Evnv2AGdMd6KyDzvFZQITDk9zC0k1oDsUWyliiytJC0rO3wd6dyupASAgeqPGgTL3u9Z8OV
EtBOXojBcUEIYd4wRrU7dTrfafstohWJRXx3XVjtUC4njkJReoUF6F+PQaNfnL2p3QxXNk+kTZch
LK+ajyYr/BgSWKFxXhpQWnwE4EwG9ctXTr47OlrKtzuB8Hhizo3QMZ5zOQfnH8yiRByR7nssPxL+
ByihTBPPiQeB0XdIrNYNMoJoLZF76DFvBHNBV8ngMq7Y1OV+zfOZg5PYvOITGaaB4VddH7wBjDv8
4RwkDijORp6cdGfgYcdOmMyIdFNsWzE9oSf+WoLqZ9Tr+McEbePELH02ssTsv5bF0SQynqZnLKH4
Tsj0gRmWl3zwwhJEiitfYFl61S0CyOux3aVzTn6iBIS7EIq8KHDEsOyEs07LMlRJcjviqt4v3PRR
fpLMUX3aX9P36mH0+CGmpP7/VfTKtM1KTt7uLmS/yQ8dM+XgZbrC/bDX5Jq5uvlp35zjTOf8pKnj
cbuESD68EYuoo5+2fSMd+0bOvXEzF178qQ/92mcvuxMmCN5BWxRTSdao4KpppUl9EgX0VBPgCsJd
8UuQgLWlvmNFyFq0WkE+jpIOu8N5ahwAN/tttKDK9tT1GgdnVDjxTh4dUebQMiTLpRvD6DhnugBq
516xrbQ1jqPmUB3bMaz2WR4QkVs/kJtHR1SmT3H1rOpQdr2npgALymg8LSClo4rIGRdH54v5MLeq
sGXaZFQL3Qu86bmagQr7NLJOXMrvz9d04SD2d98gAu9ASl2snP0NsHG80BwevWENYzgDwUx3AbH0
F4vCE0OJyV0ptjMd547PF2Sk/C1VSp8HWzIk2pwwQolCugT+DVtmo6ykRTX8CoQrbCx6sxOHPJXO
a4zkQhBMIGPpZ19obFmadpdQnCWYprCrIyr0NzdMXJN0STO4APgYKj7FXiatDzYVfandw+jhoD/f
2nWHbmIRKWHEYcPvqWCiBfAVXy+LpcmwNcQOLOKDmB3B9otKRDU3R0RlSioTIjXjk4zkfZ6cQd84
Wl1WpSw6lQj7jMUQfYDxEZ5pbY8YkeEkTq2SeUSUhRSw9jvKTrbUi8koArAHnGHVSrjM0NicDGFd
R0Jt3ho3MrPGHLEKSiC63X4EvC+rLWTHn4hfJaJH2sd/MDaX45K9IUzUspsSRBo9Ag/Eol8ydvp9
3NJrdeGktD4h3pchg938dYc6YWx5UYTOUSQRXdBkU83aVkcYTm65FYxe4HPShWKg1w2B0HlCwcz3
tzJ3dt+5WYz8bJdgraS1wp/USOH6L6rZISmd5RKWzDfMqbSJnDMJRql5uOgRpDf9az/x79AXRgNP
OYPjjVzs+4S7kBGckva8UpWUlrF1SFVQu0BkC8w4fWPmf6OjXFMZIw9vB6C2o1j24RwVf8sdIsVv
Orq8KbX41pTK9f+3jpsHNeXte9i7948nNeQbJtIoaaRsX0oRG2MDld1wBwIiw9rdgSp/ViYjNG2n
zV2LstxUY7CFXExbLzHPcAwToOpwqPE+a57kvnD7k0GVwqDnaSfbjKoNs4nhr0hK0cfI3PCbU6UB
Ra7bTuCpgZGYfN36VBR1bryxA8HxdQM5XL8tRn/Poo2qMSzgJY/1xri2scHFAVPR0g4TMJvfcZyW
sq2Yr+fPEsyEIah4kFdLTcCpCOLZxxdqw2IspwlkfTHoIFmFw6wCRlQrR0UHLcsAO3PQlG+fGdkV
ct1cYGAuN0/L1wGP9cCGSi1jVH12jdGzc4xRQAF7FxMjE7vlWT0Biqyoj2WQn7xNg/YJ/fgRJhTE
1f2e3TTpJvId+Iqgbcx83tB1o8p82r41oE/h8ptlkLZ5CVFNIcJXBVNQ48ocNkMkoIdTqg+DUhKs
5G3h64qmcRy9s4xZZELLYdM3c2Jftjr8rxerZQsKt2nWEQnO56FraPJvTETAn/tjJucj/C9xPYLi
PLq45tAm/rl6UipHA12fZVyLjN0HyiflzPPsLJ88efUmxVKRHklqYt99rcT8hZbtbBvtS25IN86p
Fu/gXIbJ57/MSUPpS5y2r3cnCKfdss8siAo5GmHzOjwaWM089LMw5M9wId4IsCFXwOKEbHwmelSo
xOjnwMeshBR7L+Tg7RcRd1C8IjczwEFiSlVRpEdPo9pC9EzkVcY0OjsRLDkrCO2dE2P8vuTpjh8i
Icq9SoH8A87aPcY+bBVWfhHClyczqOPGa00lfewqUNN+jpRbRXMtkVDX6QrGUV/PnzBiLndC2GvO
oM/bDFSTju2WHlBM6RZBmO2h37me30X8303K2otHp8NlOrt1bmvWiAVE17QMdh3eVpupxRGWU1iQ
nSLuXvAmpjFPdWQkS6WsVB8oQTEo0BkorKlgxR2BlUKJ11h4umNbaEuf73KjKAhEeDbIp0q5Gjds
RfzYf4lIxwFshj/fopPiul4XfirjHrGiBGSlyvb+anQVfI1c/r8DDBWcuRAmNsJ3ac0LYasK/NbG
CpjRgtmQtKrGiGguUF/9LTfR/HcU6f1zLkO6scj1G9TCpKvVz+eFwIf4YpgdWwFJDGAVWZwNw2oe
/G3ue9dmpajesA48TDKdlK1jxkAmuWvcIsqxuJdzxNrZParmObGE6kblZk32eOPz2x4dCYm8cGwG
FtIhkpVM9xrDVfEoFsBMBVjMFoVEdmQxXYvt7pnTykAdJiSmIxChmk0z6IcylD4t7z1kIebz7EcG
O8X7OUbxeYkHMDGQoSjQdSGmHyZVnlIEpymQmRCJ/Y+i96OHCNK5qigOFEuBok6/adKAlpmskgSL
IUptE7oAooN3wvsH3w9c/MVmM3KWtvC7hGs/8j5zqDje7XwZ/PiRW28f4+gRZYRaUe4pZSa3ADbg
JE9pNzJ+Sx1Py5wNLksKXcG7kJCij+wKGF2lDFDl3K9rb8uz5l03khA2hx42nGd8ORNy5WQL0G6Y
nqIw1WNDTDpIH3pVGS/S7RkoU8gK/1wRRhHaJk8EtsD73GhRlNgzBCIN5KbD+RL4nYJmNcvLnc14
AIo/2+TJJ3ZBoD/Oa6A3SHuW61i9B1vMgdVjMN/TY8O9lDlQz3SVuSKWUZrPQm0+bOCEXdbgkU4M
1sVIqd7cFAgCZR7FX92OHXzHf9hSB9cS2KdUKVX5ntthZJKY3/Lk/wXSinnW8ykw+QATss+BARbH
qLQd1E/LMa1D1zCvzDxChDP7BZe44mGWqC8R8xUzFMUUH9nt3UbiwN83wOtzY959wD8d39evhcnX
QL55WPtds1AGjw+hCA1IarXEWuX3aO/wUmCoSiBnxAi2Xpn3RWgP5LNLqdClV2fBvyRMrekYn2lJ
AhvgcdCPCudJYpa/qQ9AQlE6qjxX9mykX1KOm7Zo1bwRFZRBbH5cFmWe3VxSmMbZTwAr0PD9vuKk
b3OLrVjBjH+rM/CypNEJdMLXEEY6wdEAhWkCHFSLcu4vgCuoe0tuq+gHtv1wACV+5gT3Fu4Yjx98
DGydaY571hi1nfcHeyQUUAPKF5+YFNKd13gF6gbuJgf8OQDLCVhgqrWw6lH/Tt763Of0oZsSEgJ/
jBDVBKN4ZYkdyVRKGzL7VfHtCTrmtQBcz9OLzQ/dwqkWZGGUx8QtGLiVi0+xEiQj3jbMQ6Ir3mlJ
PVUnbDw32/9xgPGC2Myh/+77S92BqjfKKze9VDBbZ26zV1B34V6YNrCwGyty3GQW6JdfYD/n/hYX
mGu7OP1jtKg/XRG012TCgMeUGmjtJz4UsL3zm5AgHB9WskuahqeniPx+2jP8O++a/0HXyipqH9Ai
I/dGzbzZNKkPw40HXrIt3K/hJ2YgInTi6k2a7xBFm+MDZTtMk627+Zdb6rI4covkDR2YTZpArEsm
6Eazz4YUrn2+UFp/aBDJLmVdVuyHqiFOrMSVyYpzfF4iGgV6s3rkbJwJKc3mVmo0wRSZfMn8WtFQ
rEZMy9+EwI6ahVmMdfniqDg4/PPQEgw2mAjHmokaT78YkAqk5dtI7l+cSFc0cv58lVC9ugBJER52
azqoQmfAxkwImA07lr8qCExM6DmAKv5gbQeKqM8KTK/BhRcji02GjqY4JzOQyznQL1QVJ7RqAAuY
oTBc1omVCTUpz4KXfH1cbXTrROFLH4+2Xnbc2yA93OoE2YcvVYa/HC+j7eZSnliBun+WsN6c0cWT
ogLYcubcSv/KrMtGr9/wktW8D53NV2uuMUziOU+QvYcLbhJzeD3dk1v7QtlLkNl9wNxMZVLON3lZ
HIU0RHGZUKKAFwsD8rfOogjFmbYDTu95qznKAmwNwD2PahPRwLRjcYrRQQFLiABDBAilzwAdm3AW
a+LEGf2lcZqoqb7TKdk6kPrX+iCJ0NWtE5JCgK2q8pTMYEgUypcjweXdFDb2eS3VsisAGTm4RSrW
A0hWOGr9+7Ety4SrEbNzAk0cyI1wIyZO0ae7QsQltuQDbzryN/C1HOjEMz9919WMGjI0pXdGJK3l
6fBrtRWVf/JGJ4WxwOBDCH/FUST8PcWRLOZEr0puH9QCsF0A4sRCMeM6IXq3EYT4cO2ZEI5rWCEb
NsCqStm9cnlyabSamh0O3CNs2E3O3KhahQ/xlFK4bOeBdypvBrrDg4Y2fkj3xUWos2DWmL/VZLgs
agO9otoYlQXhJyC59cEqCtIHTAqqixYow9RE4t+pg0s+Y6Gbwy8gVfrG2iSnbkRwznAiAsD96j0f
UhlKdvJgijdGQTs+Vf85kMuJDB9/zyxufxFLy81+0cvaK+K9yM8ml2Tjm6z5X6ekPF/ST2FkNsjt
6si1LDrdSaNq5XqItTGBxlrxLB4QduMOcZ+XxgvSXZalbepaYc08wjeaXnjKq80d14KHF2KPol0O
8YKJhPsXUC/xDlwRPjw7Zi3mEBoe7OtXyn+qVQ1A0jqLJ7kdj1ab8k24DvsdTq9i4KFVPNIDehPg
S+3QtM6b2fIlUhXZZ8AmPQW2Wu1x+6cMx1J0m4IRaxnAxo/75cP9Wq9Gd3dbZwe+D/R32TqkEZeY
auJMe3UwA8Ibsu3bIYG51PhVaWIyAXN6Fu95pCcT31fXh+PDBGaVoecdgHFEf6rz+MZdNYxRZFpF
Uf5NOJop3ZwwY8oAR8S9PLJnjFUR8MiYMJjDx3XFVylGDUUdFbMCtvDfUh0B93wEkJTLcp00b8Kf
g6rBbZY56eVS4Lp5Rvk0TCLt/I6cjLfbrVyRjwPZRT+rMwLxvELIzHpNLqtebTmVekTVIk5VEypH
O+AGXA/iQreFv8Lo4uKBkfZHITG8CL4AE41Re0A2CTFg+cvjU2QMoiVf2W79NlVOT9fwhNFiv8KZ
z0UV6U3asGvQuqxzk7J3cskcQMaZXesvPnu/zCCmW5uRPYLdmy1s4iSE9zov94Z8owJ5+uFni6iZ
hAtXK/5rOXL/Rd7Xf3uBhyh4wHzJDTctBAh1ffIK8AYb7i4mBIrMNDoWmVLeH0QirMQyBDP43z9k
qGO9sWBRwRS9nOhbnCBfZLsQxxZDArwMEz45KIkk8jK7UVNKgKFfRO10elYvi/ZKy6dnh6xPIwP9
NDh+TblTtS7iJbqIQ6DxYlFo0tf8OOAxGHdKsq+CcO93azpnQ5yO1CeheyDcAwlN+lp6EiBvf89r
GHXNkRxY2nqwkK0sWeFjnm6Rp9mLBpUc7csvd5NTfOvw3wmcPi33Nctw4KlfRH0WNkBOhxy3infQ
qoc1zsLaGttfzTDZIx8s/JoEYk4lDFVU9jv7DpEgQix/J2CqhuduW8vwJQeODVjIYlKqkg2JRl+3
6UDJ7DAcmeLn3+uuXwO5BUR7xYqTpVpjoDgH+A+QAxZi/3pMlcm3hpsZqYNbAP2yVnpSLKN00YnE
OWiJ8lWoY3RTr9a2ZX3LWxga+0xzk7Thfn2PlzuM8i9gcLtC4Y5CXfwRe/+HIJYNsE2VrSXVO5YO
0FZgzjv6PdRj8SRh2oQXIoWeu/zdamD724754Qczh4wglY/d5t0UNOJYn/luoc2spqLtrIhE3+fx
II2SThU692kChP9uIEscvYYclinm4QTF8MZ6Dm2lpdLeV8GSsc0OvUGWSDH0/4H9TxMBgwDeI/4R
NuvVOrAI9TrBUVUCKuVPHuZ04P5jLK1TfmXo3GKhv0jAojtYzcBSOSzgawN/bf8qaZFEVFanSqMy
kNVpPv6XjnC961W42XkGuAqht7UCB6tfnaqjjJODBEt2m9tcrTm8IKRhwJUPiQ7urg6iLNn63tGb
82+rxlXAmZrbviqcge5WnUvK8s1HXA+cWVWliR0bNrKpqTpLiuWLLeTOK33WvPzR2fO+77BvnT20
hL183wSqv9GWzNhg6NM7it/T+blsHYQuzIWDypJZZpVf5dmujGmVYW3vI/KJcaNEeV8z85X0Qb1T
BnBz2iejHJgSRWiTUpv4jaJ/jJAINxZ3SLEvyR80ueE3q31vVOMfb8BnzG2KkQzAxED6CnQ+4/4O
gWCpTnbWXxjHAo1WW5MdNPIzBz2c3z3ksP1yE3cemyODuEq/YSTfGWmS5rtVCVkwDyCSmoJqX0F/
MusuXf0x9qhzohA1rQyo/A5iCA1ycPuX57asCH+3aNghWLBPbnU9FLVvq7WUdHZkpeFPOQWCVuIC
cg6xkVxWoC0Ap3l2H1T6X8BYVldOAON6+6dZfdaM5GNIBSaIhatAU4I4f67AGiJdvlAeSBTAu/dT
Bqn7BIr8cc+Wg7vt6Oa1clOmQ6biKC8/pd5WHcl0b9CBjRFMnm40oJuNpnjWUJi/UlbsfvZ6Mkf0
WfR6gBzgJaCHtV5ZXdRTpmKFI/ZKTPSFJnuHdRpnDNEc6rxreBEWibdS8wqUyz0M4MBUYP9V5mRT
M5UJSJNGKKTZHsr7iQTJSSZnVwWRBAB7V/Wf1Hl6/MGRedQiI8Ccu70Fuur/VL1eVITKPS2iWp2z
Ga9F8BSMxqyb8p25aEVSdhfbkGNeljOn1uRItEKdq8t5vQAUy9TjnOIOOXB/ppkelklG7vvpnzwy
arYKsByZu9o/JieQoq1fhPRyYLSTU4+P0jdY5XbxHLU+wLK2oqeQBa8ec3h1+ixSwefH76uvtzuH
P6ZFe8p0RVDaNNw5a0uC4J7TNEVvDpqGdm5pdw6m9k9zF/HAKhjw0eJ3SqRkYDe6W+3REO5vqE9t
CbUKVlymjAUAEpsVgj2pfibWhAkrGBooA39wJyyEJTIbDBzuowYxY9iGZifamdExkp6PLc64S5NW
0J8isNfrWdIcAsODiuCCUl5m6UbanKYYX2i3yQR4Pyy/aGnWh2XBcnWJ710p5fzwAZA0zLBF25Xi
k/5D78c5BLdFHXCH5d+sZFWa5wnzOfiTkRsfRYdyiWh/G9b7mE5AXvchiUHquDv/kJGY+THH8f+1
eN0ql5tt7uhuw4bsRuiG3aQr/Ue5Kh+RFLTyMv/vDsoEHB0PWn8ZlaYvvdmJWeoOD4wTO5kEnYE9
K21n+cuDt+sdL9axhQZAGyvERbnpHYCWINB3Z2uIOMd+9+5+Bm7PhlEgVPXr7VqyvgRa1BsNpg/a
juA+Z28wxnOyBZM9LTXsWJjZvvZjhPldWx2iwL2iVFwtqeilsrO3d31g3EXO1/1sQGBUoKKI1tsv
uFcLKgX85uY3ZiesYP72UwW+vbYSvqp+tXh50qEHGi7PgHt/oAXRzu8VWBC49eHOTGzAddKeiHWB
Wqz/G3rAorbYwTPtj2MJqXWQ3994iiHFP2lJK2RZWXrF1wVAzjKB+8q+gapLfsfkMUNnzORQfYmj
3mfow5/i/1o7NHqzQcJ2t8GqcAHkEsGYtpR3aKHLuurHnjF/amxHPZ7q22XXHBAJ6EdZuyR8QxB3
DtkGZZtbrShRcbdayKjmWQmCVjEcJxg57/fm5sKz7a0W07sufFPDlZUEh85TQQMws/EReeWU1AV9
R/++t8E45ua/ge7P+vc75O62E0mogqq/H0ywz5EymYI0CY0pHl+rukBOS8TLoyAJ3x5TPfANZUNS
TvbLs4oo4/dZ+jmv7/J41Qbyt0wiF8edzsT83gOedv4dI5v++o3FGk56SLg+SsAzpqzfnB1JCyOx
RaPRrDvpK8nXLG7OT2awxyRGu4iVM9nxTMc39de7FZpOxsJJQnDop0YGm/i3c+ufGJxC82whT501
VWDSSqgWA+eKEkcu2207iVQNlVvdpJ4l9rURrN62Bsox7pXkxVq6dcrbKG/tB+m5U3yhDEL0xtbt
eAb+hSyyuGrLstUeBSieFeSlFCHHu30OxyscDyYGvr4ThbOyOIF+C2LkHm2Rn3N06U6rx3QIdQAZ
40slPbDXJ+ITkdVBXUiaEEgQlblO5qMusCVrpvrOUa0i+1GPHBpZPGwRqao2hOKi3ZCH/MvMW1t6
OWCt+/kGliRdXLtOpsG3G6Ed+cJOvBN/o0bOcqwt4MnYxr9z7YxetOc5y7HHZM4ofsGcyZPSpt3T
oDQSflY4h/nn9U7yyZwRsh8N/pnhHQlKSErK6CYHBEK5/XsKCGB2j5iha2Ce6es2oJkYQisIuKnc
QjHTS+lbkW6a5BnEdBWd5hsBsVXf9UspKJUEkXlHWTxIeMxDp/IVIwWlgDj8PigEEP6W8IwgfJnS
TuKaShXGVMEkJnShsSqCp+srWc9Bf976CvELOpLp9loC0Uw7A9f70BgGtQt0JP9bMTW38rcikNbG
M1NYJZePW/akc10a0v7oJWTsomgiebNGwb7jZaWyMQjmlVTpzO8R3DX6z0y6/RICVEXn62dBSrsq
qc0oSN5Sguq60PDyPxkXhce7DpDPr8JyZlueZT6rasn/bkaLqAcRfuCqX4iMexmv0boKZ71e54BD
YeG9qMe2Tmqc2SCTDHQgGP9M8J+PrTtxkOJHSW5cxX267Sthc5Ch2bX8LyyinpZhZvINuDHw3Ls0
AHRHHryEGLGAXCLXwg7621chovuusqsJokMEASPcVkLO+6PVwdu3VEX57FyMLXORmP85HbbUXQMd
M9acKy789Wnw4rdPajPujrYK3sow2gG4mGBMLnvs0Shh5HO3sW5AV2uXyMwC99rZpEc1+rKxBUyn
OSUhl8dh3jytyhhsKjlryF+Zl1nsk9BRk+Qw6i3Zs6jfBf98Y7uNs6dovCyTaqHC4XNSSDcHO7/l
DS8vYN6xPJfcCE60Sd0ZhGRdmm3TMHqwW91KEzoRBp1nMV8seuuRmaXVa64g+s8iEFv4XRpwAAZW
Qggecjx3FrUy3FsFVQWuITChpU4XyET2qgCQ3FvxqMELojrSVDjxaeT1IcLY5SXC0smsigjqeuGv
l2vljw/DwANGPJ326+CmQZge8HY5fpMZrMlu+72mBx2dB3FWjc2EQXHPd+Hgt19BdoZsQBznGyfZ
Mzkm02RT+1lg13oN8jKsRXo7BBWJYoaXRfV1yWf27lNUUxDPET7f09mwa0Yq5aHhmP7WDUX4DN+h
ujcVyU9+Q6pTDrbadAQcTds0k1YfRGQ38giD/hUbylpnZD5yicdQhLBWpePaXEv45ESNujyVKyvf
z90BnXj+SQHSVK00P3bLJzf9HYwBeUwqmBO0v4mKgfkxXuCt7FNtDwDl/YFxpJbkNyaBi1fpomgl
sQ/L8gYQjYk3C5VeE0xUCyzk+Rf7IDDY8vcJormafhR1jk/ESFUZ1EdnRY9s4NDHRvgvGsweLHbl
9B7wE7dXLnNIlMWH8wrBBitLcyKMWfzumP40UOfId7EMydFYFR3NfAouR+YtnsH0nBnS02AwEO4p
/u6BZp68ziDrjxP+cHMxk07syN/yg0jqvNDrhTPQ7evq48iZozz77W1waexLnP7K4DwTg4EVlR1Y
wF1QRzkwl1xiTyqpgcskFtccGjgifYgaF4kd2+xpR8x7CkQ/Z4UXF7NVmK/8hnKgTmjUYzrZoWsp
yUJqmR9irQaJOz/hjUfiUM8gsqBnyVhMgkPUD9ZNLzFXDWI2Q6Yt0DykTy6umTFyMAT5AvPeVuQi
l+MErwInToZ6c3BQtX1s54OhWAu/jjUjIolCfAS9nuTyYpi6/owY2+wMCfQeQrY5xWRNBxKPToEi
p5Q9EghPw0uWBHYjGmzxB5T24hSy5wc2U+DKWh/96ILaCoBDirHPaRZC5GEz0AqHG+qovsduCOqX
ZNPJbSRO3AsrVq4V19ZSgaegSqHwuxF4qj+SOFeM23jjG0LkLoIzXLOjnG6FRkBE7YtXaO5mNF2q
E8l7ghC25THTp6IUtUuJWlp6j4zl6k97CUl5+Rxqrb6ExtUJxycNljCWsq/PtWrAFMD9CT4icemO
+R4wIOGt3X31rQhLgeBow/amW/RGrqb4N22EWwSPoxuwL+9yC9AiD76+c5EkgRMED5gkrG/w0dOa
YotAqiXaH68TgPQdVINmycLxIAWCqJ1vutcI9MOJ+HA7zu8H1F+/Eo+DK0vnwAXUqagpwKgoOFAQ
UlMY8EHdyCOqXyYCxSbOw0NTgmR5MrzxwJvgc4ATLAUuBykpBBe9t7+UAOdNgfnkmgOOxLLMYuhg
pTz5kQwdqn0heOowaxHtQytAXIJFolaAZCtVpQpcsRDfwXZK1RGtYVc6OZmQ5xcRyGorm3+76ETc
dztOu9Oc63xNS6JN+9ZRzafhh3RUIRJt1zsx7MMsxVfVPOSxluJ6JylvrfMxOLXzzkknQGfVRno1
FtqXr81TgoyUK7bY/F0N7OmzvAKmh9bmdFJfnPJqm5HiMhfcdN8Tvj1axPTgUvppXGFGcoadg+GP
zlIWWsXjhwzBHTge7R/kPaVP7Zzyl+KXy8zrq0b9m0LEOujlvCdnFHF9LCUblEQBlzxDjK9BYKLf
ypeo7hqcos2oPxQx29gcGrJ2gvyJ5GmJIo6dx0xmMhhxGZW0vAfU6VXtTbvER9YfPShmKDIDKnet
1SJl1jN1qGrsmcJ0RNIrAquxKRLg9KqNAsEVcayPRuvDsfiBkQu6OgDx8st7V993FpcyusA6xslK
YwpM72PFn8IlsoC1PZsF/jz/GFq+iKiHD/wEK/xzEMocYmw+VoIDf9v1wdbex3bye4MTQB9l3AqK
2wLGBvk6HrVwo63yjB1xG1OkVaNXY0XW1s1W/mrl94ZSM1dVw+HtNeO4RtwTNVve0GZ1GnmzZxzT
Mhk+OIFXGVNZDcVEVia8QEFBlrkohMA56u8UHAjnyWsX4qxav09LpAX6q9wQmnUMaVMoYVm9vvBs
xrx63OlS3uMuJ/8RVM9zCbrF/mWld6X8L5unXGkhQmjChVf0xM+Xk6D1bdIgKGEJzkpSbKnc3Fjt
6iVzw9EfaUz0FOOm6y3r1+axnqs/1XsQetj3bWL05+kOB7PZnR+ib6JamLIwHvQPHzzHjktht+tx
3qmhAlsz+g94sIejTpIrpaNaqXWz7iOHJQ37yWlw/QMrHVEslDuq+ygB6MsaGJTGTQZsRJAoyWm/
0XCNXmpROQd/0GJQ7haUtLwGDkZbl7b56OuW8nLBYHDiQ9nCwiyVXGbS8FmCuqE7hx7RIk15QhPo
ks8QfEZ12HGcrTYK5yEvHm8ibZfcPFUUPSGcFxAY7391i6ID3vU8/OqAmz0/Al3MPmHhx45oM93w
5oHNCq6lgOOD0FJAj/MpZIVnuXRFdU4on/fnzO1uB1uledlbvZFardfg6w02temoTlm+SoO0eCBs
nnoUQTJGHCWy/ZQxVdoYZUzt4+3Kj4ZbAkXn0WSj6uhVs8VTfuVMAF1Q71wXbG2nkzRIYB+WQrqv
w0fZjggHoZchbvR3sX0yHj90lAeSiPaFZ4xNmLXCoXqRg7gvGmV1zoEYyBJgwVTpPAi40YFhBcxp
NdiCTajUXLnbBp8Mb7OzHLX/VDrGhwYyQEauSiFkvIA1XLB0XJzxyXt9mkcr1zPlhvVFztDWXMDP
fJs3WxxBIMFXT3nQY+iVTj8M4J3vO379N/AJ9+YgIdSWa7mmpc9qzHhyPser3ZrKLIuy/q23o73U
a0PsQDC/a/bbz3U3x0HSu6uNthXyIuudT+jMbSxAnPjEjUVz2WXZorNfCaypzyFp7liUsKfvkFxl
bKeJJtc1C8w926iFoWOJ6BZWq4fUoaVkTht/bP+D6C3L+W5l5WAW7qRvyYh/YBfOBihCwrunHo5s
vxgsHY2RXyrXL8ShYWGQxHsnSF9z0N8mUCibXHskSKt3g6CxjcHnlg5VxhyohMai9zoW79JwR+XM
SH7tHv29mLFZcfJHXYAm0a75hltTeSLNbgmDqdSWRwgHU5cL1PsuKV++W6ybqaCcwimqRn5dabu4
QvlJxnjq+wp0lsJJiL7LiNbIX1ER8j9MV5cqcL+CUfvIqi0URYcyDGhyBTVdac2TbQ9IBzhAbOFU
r1aHGuoimY1XlCCjfHfKka7Ys/YaEMZvq4NwyJxIVNDFgqpfxHE2yq278mb9I010Dkh5F7+O4NmO
kZ5k+YeQs9Bt1vbNKq07GXpkFXm1UBSbfA3yBpFooDNZuM5y0nDNVJWkh/QZ46zc4Zd5ytd/oFkT
tO9eoWP1CHzeOfdVjXWGp6lWAi1mOeyuTReyv1zfuwUG7sIRUOgSD+kSpJjmRbutSIN2ouHW0qfG
Bvth5JGd1zcW2/2/gwBfVD1I8kFWQpJDOsZ4FMIl4+iig/MWYE2cHDRDCFsRke3ydOrqvmJkNr5A
HpBKnvPfs3nDxpjgZkxDTeitBnVf3ZunoEcb0PoTJyl+BfQLf+6LLudG9FHdlD92q4lq0wSmgi8+
XwNIGz1sFaecIOBKJFHoukrKcrT+V5lty2VoE6tyf1SvrmWMLCwfSNtYHKD2sozWT+fn/mOMiBuL
BI+LQWlt5xMsVffW8WDu6GDjLiz+vI0p2GINHLyCuAvMI0iTY3pHTlR90dsQQSt/fWDRe+kjXNkL
T2nnTyBbIyN7fpf8CoN1lPgEO8365n96Ln/StOODk6z4kv2EhfckHVqpbxonuc6Wm3SZAXxuKQ2Z
z04AR8x5BHAWPVYoPlQMcivKu8griLexL37LDE+kHBkuYR4UD4s2/vA6nCTOPGE5HMirDzZCtG0d
WJf8ZKAf6a0cD5wOc4noj/HPANeOp9jnot3L3xpqINtxUl0Bjfg0/L5eH42QCQgYkkQkWZBYssAw
unxONp8ZnAMQ2eW1yP17IDGOkMDGgjtOiYFqdMYWwuVC0jqpigMsLNLfSMpd71PUVWoMMgZTTPgB
E4+ttlA8QKxSbdTJjpxoCPXHs7lrnoo0GrrvhoVIAVJWvSEuQa6zBiwB0jQZSCu7gYLyk2xgk1rI
lLMQ03XLZWdSctrye6bsxXF1yvzZw3TRWrVhQTqR5x5RRo/72Pdiq24h/ikM/4iIDTw8WozF8J+F
qL8KUtr4qs/KvnjyzgCeEDN8WcUp5qXi7GKuXibMGW97J5QZ70sNtliZ0nJrdE2E4lqAMz1WFTO1
k4jSKTSE06IymSX0P/jlBjl+rktyVktP7xvHAV1BGXTIKFtZNKRy3xZx9ftk6iRGAYLdQ9FQ3/VP
a9ujyfvCaj8zKGR3mXXVm1YKZ19+boDRGtVLVbcsY37kDAl7Ux/FEJBn87XJzgWvz7Jc5aTxxeq3
BZaUflyb3feIKP32cr2xxNHdnTFQc7StGDavUQ6bfZyddOQdyJ5zgULLaDMst8ckgq9SLjWqKvfE
Gzq4Zleur60M2498BiICfQ9G2OIFBkqAUfw6y8q09I7kVe30Ppau2U2FWcRRGa5IlRuzkIsGkX0r
wNgVKzK7HVaLcXGyjV1NYtA986NC48H/ku70apaL2i3Me4Rpkxnt/TKTaqHv5pabZrvmSX6QhtPC
VKQONZEQ957PBlD3gFyt3UJHbNHH5HHTXNhx4SKiRRmJUJl4fQX2/NVDgMuOJ9+V+N0Rez8C659K
ZjGxMfd0ZPb+MxDubxhj2B2wjDE+7JymtJOsH6qpzhvZzPcJseptjZJg1M2Cb83icxLNYwDQ+MVR
OlrzlMiWDaRM4zomo4HXT264HGqh8OEVIwfeWREyTzPZCXZxeS0r1dz0owlRwmKxSB58AzMzpfQ7
3CCexrnG3jvFoE9YqyMMNPHGcxwR8rT+EOoztsjF3OeEkg1WT4yNJU6J1zCaSsfABDtREfe2LKps
uBr+26MTyV9ouhY1wkw6OgiNAcVLV/hc8nC6c1k9VbC5nh4FtRWXXm4ET28y6kYwaWj0c14Wy7mN
3LP9f1Z145CdpHaJWX4CI+xjczZ2Ze+YTC+FGPgIJ3J3m+qzPIXJ/e3X8cRSmGiaTVu5APv5I2kS
Hi4PyOP1DxE7d18EsSOqoIobgLYygLYoF7dqeAuwEOZfzRiYjJxWc+wn66f3397DbhEwZALvF3xq
AWq+n9YY4Htpk88lEsULiNx3sL9nfGlXg6msRoZlJZLrhCQQWEEjesa2H4S5Rf/nuq4mLOzW/DUA
Z8MVhoRDsYXXh2sVwpZcDQcvQ7NGbn5W+NICQYqNfHa4hXrtHQIvuryNvRsMUVfMze286W+A1i3Z
XRSCO69Vme3PQE+rvsXmlFqCAi2lYptZoUGoIh5dutlUXWKGKVF9+v6biLM1W2ojUfbsd7iNjsgE
1nfHolxhgOQ27l5OKUCzh3CDcy/6vLHjNGmm5HRWfBNwnD+DNa6/ZS/Qr1Z82ca+eP4NPgmVk7UB
r0WM+8VTZQvFJ4nRp71rYvBfhhUUrXrL8LvPJm9Y86UMIZP3iXdw8fu2g8z/7y2fP/J4/hurwR5T
WaWrO264yCFsSL5NV9gRzv408SJeHVA9k8vG3lpj9CkSPo+RvyRo9UUqmdxK2/v/MKHCaVl2lUgl
vXLtw9yARDhB1xjb+mDHPiSSY4O8uC6p6z1ABcBEs4EmHgzZk/a6YVNJLzXCY37U2lnK/ufXuJoK
w5I8H682FsrKKal2KzlFwA/y+T1JkDuwl7poZxQpHTdDoDZmr30A6i/hktRNFi8eF6VCR9QrHMKK
6U1UtQ5XDi5r5c5dOQPEq9du1dVC8ls3qjauDhW0TXUJMNl2y5N5LP80Qt/6wU/IiMEQoz1bBoM3
1zvR0/3eRRPqZPLzX6qIRvsMORKRbp+/9g4wrljlpBiRIRF4okXDDJ2MubdeF3gkzkCklHJNSkX8
U99VR5bEh3q+tNM10M83UrsJZTKxmnwszgTHGkpiD30/P6AxmmHkt2c5Ok2P6w/CtYSZ+KYa7yHt
5520h9jUuQjfIIp0Oa2QvzJDG9PKlm/BpsfaXxIXspIl/BwzQWqua0xMdHpH+xCatJM4ecOuK4AS
tkUVod3sNgADyg0j5fPLwNGczpqk7o1VhJpcg6hn5TNjp9TSELICNgyJEE53lFVZO8S4mWrMfkeJ
67GkXoiB/ARspsTb5/Dj3gIV90tiLytjtTvQ2UrB0QK5yFWbZCNx30GakzgPFrz/My88lSVAZG8k
gXXVxfQuTv/0D3csIhvGIxJQSzwXkIqf6CeivarMSzoBph0RN8oyudl0w0o444gfBEZDP/oE7Xsp
MbgnxJ9913VXNVd99rLYF4G0FlVUz1jrQMGaPKPzm1p543RmlINg0MG5jj12DVOZkfxezbX9rRqd
v+uW7pGMp0XZhiqmgpAUdZCqV705DvuTpxDhF8o4Gcj54KLZca2CjHMPbC36pU39dPGDIjP99lhb
PBwxtvruq42lETgTaiaCyvEasXRRXvqfXmAxIxlXx8cQPyrThlsvmbG4um4gKGkuSH/VjAFuXQWq
qNH5yjFtyAAV/GfsZ25L9Yza5in4oDly11K5yP24218DESNImoq1BfxlzZ7H6R3AAnq43w/XikAe
a3hnlfaVIsJeCQx6McH6mnZgk4GK1zQcIJn22iDhGF3yIuZVm4MdO8MBocwhRiBzl1yn50ho+RFY
U91mBKrxSEoW9yw7inBFY9EI8Uokz7446buirhnZPznHmW1jb0Qp7cap909VAYuQr/raCaRd6qMB
W9imEcvUq+PTARJ6GxbJ78FNooAm2AgsA/djmEuPX1GCj/N5YjdJPjZfMuhYtQGdCVgVXb906ZdC
Zpz3TG37k2Orq4WmP1L8cjEiNLJzbNnsGFHQuX87zd+yruoEy2eAcVN4qZF2sKXaoYlMJJ6tUWtS
viW90EAuNCSgl82DrLIFa/8yamIzdLKZ1EQxU1gGcb36+Xn1zXkOwnp0G4zyAcgRJMm8/KCk/ICV
+UjaoChyY51a/OMQCuuYX2novXJ5ES1MW7bSO4WXfjPZFoNhAN7274EorMNTFgGBHY4COgR3YG3H
5qGMkriHF0T2zsb6FUZeUpDRP9d5ZQJX3o89bhdZqBpXlcy6lKE80uCYDGih0AZyEEoBI5x2DtDd
9qSwA+qTzyxwUKekkrE6wLOvJQbt1atlX9JRcI1tVBkA9i7Rs3q7lSM2LhrknhfB1GAy8fO4Z3cb
mHJbCPPm0gMf4tEpY8+rlCjXaDo/rbttr8Kh1Xpv4baeIN/+NId22DDqr0m9GNpP86sMLAkAQIaF
hXFayTSDBofACDswZwm3ERSWzIOXIUoobyJiokw8C4kxRj7Y4eV/+2B6zvgSur2myE/tgqCsVu4v
8l3rlbFE93PLuJ+RKiEoIH01mfSJlZ2kV+FgeGsXZa13EVylyEHZD/PeISSIKOdubEQVA54HGujz
IUiyueoMH/Uq7WH7zS9eC+1c5pIjX2W3i8WxNXzcrjviWM+OA2QYNhQY5iM5VPNgJKj2J7liHGxp
xmuPqQxFIrwaOgP6+4yRQd0oZLR1hC2kpDbG1HWN4rS0wAY9TBfMa5BW/TDLoBrWPZ5svvdl5k68
kcuOV0QBC6/JbHlYYqx7At/C7aLa0zGhbXUesvrQylbF5K18rBEQHQPk0c7UNUxw0NOFyh+zueeK
BDTi/P32Ld3vnxEgG1Payd9bJZnKSbjf7YFuvg1QjN/jXNk1ASZAUR0vlPtNX5Y4Fj5PUzvGShW/
3C5up3IzeJ6BvLZGXY3L8onsw7bCaZ1bmdKSJTBHMZxOV2SX6kh7XuwpdHzV6tcudZDvGuNys8j4
IjMBRVJDBYpAjCNK2SprPWtd2uAkLGIjAej2m9iD5WpGCsY4PtVEndeMCO9HFfxX3rmU3eo1sqHd
NGAqomlisiRwJEaC+kIqzQ4d49zflcJ7J9gpSClsAo58PFU8tswr9/mQycdavqZeFCDQsnpWxJQ8
Wfj1pGBlT623n7j4eMfbjtnTMvt6NEPuavzGkbw3SPeQonHeeHbZeAzY/c9xQ2OrAB5bNTE3q+Ef
2kNaZBBOYQwSYwBq1JbBg4NTuXUj7zm7VbRq8IPWz2xqWeSAJRgbb4VmTrzRZAtFPPzqkWnSMs3w
sUfPanUVu+8xLpDLJhGfyTWl2mdnrNp5/9ta0qAXyeZRBjw4XmocMitmv8wLiYGjFd65EKNqcdXK
LyadibHfxDYKloFMMFuCinr//FQ0+9Ho8fXrXy/75WrqdoCeIAUjlmgReZqi8tW/yU/pGdgoIu2e
2mMg5P1zEmvrD4yB/AvTIPGvCmrAdjtjPeYVBeglq2qadqXG8x5mcQWCAog6In6q1zgFKYvRBJO1
XvBFuEu1uGOuu6xKaq2hzmDiZnkjSuBROKgmH5DiTJS5bQpMOkv4+Qa8QdPjaBw61jihRgq3GNW9
QKO9Z7K+dh5YVoXkPFocOltPhSM38U25HLu4xAupoSilPCP/1hReLPlaOm3TAUaewwBJ6LitlFoj
lPdVZyarf1mUhOT8dQu37s5X7Eu8IjIl92cto5UOR9kfUnuU0QZmoJeWZ52dm6P0goIwz4Y2xCVL
lS33/G4HIww/sc8jb9653PdfGr/BMTpFGuma80pVH0ISbYbgHJKsF7KvbPAhi/+77j8MB3WMZVfP
K5qsHkRxvrAfcMNpeN7vTNj2w8Zt1XXB2c2ubsfEIpozg8SoFKmlzh1cVUEk5ABepDeOWEpW1GGS
8WroRo2kJ924Slji+aIjTGiaotFeAX9wCGxDe9cQeDoe4MzEJSDtGMp+t1C3i+SyIwMk4T/DcOIu
svshUrQoq7EZua1ZaOTclH+OYhLiYS4fzmSQ10a8+iI4+hYgQZKoZflB54o5IpzYly7NstyD5LfB
c9lQVuW/XlqZsjgrew1ETr81lMNJ9A+K+1aFWaIsYEqnmFEQqDYR0sLRkJ/XcIzk24cuUSb7/9pW
pdyDVjsY7Uo5tSf+0PQvwN2pVugTRnwZec0W4uyiWAktB3Pbc8bHjkUSz7CQtIFHLFIkCNt8AMbw
lp+aQlUeBV+g+tI56oKrt3kCC+krQpWNgmk6iYTkAWNFZ8shWpW+qKWOCbXCDwuPincZ54ESj8m5
+xGjgLo+a0CcAnTdfMEYLjWrHX04C8peDj4UZZf6WqBu+NAgGz6NdLry1Xhv1FGOEVxT3qIaQGHP
F+bn1POWF7Jk+FpKTzCTONOBvWrCOEhxufQia8d5NDutnYeS8sss3SUZjyE8x1DMy/lxa98MnPve
Z0h4sX2qUqYXCrv252PJePcq6BX4kN/dHy0yER3xc8isL2Yuu29fa8nz4O8S4GFp8xKOHw9HK35T
Tpp8KLFWYLma47AmqDIv7tcAADPFsAC4uszRoVjp3FwGvx+lWIRn6lz0XEWBdntBKWzGUl9BApHN
7gbHwKsyhNHTQ4MrcS+RRgkcGpcFUSqItvcL/yvVdUxY5PR6IZdwBT49b26nnq+WmJ2W+EaO0bPC
x14kQC8i92FG5vkq4ecloAmTsi/umRDfD8JfGOO4yxlynRkSIC6ptsqiv/dUe3kAX/hwu6xVre9c
YouIRM+NjIOvXbAIRAlHJNoW3nPZe5UUSAWoUjRx3fnUfgCL4lkprG1mTgiBZEWtp6Dr4bqxbr9Q
GiMzByZ+7ubirj3mKZEVRbV4UHbJKqSG4Z7o9oGclDgIW8h+AI7F9opZyp3XAXVJj1nH0qqdGbVw
ZWSJWal68ox4btU2ll5nhfsqlL2jbN7tQ8KffszhIwmhLPJDrKdpV+dvXvqxoSZaIzEcwBA0rk1m
cN38DUN6yA9BebTj4caB028CHg30K3ghbI6xHJcRDthFD3xtw0Jt2EUJqrjYy5DBZ4Jh5rOTTXn4
bKajr5ahtmE8AWXy3/vjGlIxXpE+2AN/4B+ZGIuYIE/0syy2yaTLczCM0BxyfkJ4WUGPjPTX5xDy
nYC1/WghFdF+bPjn0aslv5TNr0cK+C3ridTAL0zRRQBzzznEgwTEhbdBAs4atnC+NpRxdZbLI3Be
Gx8p2zsRjFjtvZlzp8+Jvk72OURxEciDifbzJvhVyWKxolsBob2FgSQb64nWomUrSZC1yNzSvda8
0S1hoJyIzyU+0DdKr0aKewtAM/kOqgy4cP7CvT5ZvuGEmncCOOkWCTSm1Amfr7UgsCf7SV07r3rc
uXpyQpInZywRp1XvVcxEPGVlDJi5dFiStfqPWp5L5eFfzfpGrqeWPGWMKpCK44LCkeHEZnCGJUwC
7si5HTDhvN73DtEQLwvWQrzIMaow7jqrWEG9xbuRrhBJilz3qDGqSp87+U0sZwy0bsb82tmjY11y
VwKjTwLfVI5R/CKJj5IBYkiTC9M+eDt9eVK/WgTOlJnDdSXmCwW3QnQqyTvX/df3bUKeaMrfcq1e
J0URYhRSUcKFNIggsGMeEoxDatgLukcgsf2Xn1JehrpP9Aj9y3us40cNsBuQGW3+RK+63uxcch9I
aElXv/TsmR0mp/HP0fpRSPNmxp3HVAxsbdvLMxOnuXQYDF9oD645De3sswUa1g8QReXt/9ziOZ7R
WRkD4vihttospdojTGm8tHGR/OGQ4gmpbK7E+azBSPTNYr8ZnBy04P3rJtHbhB+GEz2o4Rs9JWZB
uvJYs+4dcNVU4khBWmvEQLSLECxWF123ps7necVwycKApjNPzn1PLiwI1cqSwsUx4CQuT/2nXNfi
HC4RzFXm39F3GiT5afLC3MFBPXRKd16mClbkRAG2MiiHqnwk6p3yXmn43dzhw01OHF3/eo+aYhQr
4/UnmfAMeA2hnBv+QKk9POrpmuzRIcvcxcX77FDSHfonu3FGP9lE6eJDWcbLgKYdVux3hl3izyAG
zT9JmYdn6ApimyUKKBM649rlQ3Jaf9f/mgSPf/NMUq8wWenVAJagoCkMzMFGtV05LKsqDlEKw3Xc
5MR1SE2+TDBvzSS5ovqan6KNxDf+8ZNFSABRm6n6t3UWGxVF61EEp5w97xb0QDqXR6TKeJ2pRQTC
Sr4FfGfBHcHPSd66Wwjy+QBl7cSgjvsqJKQcQAIgoFt1EAYsxrSqj1AkXM3u0JrqQI0nhhMiMFDy
PH6glUcgUeuhlJgtdfQoYxq+i7ywCFw4H1/Vmz0zV4KMYYNmWMSZO8YFoIw0Q6lnFlA4nFH0yy1h
T4KSMxnYOdsQkOhCVdUoPEIxHIrdBtjhLgx9KNhHpevRIRs6PQ4MJDlC+/NUdYRRy9Le2v8dadl7
UW+vxSeq1i3AfPTbXRHIwV4vYhNAxno93BWmJDjcZZoL8hSPRH7GmoE6o2AgcWg69W2sNt0lRDcn
OUCoR3AIvk0avTDlnOyadWZ/21ma9N0PsHxrCexUASfR1NcKuUxnXOb1axBex4AlQDPcCg35Egqf
ZyqV7CzUmkwzFLiaTxyIpzDiJQcV4a0Bqxno57Kt/s5thn1J9/JPb/J5X5igQc5W2AxeJufLP2se
1yqGlzROMDVhsc+zYpKx/66cC6FLsv5J5IKzA6/V7ZTuefSZjai3+KNOPV+jwJp1r8wyadyiFfhZ
7GCRVlTC4jYsiqbqGhYDloK5dC/DuBmDMgjy7E+gBYlbj9WOwdZHnuvwVPZ/UJ7HGgv+uoaVJTn8
BidfWxOrVspLbfbJaNLwsUBgp5I/Rb/1wSFRIp/YpLdQfG+C2i1ca8VBWRFK/+vVvBHnfFMaX8Qf
vsRCaxIQa3Ws50sUT6uMjgfxdV3LPn8jezgwBGdKdMxBSLK4GPJORT1ukQUuqUVJgDyOLnM+DRbD
DDj4SmITX1WkWDtTlrl45AXAS+Y6Faj5TDZAoxEX/JyMHCmZ5CCVgRLRK5CArvql3UKg7Xjk757a
EXvgV9VejrVKTJVAine9QKUJkAcuK4z017RNwTGJj5aswc8aDDTiGB9FZp1buRBr3CKeMspRNbrC
oWNUnVMHg5CYszOvjxXQ1j8lLx2FhYVpZmaL195N+EndsUR2PCgUAUnaDezPcG7k08uL2h6V0vcm
1yJxSI99iIpbDfIzDj25xVTY/dOeTj3a4ad5UsC/fhkoiUmMjc717rgc2PRnbIjwAOLmECgp92pd
AZ4Xh9NuHfJkM2SXHkFZ2Yzw71zAm3cCTjvC5NHeuSxrkvgmen7ebb5JjDGUkUye2xf29nj9sBRl
QLEX5fMW54bEAdfRFp5ivvT6hr1PcCRhiu9rikJD9kqqOGldNlKX+WXLccvWdoV4VSSkJ0M8jwX4
ruspBNikJL/GNSYdfQp4YcFoUfJxjmME8h7Fkl0H6e1nWcbO+eIt9yANNnRUmo9k52FVZBGs1rgc
/zOFR9lwKUCz2WPmAnIDjlp9w40YK43TXzaKMo3AEcvw9x0w6tbukfBWLLysmT0RBy8d+EbeV5Fb
2oIzx5/EkpbGzjpZunQjFWqUuoAXTwtyFSZJIZ/OCTCmbY+iEWI/HFdoNyG6zXRRSs0q3GEVD6Un
uSkwRCABv5UfhkFVwBF1sbkueOZMxqwVEGMNr6EFvMsx5RSXwbLasqyOpde/mCz3oEQRJFQvdVIY
w63RVQm/qCo6+i+XU+ufiH2ivTcfQ1AJj7bAhoHa6PQ9i6ViQJOxqL4RAm9I/zkQhWpfvyO7JzJe
8UUeNS8/AogvEkf0vDZ0GQAJahgLV9B/pq7ZLD1Ws5DLN6Herzs3TReYMyu6n3EctRmrh0GtT1Qg
xVO87PuFjDY27l4CaATYfFSznPt4bBsATEB44AlFd2MjMXL2SHpLKaVi2knMtzqmCo5UGcwlxCPd
COOWz8azArvuRJdg7Em9FO2T6r2C35gThTJeoitA7kPjADhZbSglFd73eEE/1y6vrrYL7iyyzdxU
wl3Hf7I5CXcv9mpaGE8mVQe6xesROKvU0uQps41WPQxxidJl/Vw33iSV2DYhwFDpA/fqt0NsIytT
UNOPEWH+XIywyofFf3WWc/Dwzhkhie/49CLJ9Zm/Ie7o4UVpXHYNNrKMaA06axtoVAnAD+jHwknd
vBSzR+RcPZXV6b9sxeAJ9aKB2BzsikEbn8H3IKhdRUKzBzhLGL7H4nlIbWKTR4jQE309lXZZSAF+
YZYyxGwjNnAvVGL6tGT9ltQhZMdXfjCrJfAiey8TCdAPL52kbL0L6GIah6ONjL/dFf3HdEHzSQee
eL4kdbBx6uLZ+bJcBxJ5gCxZ48ANLOhDCaq0oMNO3OLNZopKbJEmqGw13DxcDJlN4XuiTAGF6CGK
aOUz8DJmpZ1eykJvIqt8+td+NMfOZhx8wbuL0e4Re4fDmxzir6m0vzO+f0bUpnuIi+owr+DREBBo
n+obbM9PcOXKkTIZ20IrFtvruZBA8pPHRhsBA6RQv68plVEhmcTyXrZ9uzbY8+kbWnizai23qrJ5
Fli9Efddw53OAH9bpd+Fb93o63kHQg6qklCVIJt34y4TEY4EhvK9xXky7ZuZOnWaCCUWnVyEP0Pc
DiysbCzahN5tn1P81I6CMLmMwW6mR5FP2y5cVP0H41TTXlia+ZSOIoOKxI6XkXuZtWkOTWc7ZBCr
JGyiMJx4AY0+2bGXBmcGHKrVCoTbDYukiqPb94Po2WrI0I4AAcQjkXjcKZwQW9Q0ABSFT7p9jMsH
FnK4MsJurYfl6n6JYvwiQ6C5d2qUpk042dJ1sNL2cW5t9UY0sKxqlBMtNkmSml2/v2a8hmSLZUCk
vFLphi0YEbMpWeF4kZD23bjqncDK6U6we4n6yecgv1r5yy2tsX+pElqJK7LJzO64Y6GrTkiQQHnq
kob1PLlEe6bK2iO0Z4mKXoFoNymc2ackVA/YaxEAugXo7m71rwEETJR6QJbMBv9hrxbX92LwFfxq
6v7tweIM1/8pISBok0jYCuX1keqA9cetBseHqEKgSjg9sT0nJYV6qGfHgICowIyGpYwCM78dBO87
7Ow7GOAVSEdtPAVAyoocBaO46KKqTQvoMKUUOncooLcKZpUyE9JmDp/o9vZFTjWbVOROGnHBuFPM
9TfI5RJj/EHhs8ITQGqZYqqwlK/obzwLtdmuuxDNjV5hWbSNCNo4Nv7oZjEVhTe++EIJ5xOEx70u
7ZMMlQDzZpU2iCx8kep6QU8qVxKo6MQkRY74Bm/HKLfSCK2ddXUc068sZ/V4PksCAKySpcvvmtSS
baS9wBYF+SvVvSggR+9SB5gQfW9nigffv3jKmct95NVMnQKuS+xuSY/wxYL3QPAYvfu1E4PbyxnK
1KHc+C+AN8Z6wkZYjnuGygj3FrKyX0dqPBCfmJhKLq2iWFrYzNl50rXpVBNF1n5tsz9ABX+vCK5t
1Tq8T+RNwW5sP2HGTnhoieOpujXR877xVLARxqsPNdjtqbJREfBY3U6OP+5vVgdAWjFYQJJl5wT7
bAMddMCGVX+d9wNI9U8Xw5x9nKKI6tPtXhwl/j9aPtsBFRL57luWiwXHD/f9Nl5K6osL6o5RIurG
xmlydseFmR8rVrgs4Gu4cA5f+tHAoAyEMcDzlAV9BrjTGhFuhl2zInSwU4Co/xphOqvJ2i2s7W39
vSy0nt+hueNc7yIeHJwi55rWWNXrU6nwT36GLFD00pyrEU9Ex90cTUMtjS77vdHtfRft+z/XvnXY
VxCOgoa+EsACRj80hw5JyvW+fp+ri7MpEMT0dfUrE6k0v9Ki8OyH9NYbgmuSm82l+Y1NJ5tyJYOH
fi3EKhIRyOAL3vaHdh8Ogn2DG+lFbHBsXuO1dkilBvdjSuUo1hp6ill/hc/JBRcEWGSDll0V/oLm
w4g1n+qYQWVG/f3l7sALiE9e8gb2SyHwWTceQMXtHc6yjz4azkipwcDiMl8DhqMOBjsI6PnCTrFP
baw28o3vE/zuVtET/FETQcc4uZvo6TZcT7zktJrTZXBnos4JfuILdluNTY72M2nPJ9DwhXai4o7E
tF6f6nb+0VLZMP0NkJcXMppEFafno+2GeHDZe3F2UIq0x8vUIEWB1qgDd+EPH+ZfUB1JFop/Te3i
BcZVcbPBiAzX3BGzRY3YLaxOPlFVLI88D+RhNU4Wv1AWQvggghuJ8SyXxOG9jOJzk3dFwKEaBIhD
HsZ+DklJRrGub6OoFNVKaZKDpDqMINz/Ykf1fgTavzn6Q6geDL07Ga2/CAJR5ljCsFBU6Sje7uan
vqWD0j06/bb50ERrtWFdSp9XbGeCwP77VYu82G+o1NUC1OFevlieQkyfdgE6Jbg+iUJvzktQjlS5
0Li/rbEZEBctv8aRp8iv0qGqeqyE8Af+IcnVvn+cxrcTzzeW3NzvtFuhF5dGSuHLGqh9N0SIb6ZW
2gKYjIhumgCNaNZR4IuBDCdmKzJFcB4NQYH076TthWY8zNYRWVSxITiovRj4zVxYQqBcJy9XcA5T
KbWebmMp8xDAtupje3xFxGTqkoRicHX/XNeujUe9yuxBBZWjZwqKUGyvAqUmQAVYoElfWpd2AoHo
qIxCfVhUXlqBPpuTM2t5MSt8WXk44aKSEk37H8lq+MiritWqYDk5kHDuOSOpnfZFpGyBfO0FFHUG
naLi9ZW0709wTRtHV/akBTmBe/THxghxIqn3E32F8pVULZZkX0GMHyHRyQTZBePaQ0rUjEL+F3Hl
P1X5FEiIINQSKZ/NPmJx3RJKU14RavnROBnCn7ZkUAC7dL+iwSqCzUCAMjHutVTsm9gNP/wXk9SC
Kh4wgsTsWd8e6AG8hhN/uW6FeAtGCEJnP3fgzAtFEwO3qW6rNAfLPNjcIR0mZz4gw0hFi46oZzNv
YrZ/Xb7qhEEUKHAKZ/2jRd07TI2yiRUn4BsHnVpc1XrCNb8yfmcchAI6LilW4PkyclpgBtEyCnW1
DRSwqCTafCsBE7tea/iPsxJUxCs4vpvaBBwSvWCKi3WgOCom9ULT4+18Hnf51JQg6apX/v2FwdlY
uIwzzSYq+KXKgmHU6e56qMjXM1NDkipx+egnm3O2MMvqmMkQDv/PZfaseztsIVoFHRfIyp6TNJ2f
7yLGIbdcl7/VauTM1jWbCgrD/Q2UaBZBS+FqlkfwaDgSF8xFhTIJnP8EwRQeTFPLfnZdGWYrUE2M
59bz0KhGByIxJOE+uYjNSSB3TBq2sWaOpukpwJjeLTfayG0LDtbCcFbrQYNNaheCMydbeTkn10EV
ky25G/S+bQSot2NbBro5awf8s/JqLY1jYnrAwF+DBhTwk7RXVDeA6SzxrM8POfAmPgQ0f1kGJyGZ
GyHjw90iO8HW6Sc45aZliqRx4YSmeAEQ+nChK+zfqVoYPeWp+imECRmoeYdrIBHVegzLz3+z2wBD
2S5Huox68xXm6VAMoRuAF2fLW6CI39PpLTkVpgK298mFkeehUf8geLPmfCrgEe6heotTnKu/cZrM
d1cMGVgUQWGYaR4wIvfE7wYOmIty7gkxdqgwYX7MJ2Ec6OpPblenP1VJPHs2O0In2kUEVddgOKiJ
1ZAeNtMtGgf+D+scQkuI1dc/Yz9PWHLs+wc/aQ1ZbTL+XMLfT0PRIQ0Nrs2Lf2lCfrrnZIaafLvQ
GHRurM/WMsQtkCG2QqVHSUz3CDEX2XvUL3gl+7vssnpqzPf/DmxbNW+ffMg0yzXhcuI+77ZsS2or
uME/6u8ZrLrtaN+DwkkziH9g4s7pSE3DVnyEuN2m1HtDQfK9O2NJWWCATrmTasDZr0dl1/tEI5fZ
qjcmbI5Ah+PQB2EhQJaD9oMQpJrkgsskOgAKUuG4P9tiHfPGu9fYcpgFaJnlvq1CX/l/DjeVpiBu
dcPpPK461T/lbsjAXPZqlIbGy7lIWNu/4+bjIy8nWz3nK+ChYFDuNLhkiV/92Z/Hj53V02ozxkkr
s1WK6RHruztXcwSqKmrFELxpHx62ouZA3ro6DVRT1Z94R4+/CrLD9qDVczhdF8xvs5aPCNeZuBhm
DgHSun6ERGkfr1CGMjq8QuoMAfHr7MEN8+RgUT3mCsQBC44z1HHsQeKwYpdEhIIq+cOCjuIBbPMi
qN4ZUSr1OYwqWt5XIIxTJag5GxMpWWrOUmey6ZNh0DJAes0Rufx9sDf0ggm/zLhKvlehAdN+Wjmh
uJb0FQUapbzsrYqxOBTyOBitSE4YxGnyfT0EFuxUqWn1vStZLK2Nn6P3cdi6vfgKZGhwbnWwcSyG
zxaVmUnTt8pc3k1ocHuSmCLPD1QXvfX34VRLHI9p2lWapJb+FHm7Fwig+aCwRHiAYcHFWgIWAksJ
TgBthWa1qBGLifCk6O4mplJhzo+rOJZA9O/2Zn0s4fQKKu71BcVe8fyeIsFtIOOBeKrdQ702g3Im
i4oaNZXeem8NL7fqYMUD7VwtR7qCgmgBsPeAzg99xE9tAScrd1uNhJh61zLC/FFyQ6jwrq2pnVRi
H3Y0sLlsA0K4x8p7AYDGOuurSl5mzBuarvnuUpGH5nI/q/W6LkVk4fD0p/Q9dCCJMk916fgugrhV
tGYE6OkSk8rYzDX5+Cc1p8l+YfETaw10tQ3t9Tb4TGwsenxQ1/SMDfGuPT4T3nsYWq2TRUE4bzKX
OTfJUamGoLB5AOeNDFYbQoDTCAx5QH47v19r5R+jTCiFCO0Yzo8PfvB5sPtbwtIXBYfA/a1WB7SB
t1YKdS1zgctva1uHdFoWbQ9uGUoL5b0tJU74zysV5MDSblRfK8GiTt9w+Grvjt4Q6ORXuz34nGSw
q9/znKeu4MuZIXa8U09BHK9v6cZIEQE1N5dxVrNp71TidKnOCpQUxa5zANtuieXzgB53opBZxxEO
9roD6Yq3f8rZy4K6aUSygAHDRIbTLGikcpw0m+q6AL9cxYVH6vnKFTOvgU4uGWdIMU9o+0uA3zgo
D5rBv7zNoZ6XA/Do8b7BEHHF/tCJm0dd3Tu1FYiaFK7K+0WiKZbFwB2TipW0o9iucf68tI4sinM+
f2Guhrl3SgS+vVWQiXqXRWi45yKez4HvDw8vBqhM1TVGl5U6Cqz76Rbrn2Q6B7Y3pwFWYgVvVorS
FKA4h8thk6sSK/cH5B89W0PpSG1bbeLZEf+gW6NNV+tTHJNvXlao4gEhBetdEsAL/IZgsdvPfq40
QnghYa5xtprXKrtuwgwB6fPm1deBISYdaWEeli0ED+OFTke8vYaIa9QSdK3yoPUKLUAq6j8792rr
429PKvwhhJiomaj+MLmwNWDEq58hxLY6wDJjXNypyJwjscopplwrBXJuV7BA6XM50U529MqRludR
wEjm4C6AQ+4MgNGUsm+dYobzGYglZgWJVspokFO/DT00MBly2eSvqCVvhMwcrMNQZQEC4z1uwmGJ
fUREwkk+F0ziihmfoY27REsXLFEQIysXq8JHzDgiizJTN2OQeELcBqjV4xKJES+FqHTFnngdt0KU
nixLD76EfDAb66dSRLnT47N3nCRxjIhng3tjd9iw59uY4IGreFj/NSevJiXLBvzT+t807tyE9igM
Zyfn5IT44CXc4/eTYi0pHjEWKW+oTdQs/lg2V9pH/koRbewSNYslMus6vTLXQ9wrLPoiN4x8u5go
r4RIwRuvxImviiwfu5E5n1Nx+uTlAKYTWk01A7QlXttCS6ujvfd47Ld62zUmJbUDnVt9ZX6ABUbC
FP9tdbBWNcRl4eKW7B5xCHO9/M3LzAo2gPJOnS3Ruq6zx81fkH/0QOYP/4RPRGe8YGrH07a1cn7q
9qGNHVvDlRU+JThl+at8/ocXYMxdT8C7MeVG/75HG8xyfFmcA0X6jk8CnoSlgcXYLCgrVcWLIA4G
rikRQa4u87TUmnLhHxP6ogMUpc+q7C0blMHx/6bajFpk2vCSupUQDU9hX9qkvBy/63R2phywfU+5
p3gKGMhD0pWX846ss6sKS+0tsrNB1zT/HxSOHXGu3LvO5Qy8CWuT2U6DlIoBkfdWDICMBk2ppbVT
2no/WvAlOqRisiyUdjI9LnHhnxlMYccUj9WgRWtZVi/BsBNsV+Mbkk48IkQ+K09JICN5NxYka8P+
w3Y/1z85N+Q9FWEIzyrvGbdwmeUAZX1BHypamT0RA63ODEkosTVXlK+S7E2JF+30K4gn1q6d4NNl
WcCe3ZsK+hkntmEalWm8b2wK1upBG2tnKX9wNKa+/eX7rlDWcH+gtC9K4L22lh3wcYC8T/EuqJ7B
9l3ZJrKhLT3YJCoXaOcCNWklRQ7b1qH6f0WcetCDzZvE8eyMkEiqOy/zIb+F5HjmnSW+2nsRdCsP
xmV35ixX+LZ2mSlxH1rknA7EGynDYUICvwh1fhC3fP+HEj62DPdCTc+i0s+iCXKlymYTRXmnl9Nb
uS3gDu8YN4/eKb1o8nUUyQ6PIymV4gynVgN7CrNFHyPxhTdWETynTD2EOu6vEmlg1ghsskffhpMf
ghpFUXJRb7wW3ILzVqo/A+vhzwzpD3M3hlUzrbqrVxaPxOqfdzKwZNGaXEScj+dN67rk1H4BIrZe
WDRZKZazGk7QglGV4TYIX1At/nxf1JurBcUKkRziMwrgKx6lLmlIca8jH7IM6UWmd2MXWBEaRyVP
i89exPca9pF+VkHn/LdNQ2BOz25IRa2ygLKroAGny+I+tjwFMdDfbtGYiGrGB/5gTm4/xgvXbXRR
BoOfezAwUIn/X5BB5uPRoBxCL1OX5lxpnSJx3wUDQYLz7U4Ooo52ytjIRu94LEtO5ZFZ5shHPQ/v
J9Hw97U1eFIjFLYV8TBWi4pNaJB6mdj6QBIb9sqZCOrkzIHs2l80alG6RxPSU+ApgCnVP3hPJi8o
/lCgtUFbPluISg8o/4TK+rdu+KHtBZn0/5DqehcWsMPwXO+DVAWppKABawMvMJ+kjMME1nVVTmXH
pFvkogjxtppwRRbo+rMq+kzwewxIRPOyQDJ8z9M37AeHSGQn+iUWB80100qj1KD0oW9pw81vCkFf
2w0eJfbMAk4ipucoybuDo82spscOowbpV6+Iq+AjXvNqUNy8QQz+xjDmDdIWb7c1gpiZRF4W0FT+
lUbxwYDZ/uAkfjZ6NrxQQZ0HW/04vWe1fFDE7mR/4xDXilv1/f40LH9Q2Ju8OwBXdcTWsea1blaR
zs94ngJ9q87wKipvSeunlK0dwcu7BOXXGZnNefZGLN0DuWnin2LtYxiR6gQmcYbwH6BdZaxooYGc
Z1B5Bbm7t7b3MlRdptMYO13qT63YZwOvDrVBDBZcsymo+3Gd8JzAycIbA2y7ETK0tQHRjAJUEidN
5yFWeIKnlC2GXzBUwArOQlA5dwNpHXzAlcVJvtuSBc3EQA9D7GlLtVl9S1cXFosmd89ivKRnNYeC
brMGov5svKVQJVRjFXHWgTbxs/BQNN4wurJp2FB7snqdbWZe2FN94/glP07slfFjSEAxCqufVmKn
b3P8GY2CAAqsFJF3ZNNKZa/HysXYqeewlzNnXJYUGs7iR1vACWukf9RkwK1yBGQVgIiuAhks5bao
MrYO5bGDv6z4w1Rftw732H2pROSvFQDphNHfR8abLOvn8d/S4eWmgVqxBak6UMvG7JVvb/FpYQqT
pjv7FKvmrkTtGK/Z4kpaCw+qUpXV+xbjv1VizD3u3fiyOmrtJE1R0dEwtjKW3yH9X1najbiVOjkv
d2i+sRNgBHzReHH6HTMeB6oFkYVqLShgnTT75XnlhlHjzM8VPlctObDpYVPCejWDVXWRiHu/JDaw
0/GEmcpCiRpQxEUc1+B300zDdf8P72vctEZk4sXYYlrOSd3bAL07H//uXxI1pxsT0sQkZUlZ89Kn
qAxxOpBbiknfCgvTGC8dnaqxqdKi1hH/h8+jG4+ATMRwSvhAIuO7lax8NSjccLdha3q/8sEDK1oj
L1KpljiGdHCAQCUjDHsD/mge/naA7Td1aplFT/BMhMwozBQbme/xTVA45HcTTOMajNKxlCgamwAn
2yGm8WQ3HhYKbehcD/B92hCbxL0pJJZd2dHk1EkflzlxhACJYnts0c2P0A3eP8kmLQdV0BFPkNTf
KIQ21Dmfcfz+hrEEPD8eN2+vNR6Rv7gIN2pBjawhOZcIoUPThkgaNbYZvzM0mFKX7gn081v2CVmp
OHcG8eDMl8kvOAGQo49LxlenL1INzktsSCd9jAv/AF+ZNCBNRia7eKJMuO8pnTcthfWTTMwT4WHI
/O0LRepib8UOW71xKutXgdAodsoUI/y8qTZEZcIxL2kyZ7oCvCHjOzBXbylPxZ8PqJ8pOFBL9CgV
rZNOdGBdO2UzuLBIz/6dy4BbtzYRX1feE1vICdKog7v5Z8PrgsVQRHkzVU0fstcSKPPUJf3Ioszq
0zGDq9SnABM1McLAswD+WF+tTvA5yEXKyzdlxZToXRgfP9kandXNgeV7N4QzA38vfKasjvDONxcZ
uRCPocX7eyqW0bt0oOGQcfPyYtyStHX13ThO+ovjaSi31tdXwF0TYp2D1jru8/5DZFJT2PAQAU37
ZtTrki7H/WHWKE1xg9L0+8wrGFWItSLzaS4Nj3F+dyPL5Pm/DBiJMdRZh61OXlfXVeubIsXRDRHn
7VHYQs6h1gyJhUc8yi6/vXTEXU1vbYFybcDLCMW0IS1w7hEAiYX8EkibHcEGGdp58YnGeHc+pacB
BN6Ni9dRzGEe7N4AqjzNhFO+aG5V4fd4rSsn/wXgoMDdSL27V0Y2opWtsYq7SU70G59MOVC8Tb7/
6PB2cWYtIHhS5Qo6xYIuftb36xTdfd3KjAIIczTNuoiAAFjLo8I09ioNUk7foJc/vYORdqiQtyhd
8DqG5iw53ZD9UCtJbXkAsaLryJATMOT//f4o5QLNSbIZvF7B6eaW9u1qozsKhM70mvPBPTMG5F+Q
LIYYg9RDmuu46xF5okDEwpgsIA30JOfYyNOy7tKwhdgzXPuqQpH4hPT5TAv+xQOTWNKQyVEyoU0b
zE21R7YWNqT1dNSygBIf3LpUI08JpcM/HSU0yTdkEW/RFGMbdjK7xxXVEvfivkbZUpbyBfVGQ0/4
qtP+8OhP0qIbI1tk/wrUp0zWhzzUyT8FiIuv1Lactz39hpvsJL2DBEPI8c+ONGOZ9z1gmeEXE9xU
REMZINkt75xiE/3np2tLDaGS/YmgBAYbMk7LsUI1cL084IXYYDiA8yTjNpPHXO3ChHaI11GQ9RDk
BtmrpDtD4gm/TUKtBCZ6v+oZov/hFMGXxp4rbqqAA9AvTmQBLBqo2pCRoW8Cs0sLWzLMWPkWoxFM
aQ/IO201FXaEK44asVludKOCscFlGAm6HnPtazS3ZswRnpECkxojgwuEkbUixmhEVV9m9GV6uOQq
U1YyPd76GSUYekEa+Ukgi27JiO1faV/ydxat4SFVALsp4z6L8bLydzx7KWv+6epCNjUDfnwAjsnY
nAPQJHWmcEJPtx6xedZ2xZld/lPsVKcJTc3rk1pjYJTjOyvRrQyQQky4NmJAm3TJ3HMrwweaZLXt
aasUYmIliDk4wYuuZcr+cKrBqYUkod9ypFALucdaYle131G8BoJ4/FOr6O/AOrkqAp90IfRthcyI
/R065IhnpCH7cO+0e31ue21NtaKR6dilAZUMMhuCTLw/CiSwl2j969g6IzQQW1Xy1d2NuI7ddqRG
ZJ0mrNjlRGd96W6q1t5jaYWItCN3WQaGHc+5KDLpRgJ82PMgkBhVl4gfFiGaW5PrIeoKXeKRTzSk
IRFhA9C9bQoUELOrPK4659+Vz8ONlyUPUt7tDULjHYAwQqlh/wNOoln+3AeenmkkksJ3cjFmYMVk
AiOxwYMovgvurvp+L6obaYjpB2vvwpMjxalFVynt7jqtsejV/skiQwDL5l95VglymYn8FVGigeoT
nLpvy0sdvUJIRzGmzcNmezw2yAUrE5ELyFwGTC8/+Vk0ymevqqnri/nxrkw1uljG5trY4cmDjlcR
PeDaJa7F+u1UBFTnzVBTeK5LswpsbyGhqhWUcI65bi2geVkj5QxOcyOo3jgStp2Y5nIhO/P62lrb
0V4mlSnBAdKuvStGOMDf3Mpmaly94DcyYC6NynLnUlsBwbhMQasUvUNIi4fjvnHdnZIJdVfPIN3x
D5mp3g3FrrnzuC0VBSsKebpmc6LK0fhowtgTXfVmG+I2Zedg8qxZPiXQ0WnrStvhzby1E+8ouMfx
lRJBM8nlQDKxCu1yQwFv7lqrz8xr5U2f5pRJ3esfnsS0OJs7FDYq6p36lCxOmJPpTrEKgPeklDVE
CsUnxbP0rrUISbF0qd3MZGowJOYUpr/g/2X47tnfvUDDk7Slg1fAcd1W+fvarEH34ikiUom6SkpJ
PDl1VlFAdQWAdqKMWgqIGwiM5wAg8twHfgx7PzdSzBUri8F2zkm7yiywfwG/Et3rrEAe+kiIhpjH
VoXEsoez4pR1U2Smqj+xWpe6vOnVpuFVPKNWTpA5HIzqdpULxm3ERQK+KM4Y6IeqJA9BENJrEgIx
lenkVpD/OWYanseT6LVmNnWp13bKEczXTwsYdIq0jC20s0Qllif/F+bqmrxcNOlsDhwspdnPhVjI
WY6qdaRzW1Wf10zJWQM4IKj1Pz7D2nZ8MJMbvwIlU+b5XW63mwB20X9R4HXy8ITJZaUtKw00JWf6
ZuajgSvE7hT08sPzcS3fbMNBZrxSiBSzR+FxRjgklyVlyScU5vCFVUB5TS3Vs/s6D6RfqxPDBblJ
jBvnQGiJRTbMXJkTy4oNKhvoREV5gRZexBS1beVu9XPT//qYeprhAF3LxE2VBcAE2TBXz4EhM1pV
4iNTpjpmbFb+TaZIgFlzZ69vKdSbGBgvzSlwvTeYFWphJ0yy2bNAvO2Ln7288hDxpI0U85INd3tJ
u3Kj+l3R+cQ+mm/ph7zUrvXTJPy5mLYFGl1RZzjZKU6sveGzLP9JDNOoReL9BZVO9A2GZo4oyRI+
hQI5E9Kt7WXbQKVwYtMuVKqIOskbvqOm5UhYrNZZmAcs5jaJ/mL+Pelx7sRubcHOsl7KI3BcCDOb
k+pg5ltzSWFBn5hts5TjzaYAFg+f7ynziDrQ7o8o/ScRqxXUHkqOMM8i0wRmSxzlFO0BLhU7/3gW
OjFmkKkBJa5SopCYOAtGOsxnDTQ0qP3XI3890Ot3kcPMeDALWlCLmJyfN4AHd6kBT4iLB1nOtirx
sJ682LUV7WXLUKf0l8w+j8l6sXPscARiTgo1JHbhtyQLXuZVTMwSkXETBg0NFC0lwW/3NZU9rXEU
EUwRVhJXTDwjp4TcdcySazqFzdU0D7sM8w9jnJqLDWEpce+xRoRW73q1mbq4dvI2IB0G+DYU2mC2
LGXkufo60SbA7xISQq8p/UTT/7i5AlyCQLeuBY18dIRGgL9UXKUaGTl9In1b6MFoNwNeCsOYTAjO
B5LzIItS8nIhPGsbrBBI+T6jvA3EcB4uuSDiWUpA+X/HC6NbcnT2QGgU6zg5oaLSjzgzlj+iOcWm
hIa3iBlvj+0hFdcsqPTCiTEyviXtPJ9pXJhniPGEpJz4oR0vNUS6R2X52CYqgE+o/OIwHYhhIWzV
g4VIPotqiBYRQITBQuqkcSoxnBfPs5Rrbmgr5uAyJG7gECsX+6Iyf6ufnCljPWqlP2yhRY9xrahQ
Y+cjEXwGTOLnnzEjG2eB9LNmmxatlUClqmw6Z+uGLs2qSEImvyRm6gx6oDZ5Y3dyOVDlnS6/qTIr
jjZMYQpemKkdhZ+GnWP5oRL06s5X332ed6cqYaATpOGCSx5FUSl+4pNe7d/qA5dj3ajDj1woabgm
d/O7E1J/mjp8cCFgt2ai0kh1NPHVEXnfkKn8bMPcQXX1+/wOQk2AzwjE2Ctf1hRodNLm/Q0tZKG+
+A6jsmrEhxCWl/Y14UDEvw70JdQu1iERKt1fbBcloOjYjBS4aE1UXxr8KxNfMDYdo3dX5YnCOkW0
dnbhtcXsxWO441F7ffy7T/9xVu7kB09BCxCKunxxPtIGn+9if2KtxhgxEhZBRDia5PPClkCL/lvz
ES6gXQm92hgEz6ZCbaSGfn2Rb7oBO9DxwOAO/Fs+SlUYROOM82JA9p7lTnBVdRn8cNqV7Gwz/0zj
Dyqtxx8EOG+6GZwxMfhnS/PSxbZ/EKznJN33bcet26SaCCzhmBDrYNl1lGtS6Z2SnCnYmfinlkSJ
iGlmdbCSDoe6DREukbnKaz/55spprtZz66zJI7izc8aw+W1IHBm7LFNv1FdBsVkxeP7EBR0Y6s4p
lyb64L515QsDOAyW1DLKr5tx5fvi6axwpf9pru8i+w4/9zR5QUkgFhLJE8ZGt85mfUA5dd1lQGi6
Y58RL0s22eg54uZVRstaRbUeYwNlVufQ4qO9JvHueZjLbCA1PacKPR3b4RcAUzth0yMt7hOIBHTs
Cx83v1QtWHfQZrK8qHupt1U2NAnb+JyzDNbgIlRFoJ4+GvouJzplJo02FdJW4b1W/ZSdvJcwvpAa
ORMkEGT1eK1E4YT7R3DtU0HHbMapnasm1TI3/Bv/I++s3AiqVtaioev6a78ioqpk4+FE4S3yi/RL
Poc53cDeLRTUG/aqRqyOhoGz97ap1crk+NbNlcHH8mbEamTytjHAQi2/Nqp+EXVygAJgt5Xkl6bZ
iQyWZxNUZ2hFDxxZse4dmse56oeuB5Z6oNsLRrJt4iOSrjwo5qhV20o6F9xBkB4a6FXPu8PW9Hii
AKGj52mCc6dFS/6kaT1lzt0bQKL8h6rcZ3LCAkQn7vqweneHf+r5DkC9TX436VZkW7I/5lOR4AsI
JwD7DRXQGC1a4vBD4NPfoAu4x9nag1dzASZaQb8h0F/KN2yBqy1MC4JcNR6CkDvT7YJ/o770DXOM
p1hQ9L8hH65gFc4xf7StAr2fgBVF6sF0A3bkn82EgaXMnG3ZTsaepYx5d/03q5AVHk9efCFe67IS
+SLfbLsm4KdfAKy/P19WPftARuro9tvWSeaSboIcKWLzRwqElYa+Q3FvPODF1ImefgBFXvt5FShi
CHq2uupA6+D7tfC9exO+HArPQRpPGbs0t/ZUSMvDMeMG+hLvtZmpNlmld3qqPLLXNhqSUlIVi3PO
ORqeWP41QjaE4hV27vPGlHtKpa+fUGdpfr3Cyr55RKAoBzD6xENYCjdVnoBK2fstuRoIxSKI18dQ
E2ixc/qCiAbz+CCTPQBs8RXv+J0mgrNG4zctyWFV6fZZ+TK+NOMI9+/0jEBKRcFDUvmswycKJeB/
wK4sAJuoQwwmiQnt5S3/w0mgWZn+FIpAl7pEQqgdKRId9mzutYmAcv2QGBe7yOcEM3RacB3HenNb
6hIGb5qjRjNyO/bfKmKUIKr4XO2obi5lS9j26XGQTIfYS5IbXfqlmczpob4AEDc8KeTl6Abr9Sd2
6WJTF3pLZR4k5XSMxXhIWEN6a6BsaKdlAUzTszaBFX8Z0rYG8yZ//vFY1a354yl4my46SyQsjmhL
8frjaw1GXXOIRE37r7PeydEKYwKxsk8Ac4elT1JFJHAF+x/6bpnrmiefuesEzVPaCJWNkcRvcNbk
NyS7ZZWIzv55PqKPAA/4mu6vaqnQYPkbfqvGuirPEFAiOGMMJtjQpvfG18gxnBKixfyA4tOOFSw8
xhhQj3wOSafGMCDO5QP5vjFIozT18ITQ7NR9d6Ztfd0wXYf1NMDE96TR+E8r/awb7VUlwQ/T2MfC
2M1SxGbXw/jSQmfkAdoW1IDsR2a1ufhoAy7vzK45Cxsf4BI9WjJ808UofC0SYUt6Xf59n/TeKMWX
6H3R4kwoCP95TW3TJk6p0rXyZtHRvs0zVqnAo6taEMCzP6wjDzsRfQJUegQD2r0GmDJ9ynae58Vx
mn4ht/8+gpZQYoWkudc/C42bLo9kk93Ba3lnhwQhz2J/PuqRHC3cequbpkRgD2XxGB+NPOwH/3tB
tDHgcWyS+ikg0NjzS9XypnHcUmo/Jaut9PSDbTK5UejFVH4wXOpfkJNWRufMK8b7nprKuFuw290h
o4Uazo4/bKPNHGD06PfL8j249ovcViEIShEfHLKcj9BiSULbhP/9oCh/4H9wRDiskrRha6qgLOeX
RSn475DIFpJRQNDxk+7eSE+UpNDYytPVPt5lf/MPCZZWjsBixwX76CEj6i8OBsySUHgx4R8ZsrcF
ULLxblBwgoELidwuAZt8vBl51e+jivf4zfArcptVeoPoG5dsgCOZfhMM8MQo/oV5QKC579aMU2sE
JbBkTUT23/ObJMecEwRFVfFnEb6oQVNZ7Spx65iiVkVdJeR/HLAeGsLToIdkfcSCtcIYKQYDRT2y
7ClHZuj9xuy1wfAl5fcyyOdDAW7+MNBjjNZNizJmFvtFGzCmCSjhTJzkkqnWY5Mh33MDXOUsLoiL
5y3VLgwr5t+OsDqp1OIj1tC5EmCnu+pWRHg7eejgo8wQHx+ilSXSuHOPjuorywtwYx2Hfn47YZq3
W+e6Ievpzt53JTAEElD0Ht8hnC7N09nql2StsppfO5zaAfdV/TYNRb1sEPaT7lU5mWVISv5R5gT8
ijWXywto4F9lTfo21KZfk6197l/RZhsOq5WTeufqtqKjjbozYP0UoPpYiW8QI4bvRm5lKv5WeBMf
1c8r0cklLwBGJ7Nmpo4LmXtodXEH4ISnAhn2UDYKPEn3TIo4cf27IlrwOkIfr3pAvzapSSzT8Pu1
TJwfVHzN1QIBJoJ18wagLGtwPxOUvbi6T4vBm9Uq388cSfOFGueJN9fiPwQYBh6L39Y0m+XO/qhH
6V2GH9nm3WatFexUc8ofMBEYDW93B32A3WjVxNeHvWc0fVtsaQjKduv+LpM4sGBXepYU2EWB+Crv
dRHW1Ynu2kKXLqISfobsU12PUEAw5jQhXS4DpsF5WbfcL6DYeDMOlzJB2wy7BX54aF84VTv1EtqS
TfFIJxc3sfkcciVjIGhbW5UTd4Phq11nZSqM4LiCkcga5jyIxtoETnhuL1liVfnu+9rRMMEFYkn4
iFr+fgGFe3wuPyEb2zGHhtZXGFQdWDnxelClYeHZjdAVjmvVF/EE502oiWqpjBrAxlrxrVMzJbhX
4s1mnimrTItXp/iLRScOpPyJu1Ec6AgFLGwvafI0lgteQgqNIGg4DcTmVYu+kNAolm7P9VvIrgxL
OeBV6S408wDHHtACyviZZMIMLQ8cglDGFHrrnrf0Vze3Z4aKcU2satoSXl81GeVU7zBJ6rivnfaG
dSwdwlOX8b036RUHFtFNkGsQke3P1qZGrpk2q4x7bNIYDVYm08RLQox6nqjXygMV08qa2T2LaUJy
8d9FPJX3h2MqcCpRyCTVZ4vV7kP+lqzj39LJ00NKdwKpgC+nMpRS9Y8knK68aReC7Nbc2xzySy8j
P9V4yBDaiI8h19I9EACD1St5iJIBNqG4vxSrkVuZxENh4an6ekMXyoAeX5/hyeQhOdkErPr0QIa6
seGGSjBniV7kh2HkcWMALN1IL3YTCyr4GWlCvn8+csMyxaWFDjKOZVJBHU0AWncLuakOFulaNcLD
h+Pzy6M9ZYPM36qKa0ZjzAhF9p1WgisKGsCWUEVwq4GaTbV2S8UfS6swuqqme1rpRrAgzkVjS0mB
Qg+SVe86FLh7jYMZ/XS73xS0doNQE1hiSq6cli9cwWLuLcvwA6nIXQkKhvUbgWsCiHd1CQbrT/az
Xyw489nyhTkJfAAgafzIRXA2v5kuuqnzPbx5ykQQsAMKYZqXEy3OgLwyta33U1zR00bJbPRdw7D8
6+MYZePMTX4u1TOSHdUr7751acjDtqrk4zNBxE4BrOL3yzMYODtusmtAu3Tcc4vX08xLjadOvfwE
PzJ/5l08MvVPUV+IE30Kanuaqw0M1eDn43Z3HHS+//z4iXdBIfgrEqztapJmH5wpfviwq+SFYP4a
H/bV9eJKK3bvS+OpFMStRcUzJAtTLpLLEcLnDVL9hPQEsleK5o10xtpF0ITVGjc0yEZrBJFGCFaV
2b3x01MYRGqAShBmdeIEOZ8mxo1wTqauhYiCd0gA9OkhTG6sT45sy0FlSkvJKQ9mptxaiOSPmU1N
CGYaMMmEJr+aDy8O0lbLBb/iw2a8DEpD/VUXN/VTlILveiIxydMc0Q4mcQBe/3ltMyAjtuG/dT0+
FJgEBqvzLbK1TjlnwMbV88k32MdYIybmFE8ebUDFTx4suDopGswZnDnshXXHRrLTAJ5jbCgkzoIJ
Xa1aw3gDcylOTVzJOQ/M1rF8JfOyDkY7gP+Nbs5wq1fjCV1Avt0RxxbPWngqCuVUFUMq6o4/EiNh
pqaEqKPuX53N2oYdySOvy8PV+P0QwsPh2UHxEdCr0BOUD4QlkVu5APPkanE2ok5K6FGdbl00gr30
ACNiKUQeNH1gYPgcfduYs30aCucYimCV34mKjrjwBms1aZ4ZwOiFiUo6K+jnhs3YpUTZmazZyzNv
o7p8/tp61YS4IYfUPMvYqkKqvL/54OOCbP0911yw4kJ23iYPRaT4NyYJR1sVhlAfyc67jvcdsNEr
9AEPa10Q5dT0DHM3xsKCJnaIdFncAT31DtrEneN/Djg/k6KOB5QgSf61JVIImRr2aA3bBC1XgU0m
K747jMQDPVTBF9UCx5AeKtZYT/jx2uUUhYDs06cXcixeRx4CyrwOkpAxyuVmC5xmZNQgmgoGgcHW
/XJ5XbxL9lM0gFCkK6XZPX68aHHYCLV4qJoCWJMtkPU0wbV9DzBcipuv5AwZj9ZXvZ3ocUCD8iG8
h9I2kUNy0csBFJ947FcpnmrP4y/B06XBcBaQCd97foJVKP0eEhxJyYxEZoPvD+rG0rQz3se1ZEjT
t3hrZ/IefpXkvAlewK7Mi+Xu77yojM0E3ZVs5jP22AeLTN0556ilz02+M417JpM1ySeoe2AhnuWW
6oeHLCZBeEg8uE/zDZrlzre81hJToTHKE4fnNsAb2ak/A6TmTs5RixfD3zVGWKhHcayNsAz9YGwu
wNPIt+4nJICJWOBXnKgPsppu46P2dPSXvbhs+6C6B4y3IdBYx3J9NA9quFtSLdmrrIHQrGP3Zdpb
3fB+D9d7mUIpO0H7cPVB9vSZmEeU/9C2iyn5ufju1fdBopvSaLUFasCB24hIG4ofyKES1HH1zqI0
mO4YmXbB2CYm4K5upzjJdNm8ifoMuDM+4W1Yv0ig6RcMtGz+DgqpGa1nejJx/FvMPS3t4cuv1FAq
dFTNwEVSuDWwB4zeQYQ1Xz6h1kh3z+BEN7WWDjIaI5WrUP18Zn7twMP8qlIMIsF1Ap/3jpJ9/rOu
sPDUZClRzszlWQKyCzUElemC1aJb+rXbz9Ze3QPXt7uWuBtdwPpkuRlHFszZBxlP0iQ6e9KnD9sd
EvIUEoyzgYGusbFIAGr8ZelCjMeVJ6l2fXUe8/dlPMVf9AcFgwItpLKWCJe1uUuStNt+QBuKsowD
6UCln7umKR28tH8qvuitZ3kRFBx2CDlqLCwFaRYYWTVmTzrKQyKe+uogK5eS2RcLG8W/w/uxr0EI
tmWXRd1tcguaLGXdh6K5V+Hgjb5sgVartAjZEcSD2TiK42riDEnjTPs69kLxEkvOKuGtU5lsnfm5
tMFy/RRE/B5id1du3auI4XuyoZCorhV2uy5LPtDc1BK+Q3az+/Y2o0nZQxQGJ4IJ9kXg0glCvIkW
PYhAt60f3GTGye/HFdzdlwf/VAjYlGlB+9+nBefr1Pq0dOy42rLD/USddBhLxRTru92PDBaHWOq6
CC/XJboBGm5KgDfxW75gaAyOMi2+VyAp9BEWeE+6zqBqgs+NU1oM10IoHw3FGXCMQLd9Jf1XCvF9
8RViRaZcuBe87QU3rc4hkRx0nEmmmLSI/sLOUWEDnP3JzjVv1N8wy9wdrJu//bxUmh7MKLNSjxM1
YkiR9I5FBFYYqvFVXZfm1xNo1Y+o0iqMTOz4XM9KRF4GVpVyetbxIgzHXTdJYpJUBpyKFTAqHp+x
ONJeVpeLLECCPzmedmeO/l6bLHloJtltuPjnLdUMFW3SKaI0YuXlW2EJVoQj20DYYlfBTa/3KXJ6
LUn9Vn/KVWGs6ALP4fIkttssY1C1d8Emg7rW7GiT3o6124GyVcyr4TeeHmXwLD+xgXjY5CPi5SCB
Ugu6BVO1obET+sOfTpZ8Qc6K4m6ku+sAE5db6+OPNNC+kHiRdJuLbC7eL4jA4VWoDPDQbNJOvxUW
ysNfnMx9vmBzmqSrNXIcNB6wiGRypLHqXAzV8UTTb0eorZI77Db4J80h9dvdD/UUliuxVjJ7//xy
jWCW+gim/hE4cqLE4JK6B5Emm/5JlKn9kTAM3hRO8gq0K2gJZcegmP4fCxwLguG47kzYUSDp5pbS
KhG75bK41i1tBZfGk9iTDA2ehrTOHPUYpLc3v6gxlUt0kP5+QBz3GBypG10vWQMgxNVtAmbAClL1
EIoM5L9gy8TNdV3fzWxGNysVycEAogKUcN2DHd7eJU4TE5d0W1ygw/NfcjFV0WPf1J6oGNa8V7Hq
dXhbLPCA8TpKSC8zl4xUgrWDMtagipypnEiLhGey6zhl+7KaDTvspslyTbb4gwvEJLTyjPjVWXBi
lepT6sYABTP1Z6uMB2DarrOBGAHtGdjxy0+MGVTDlM1K022aRMFEpLlFDuAXjPi0mkRtKpIA8Ah9
+i8mciM38HZOT7gXbKrPymd9PGdXGp5ThYdjQM/sE8GUsESeISMfSbDffX0Su5kWD3+Ygga0sgbp
cu91UCF2zdDfciFAkRqHbaF8TF8NRBIbGKrmP1F+tYKX+qiIb1cRVBjfwcK6C1qfILkD7VBCc+L4
I/zZyt+y1znIRTleACt3oxxMXYF+ZPrJoHeA7yF/1TIgivf1ILoI/NlucRjRuNWHE9c9UsEa3X5u
oKfkk6Esn1zLTsYUqaRlkhM63DHMr6G7efHjTV+OIZfwv2xmRkZldqHFd33Kh0HF10xNJIN5h8gD
xxwJva7K80ixRguidzS1iH273csDT5gBlpqHRA4awkFRFmtHLXmJ7enaW5Zp4/BTwsKerjXTu8uG
yYLuRyqa1HlK2oQvzAcT775GQjQOUuIyJBLdBbhOXgpYnuGy7HLnx/aFmnSs2j41v77EyABySD9p
dQoodh01rAVVGcRY6D3uwXxxGcXuyTrVIapJZuYhHRgLt13hZK50NCgLHUBuZszgki7JVz6msPrx
v776aF8nCqHKjpwoS2vEyNRjahqjRYEQMLIHgAGILxbixM0e3tsMEjLbo7kO5tc42bw6b+Ova1YU
NTvdYW4MDtAkOa4hz7nazGoID9cg+eCaIAMEVgQm10jhsV7/IWCdldIAwFvBARLKPMjR/bK89IIJ
2UWXGEqJWI8hTGNeyYHCsrF5Ord8BWxkho65grcj4/wi4+f04aPn72+nl1/iUbQBzhbQtS2FqDtN
Bfe4gZF6NC1CRe7SwyzByd/x3QtDOgk5WcdV93oiLLalGg8OgNsDucE4PD4k3+nJZh0J41n87v1S
HWl52giGFTnBaJsGvMuLiSkNXSETgGEhKvEXCcqqNYdI+/OdNzwt9VanqGBAzIFdAyXKg0LlQkTs
cCj7qn3Pvvm/gEJ15eDSKKLEeYMep/L554oqDpgGCJoChwutlRz0/n+36JKnzF5Rr/Gy3qYhxcWA
KJgW2q4lm/5kMTaGVvo1Zh79FsdscRaSI/Ho3DW4wxo/7WW18UyqTcQWXbNFxz33Kbk25K7X6SWu
or/OyOiQcj1hudWGqQ9CH6HQFzpEO8N8SM/B16Rn0cF8mWxbqp5gOFgsfh1YUF+dnpp/58K35Bwx
vXwipobx602NskVxm7YenHs1MCOGjHA9po3z9rHl4sXxFGTKQVn0go62QY3JP7SpqGXEgiZR+LWQ
yQMuDM5wAHXixqL+WTl4TSuowh9W4WDc81t9QO5+M3HrbMl8dlzqIO66aOnavA5jeOCR6vDjSfUd
N+JdYKFxkOEZVFwaVNRRzcETvYJmuqiKZZ/EikkYUbipk03mqvhW0WqZ7sbhvaZVM4ikbydQCV3a
FGldcGCMnZrvtpjMAmeoTMVFBmCL6S7mCdrZQkGAVYUg4wq3SRhq4lZv38AKKO+ymtJbvIISTpxF
eLh3fY3my+v+wgrtHTucbhgd4vsIjEsfU8E0nu9L9Egm3QmIiaxEhxVshkR8Pq3n9AkE54BEmHpG
1oSf2nypaEsJWBkB+k95yK3KeYJN96u5og3xMQmgY3XAJTuSefTSkgDNkBEIqfdtRU1UEJjTqiIB
GLx4Tt8n5W/wl2DRtP/kym3UP6n1oe/I8DaJKoPD+ltqmtOvHToem12pwHrxF49S4HpmqYDe7mgY
hpOpfC0jd8RyuYY/RorVJ1eiIeQ0RSLSPkUMswEWUer7Kf5bNix9RdngM8Kz4D4SeNLrM82aMZ4R
3Q/WoyCZqs7Ys2VuooDV9owepN8sSHoFg7/CVRvfX6iICqVB7/SbFqw2Yjp52nQ0z6NMnVJ9naHn
Fod1ooqrg+VydqBU0AvJWSPEbl+4B+UXSVqQdSUH905VoPUBKfyaHjudvQTcIAGVav7FzzUJZJED
eaEjAziD4ZY0w1JKInizdHUWC7ZjxLpqazBzt/aUk70mJZOwpyehgq9OlBKppgZ/9LeC4s3AKaD1
QyZMr+IDVWRIAJAuG7Ll+aGTsywa978UzRxAFkobkdsLLTZW6t/R5FLta59xVGko2cpA6Zrrnxy+
qGKa1pMP/3h/deUXx46OQxKVBrva2cTX0UG6Gqhy8x+MbI9P/7ZlszQT17o0eW1Vocrb/VH3DZGE
tJl7vNEDZDqdySlojuz+aueIxH9C708Q42jDWNPTE4sHDJobdli4emVz1yVs10G8VWExoG09PJNx
9gW8cMXBetbfoL1EQvfDi421mQv+ywJMtHeANgS4jKCrrbqkOLavd9mIRjU5UFQ2P8+Z23E5nv72
ezRIl4IveX6Dc/V5Gek0DVqjpxVMCsgon1Sk8J/kbaLw2jOnlOEy3PjRdyMhTxvW/aUwM5Ngacpt
C87bAtZqnuS5zECtz9gBSr7j03ERZ70d/eYKs3ssqdO2O42yan6u9+Sd0nJzPIYrfSXSsHSH4sn3
ZGGjbX7yovjAw2aTunJqKWL0j0LC8uCyjZU1PoY3tZnQIMy10UXPxlAVgz3gc0Dei9vVeR7lYQ9S
1/cgoayuzKNIaCZqhnyPLhmy1Flgpq6A/TfS2nEjUc5d3CWFKwwuqOZpSMq0k5YOAGmCnAkhe4OB
snpv8Mo6Bu0FsIfMQIRb/zIqP1qsKoUQiYG/3oKT0BXuE5O78mSEyGGPsMRQ4EMxRyzFDTg6m6yF
iZ7ykjcmQo4IqEmZjKhmq204fgNNze5/FwSAg/X3UPMFwYdu/iN0BaqoZ30DLpc6nX3le4PxH+/g
oohGE8vWRUHEeNDXjylOrT/x/Lv2gWNvDQ3iNBxVD8xhAl3YYEwKC4yP1vrq9eD+h3bJray89kW+
ZRKwzyuDPPknY9gbrlsyeecgXGxS2noVFV7+csCp1njJ1JdnKg1ic06cNYivCSPD71UJ6fCcqD8l
l9+sY/etOOwP6oxZPxz2fm/SR2M7vmx3oUeWHVwow7DPwKRMCtiaJZTktsBB8mfXWvG8WRTD8k4O
0N3cQ91956Jm61F0fVWimoNVelBMZl9XK6SlC7tMsPA2y9Yb1n/7xJRa30blpcgp5frSiSZJ0JiM
GKXElaIDJzojNK6y6NOnmMlf7pVKTX7z3ItItFu3odDkV29qHx9K8pcua0Q9N93zY3Mr1uC0x6gE
RRPRo4CQFIomUbAuzvmm47arKsD9MTT4Bdn5ZZwJFJgdE8Ljqd188I9nmWeymY5RKB6uqZLk/8Ya
iXJJTx/ukqBfhHdrSb0phM0fU3a4CBiTIJKMeJUOtib/Xw99XeZErV4OPz7j90BgiA+UeuDXvaSE
9FkZC7XGNjY7rspCPk5d+va40Z06ORhwqTi17icJP9v+I5GkC4Jw2sZevgUXsZZfqV5aA0cCuiry
92km8hlz9fRhIoqP/3/ap0+lwlP62DpxCY7et3IHcqauh2YIst9IcIvIGxE50GDzYBKtGpl9XfFg
C9DxXtzJs3tvNmMrEIa2KCHYIT7QyG5+fa7LR88NC3RqI+FcKHZrqBr6i19H/5yTwGEPRl1rEzgs
d1Q9TyAMflyZduiNAvuDPXyBxKeMYmVWzB8+e7QnOwUCI12I1X2+aAze4q4XGViOvJdWji9DgRUy
T2HeuGl5TC7USCGMTf7D4iulX1WaHcjr/M8H4dBmNOZRdwdPICDNFMeC5dYDZG2zW4+aXc+SbYtT
aCQRc++8ZIEo8r0gmOWxE1siiTuxv0889+QcPAHKk5EY/LfZhkB0iPellMujRZ0yXOdOPKyEX5fx
eXb4Fhy+hAV5QI0IgsT87nK20Rs0SolGtbJ4NK4Kx7LMrL56XzddKRiqUw7S2Z6Rev+qZhr8IHj9
r1E2VT6Ufbb/souN+mrl1zNrdiPtKJCG+yGm6I/Hp9lUZtqx+620A6XkyK1zc0+mYJaoWZ4UeFYy
epXK8R1nlvJHFT+RPssExVmbqNZJZIRgtEKAJL5qfOm8C+wTXvI+r2NHPmO3yCyCpIBe+og2kthY
hSAdpnLUXbp28lXqM+6P9cWHUQTVgK0JJpOQaL8dtY9ujfiScdDyDEA/9gTYRy6GRlAvbe5+KhfU
rFafSo7jNrhTotyOoO9D6kzGc4lXDRYUzbOSBChmUQWwyRiebS28JTqrjm0/9xsPbeZP+20i5M4g
pVjs+ZnI2qlknvYPM6PXv8nhbi2EU3HxDZ2ChnSZxkeV923inzw2LvJg3sfprQVBK00Jxq525nBf
ew3LvXU6CanHWSEbGkEJKpf4eDOkavgv6buv3hCvyLALyb9LldoWUNgq/fcflPout0fUA+lgi53M
hwKkF89AJ3cJWVQ5IOk2wK+vZAloYKM/ltDVCLJXLKIRlwjBh3hJdMUXeEaF40Ty6J38fCaFL7N8
rSuWlFX7zGp+fm6ahyp27YGdINua7q4GDAfn+C0tH286oqbWffxbDqHOSmrkhw4LTtxmV4L3LT/p
Mw+lzvpX/o/gn2p36H5/T+ChXXP43pS6v6hHfuBgE89ciiPXfr68amihzI3p5d9xODQArdTMlaOe
CjbC9ocB/GXdSnPha747md/0D2CdKSDNWyJa74eWxGiPe9n2JQ8T/d9OSTfgHI8qxQN6ibsVA8jF
40ZyiIQqxuMgYY66F1FyNjGRrFbBIl5bXG741X0XsUV+P2pbBYctYlaGoYXSw3VM0VdCQ85CBILh
NMnq3c4kmkIFWgjtdarB3lkDkZpPVOL6BCqDCt9uOEQAhWjABuDoKPV/DQS6416B6bQ2ansq8tR7
C+SMxH6kODUzMhXPq/xndeAZJ+h3Ta3bZl9ZqC+Rq0+lp8cdXsGh4cL5pkSWUFAB3XdaRzm9mAr0
Li5Pa6ClUKpVNVVe5v2z7pHuehXVAmZs8YJrbZuAJJf6Lfu0k3zET+z9+g6bGXe2uFqRaHaYvOtc
tFK/t2J7roAIFYrl3M4Z4a5A53XqqXf9iFxkbLhopph2Hv41V+P/JNo+knoo5av2LmNxRc+LQxIP
d8IehGbeX2DmgCENOPV4rKtE0PXQ/2RbHrymRFukB+9t9C/7nBrwwlVysaCKRU5vuUurnJW4o8vl
9eNC29K0mDZ1eh9/sbHLqbsxWQrPZJ2waESYOfdwyikySq5twhYiRn9mgji6LLkAZYE632M8vazH
2Tw5wtOxtmoZyzbk1foVs1yMfMzwQmK7wsnSxjqdmCmuJH1kNf6UcxAbdAiotwo53HSRBLwA55qz
fD156vFFM6jeOI7Oy7hUfRrBKhjjks/L/4C/vS63Y9UoYb8K8yL8M3KPl27DIT8rBkhemrraqFle
c1ecE2EUk+SbODD5wJmxFc+IblgjskQlU4xThinJ/2T/AzfhDGQPYpRTFfev99xykt02dB9UYq1F
mzNqbICfPk28Qk+ihAGnamBEzeMMLrgi43DxmTi/yXnaLkEuZl1c+5BG245VqkezVsgJU1k6QIsO
6g0Wfo/l76qVQp7hvf8pVnsTs7anjsNkJGHPZUIfCrqTCSm2udWHni82VRaNBpxmWOLpiN/LtL5l
V1IWP/G/2ZwfTsaF/KE01Lux7SjZpAKPh9SBHAipz2aOs+lIeVmzZEvD2pxdBwXEXzafbxXXrS3w
phQs0JW3emz8DEuq9+St3vS02tw9BRh3sPAzwUBCgnxUu+K7G9lZRtUD+qrmdqFdDHm3vyKcfBf3
rPsAy6vadYC4JHMa5/vi84Md/N5yvnag0Cz9IXda+4Yi5XIgoD1e1zNtzVy0KuqNeRagP6117Xe/
G9LU6N5LX2lwoSoMzxGCCO6R/oo5LImKeAeCWl9lBQ7jYTwDItp05owUTKAasyed2SQZlj8gf8DS
OnUF/DmgfeB6TcyJUPbTG1vz/rC5E1z8Q8MH0OirXy+jSWN23jgrqEv5eSt1ZsCbr1wkDzERQn8k
YccnNfGudNNXAOm94T8OCUdIW3Xi4w7nUIEsMRtQx65Fh5qR2d8xHGlIc68k8EZadrLfLm6u0Iud
t6ZmxAy3F5axSNKoWBHA8Jk+vqiNfGYC2e0WpYdLMI8lKQglqbMFj6VjoDIXV9M42Djr9KdI2+KR
u2gjUFoSPN7D4o1YMCNGDeALtKHyEtaueTikuwQ3aQzKArEmx6DkbSC2bgdFmsBRdq7tHymBjhZw
6mSAeY83a7IjjQtHmBW8tG0nMP1ovT9j7uoUCWnML8BiKB2X2NtwpYYLA1BGUN4c2D6g5c3+UaBQ
EtG3z4TZXsWyPCtMXU8L81WpeqyCgGZ632G78CG+pGPf7pxCXWpKAzzeSedjRUsX+2Z26dJHS/PL
giDr9Z4Su/FKVQmztBGxnAs/6ZEko2K3Bt0/5EJRsT4igjoUHxKiIBjqZG1mRlMrnzsn8lyNa8Gi
aurQCQslhBCwDBkXNQj9zzP8634Yvic0ULPyd+bDrd5PBEfRl1L9ILUlhQuFpO0db4K0oEG68uai
LTjp+nnnm0b+JCr5UaUW9qMJGWD6pksCdDsihGEA2pE/uLKizj9B1GJu1rusFjjrhsNbI4XlU7HE
tUTJkRbRuprk+kMY3O4Xv2HI3aVQHD95JSFF+j5uwlth1jhtPZEDSLk/EhzOliqXI9f2QEIb80RW
pyfyFX0xIEfczpwPNEQpyItLc5sZYburib+vSBzVND9zrfIc2ASSeRWOUhRGiB/DoZPX1iHRj0uS
XFW/F5D9ou/SpoyY0IMa2YPDUo+qWtmO45T7Ng1s/gT67rqexMw84dShU289N4+R++MCcxHSATPd
9uw9pG54VGbH8A1paF3mblRMcVpzBR3djRpp5mavTLd8AKgbJ/sLiaFSd1dZUY5DjVqsvrbSBu4i
mRc25oa9tVgq3FhSYiyyB6gxYS6mkcF2b2oyzK/U0AjaU4zdujdxesR1SFqaG2PJg6FD2t8Jd3WZ
mfaugKIEGXzIRkPCIWoUtM9CfbGSJhVsGRK0yNhiWMHejWcl/ceIvhwr9mYBHuyhwfOF/AWGYyCT
vGyqrUqSYrU8pvehwUxH52wnNY8+jkTX5JaxJPzhN6ewdTQA5L4Lp7LzspOrTlhow48AlM4gv6Iy
6nLK/KW115Sl7esxZ/ppLPtLxpZR28Q0uut9HBS8Ynrp0c3GBrjy+zyF5K9EjdT4t9pE/jPy5vtQ
N7P+fYph85hcJTpVFoWriziiZpRWyQL2j4diDBT2gt1tS0kuEneku70DQi90pe7oS7KhO4ISfS3u
H79if6ulvXwtW2oqFJz+U6rU/0UL69xAX8wuwSJtH4AI6JOycreMiK2viW7Hjjl8eGNufrgrG/tm
WafUOeH3Avw1UbbBDfE3l3u/ndGrCYJ5jlFCQRAmNtYjRJYfh2RPpiI7ZdLSGbqDQMF0CBzUvYqE
nxNy1ExQHBetdjmMDF7CjnmYLtrtzu5P5XjtIvlJIdpxSqY/Wv8jgXUMHihJ6mXo6aEKw9+jLPLs
mRzmd12w6QwIb66/uSjPUusxtobHIyUnGOAEH2rb47pqBCTjHmGkDCWPqWVT2fIVp1nb7x6+dgw1
oeg71UjIVBzLGUres3SSjN0ZGJ9xzXwANIpj0C44kUbbuxriPn7jMNp5Z5CttUDfcXSmzMxoR3Tq
7ljObjpNYWSihpO9mFMo/3EnByLjrGyqD/M5/Ax8veAqA516pl5FgmbsB2czZbnumtWSAOHxQekf
1FQZBEMYzDB2A9gZwHjL3dmiBvLQVxtPS+HehY7/eXarUMXJRp/CZBMBQN2OjG9VaHy3XUobBdks
VAOrXWZ2/v7OV3tRrfVPx/2qGCZJF9A1+QxORnqUBSOkzNtAq16Ci+yXchUEKXGxrEOsvhnNzcL0
/s+QE8TobbV9q4hYbvqHPyh8d2iEELIzZQ5czsO5WMwRKCpa9+EOlP/csc7lrrfTr0VVALMEAA7p
co1LyNRWgbzH2+2StTis1VfYyfZK1QChEtNuxgiG4T8jNxDFbEpJSYaStS0F3YWbJbisYKw1hgRm
NPc1TD8QCf1i9PE2R5tntm70IjfosD/C1BCZelktkVy2eLhTmSCPJQxhDw/6lnGNU3dRsC9QAeke
gp9u7KLyR5V6zrmmBAyqXk4xQtY9enEmAf9GhubuznhKnG/WDXsYVexSoGM/0xROQGfEhT/OzGX4
z80CVx5CLzZgj2eDef7GA5vnh8fL0eoHW+pmoTLNQPj2/dnp4N1TnE+2BOC51Vb2MNFkXPGQ1hc9
+8MqYuPXvGmJ2PQyhy3+FWHYIE1yAqDlNy07wfXrvuqFrw6EpUuXl1Fio7G164sFkWK3/mdCZ7Dd
b9XTeZPt9ksNJHX4z5W20L3l0CiqD/HBK1Tu7q0rJBSquOpjiGc62uzbE3d1lKYO4hwqPGFCcsmm
IHJdwlYfNz/QoOeAm4/GQk5Jqws18S7zGuidxpEWbaY4e1/DWoyKupqTVBlEg/y6CiMyBPF9MXpk
CuhxNe1lQKbJ/F7+aV6EeKTtP+oAHPqviD32QyIIqNxVW2YNn0w+CFFYP4Ei3BKAFXEmw7PiQ6os
YUxcqxqlMtwA9xwbn7wqZK/+nsm77Z7f/cR66ajbX7tMMwaEPp75r0cZNbw4IvzCiCFmsi/fK71q
0Ac4V1WDFzyHIMv5g7EluxYP0SLw6id8mNUB89Iwj+HOajjaUwUUGxFmTA1QjuS/DZyQ3icL3xNv
FUf8ZxqmVmel3M0M3THVJ3DD/ZCQ9GbtG85GJYyIKjhRgWwoxMwLlNKfITZBU8weEUZpHVup511I
BeDmzBrkmx+R8+pLUP24y5N/s79Ec7/sJZMIqQLd0/Asw/c3aHd48udKoVrlQk337tp1VdEkwJU9
21qkDmnAQxBLzNwQLNsXc0uoYRBQPS59a+S1wWBK4ZcV648CYNTW/4Le3X+NoCNfyhE5glzxWQdQ
7lFeJPzrjJGg2GvzvKHXBdmqqhr36IHH7s1/DD6fp8ytx5E+/Y1HcLKvWYrGEc9Wc/7riLnqQtaI
e9FQWy7Dga2wpeDKWL0o41ANrrnztu4ryHNS+ZpfcLzZZAr4O07YKB0ZICT/MMrUVgRuIB1KXE8n
vQmsvTlCwRG5kEyGHboI4oPMY9T0uGulWMnPJJd8ZhATqjfUJEl0HrEf5/T8HA0XVgn5T43t+duo
z4QeTrhrlAFEsva/Rl+S2WUMoFxiUXSgR9emj3zg578luUXccO5eu7dIiPsEm7SanlrGZxNGSG8o
APrOGmucxnyaukL8c2iOAUXT40O/FutVqt5ImJzicACNd8Z1LqoRPBjja/oZ9AIui9EOeonk8p6a
ChbnV+lzWltc+5lFEQnr+OtpnQZ5LjmAnaQuoeW/sq6PkWEh4cqDe8DC0j5AFKjQZTKqXDoArWLO
qmvGr+3gbgzOimxlHj0XlRrVYZhERX2lmNG9trXPygLcZQD5U5tMpE8WwYvnfzuvJn2PBha0m70f
ayS08wHWAAp/8oMy1IFeeSbry7IErVKY/lTJj0NbJLQ1uT1Dv+cX5woXqBkQfutLYibdyOcvXDbI
NhigSjFETScFnBGSZ8b18ZcoNkV2452+q+DDxtz/V8Zemk2DWyznWUGfEeh9SLlngmWiWc7glPHN
6W6tfAEAxQJyJIkTsyZQFetA9XPaxznCm18v72o+/NC/Y3IkEd/SALdN7M19DGlqsJNyes3ZnwkK
hQDjwAp/Wn49GGYEE3J5JYqyyzBlynrmeUuoWG1J/cvmq7nVrIdS4CNZ8MKyUfGyH24xYcwDPJyJ
4qhI2rUH0pp2WeEi2EFvD6JTmOol3bTHjtcTXXMQYd2jltg14CBzYWw+SrnGfayuiu4lFap8LgTq
BkPgqXXBOmVVqN22ZNBvksCQ/jxCya6PYyDkGKlyYIToBBJVb3t9Y7QU2D+Bq7RRDArNN4BDar/M
tLiuQdgl819DWxRzWC3y9Ljsfpawyb+m8bcBT5nNdIUJdvFpLUdWyJ252QJUGiZHU8ylbMTyW+5E
+uyg9jKCy7XLeJ4PrZFzFkwE3LXjpiUsMoIKwHDJUa2Oiea3OZ5Kh6yhREy3waQTpRunFZPFdBB9
h0FqjgOXpAXxiXVlvJvSwJ/qPeF/UfJWOlsMWE3NsgKF+drFJkWfteAAciWvVGOeGEmPDeeKNaTZ
8nqN579GNah1O+BoT7zAjSdRSUKmySc/nrb8VnKS/VL+ZKbTIpcyMr3ipSZTJwdwcLQRcTBJ32I7
yarcbFXKx3Z6aIRiH2aMpITw3QOFTUj9R0rJxakJPkiiplB+y22C9/cvcdpc3oop4jFTp/C/ZDhE
6i3QO2IGXz1k/j0OMAtZrdHI4HPhKvrBgVc40vBfcWvdfc93ByRDxzDfmV9xCTWujqFZwuY+5hw6
O0NbnzGcTVlMe+1bSr0VX/6RglTix2VCY3K8Y3n2PMV3BgKNzkN7jY6UWptx6oqlfrcVOW+gYn0S
oBb+x816vW47g5wJhzcF/YbjkAIUPz4XjoRLgDEfeEkfSagPkPsQlFMtHe1CHEervMT/3qDQwh18
JqolSlfXkHPepTnmtTzmERU69ecPc0IPdb7/Y0ZMgRpkXCvT/qN9x/58wCPJe0jV+G5lG3HjSdiq
6JsLqbPtGTkdmB+694ExqrfvkE1TG90Xv/oTqPFAZW0s9dT7MRUGBomEFAx2r5gIZ0pYWAGTYaVw
7aJ97pQD8Va0QFR7rZFOFLE2cAPtFD3nxClzjSSMnbko/zj00sBIVmAC857QPn//FWnmn8OSCdH3
MjPNAJiuVCYm5g9dnxN9ZjIm7ESO/nkEjbprvI63ZWKpXBYIc5qFf39sdOTtpJr8EdUcncNlZSVe
V9zH34xWLsbDOP+TKAW3UzYTBz/9qGQUKtEGiQpCHoRhzsgT8hVP7PZ8hd5/rjfsTi1BAYDS08bT
QEzspX2Rsk+Yq+1oe1EaxwfiDZ4TFZejzABOK7kIhqBiogbWLDbGKGVqxauAVmGLlVaesdjDm2MZ
dMkZgg311YfZDDD9wvqkMHQ3NPEFKBV/sHMETFMbozk8Rf3hYVeK+x1dGUchfiP2MgN1hDImmuCK
LO7ogJmo+zhHTqqjgdejLx985TTc6AgD5+0bnypD4qV03P2iJU8Yj44Z4bQu9nR4X+UbFT3bf9XH
VatMwY597d8YbMQTSIHugdC8JWwSPh8LQZYBJl/5GGtO2wFBZcdV4bk81hs6cNIVWo2dlOcVj170
YX+4eblmpzD+v2IJyGeL6ah33vF6SX+wtyGfzDvHtlaUCcLGXH+dmesk1HBSqdiRKxG828cVcz2W
kIlm1EV3hgkzsQiAZ1QG7rw0czjwXZ3GH6eGgzCgOD8bRit49EY+h4jp7u5yAVRJwC1UdSxibEKL
6J5B+NJADqVyQ1AZ30eAaAVUorvyvO+kgAFOVNTzk20SVpCwjeIqn05NIz1yWbDlKJcrJubZk0y2
JA1MlwaOVQvtsQZEFqN8lrBybo9AJ4mHpYsHONoQWGoWxaN/AAeItw6T41YsyxWTNrEOSl6O0uME
VMGA1f2VUZYEzFTE2XnFsWgHTbWk4EkPfED0K+Vd0GTqQHGBhskOyNk2w50F/sU5PSb1bfk6TCww
GEwfvJLPejBoPP+t4y4GjmDc0TwnejVxlU61VhDUKoq/TiV9DLP2BPzlMNSmj9UYZ7CJaTibYmqy
Kx1s2iIpw7dsl5bUPTXUEuWmmuR7YXAVXv6iigVwQS3g3n+I6Ai680pQ/jbtRH/F1AKZN/t1PsFQ
GAlvqAN6CidekWGX26OYiimc/joNV+OJVDhcwvijgYtsb2FU9K7oUV8psVgP5XDfQ8814vpZrc1A
R5awKe0LSkXQTdJJBABBuVkMcI/6iSiM4S6C35LQ669Y8/28D0dWNEoovkvphOFVYlSlYYdfqGsq
9Gd1UCJx7fQwDozR9mxsHlAWTT3ofjGvAvfq1SFOritByuk49IUhq3dxYte4uqZ1pr5wY3oylMmQ
RCzy0JSUQtQZZJT0Y6cFPxF1ApaDSzAeDO55PRPHs1hmEgt18Rwt0dwx8CRbk1HkyEwom53V+iBL
uHdcvBaHmqlV6PNt6jBLsID6vraQ4xl4P0A3D4dYKKKoYQeFlAlUSwRCa1qKZkUu0sjcbC3MaQSB
UrjZq1UqkvbAdfToXmsA2/wDiX94wM9D02pSLL0XAhjCeC6wMJCDFSKBTD98XnWDzEeJnZa/ZDao
lgArraF4aiW/VqNEhBZJ1l4KAt3jYViOyX6u6G7Q/gptdtPe1+T82jVkrlxxUWL/ryDKcCtKvcjH
vscH7Wy7Vem0LuSspMqxOv+SPp7XSi2Y3nWYK7VXJOw76hRto5/O6VJcWchrEHwD4eiIAcH/1SnY
Wnp0uigDEs78er+DKGzoyldCVvw0B0je8GS/848Uo05HhdP4EQHKCQLjcdmGFb0IGFbrynDbXvN/
enorgdaFNUoIdJWpuFtgJkffCa0AiD7qmIHiIOj+iFYYPcmwTAurlgnmJQF0rO9/tpoHxV88FiVa
1qaJlII4YO6Dnwb1jajIZFxsBtjvnl9mdEYaWsnsGevdkYA8iZQeOZi648nuc2j50R0OTVduneKI
l7L9Pa7Wytph6wHx48+ZlXSGRNh6CSkRrDCpBugYOPcxFdAHjA07VeqrOWc4f5T0m+CZ5MtEVlT4
p08q2xjC0OHEaTssgq8Hv4Nba/OyhdyFmSi54QmIzGa8KhtpLx6FVfr056HzWlzaAmAvn6K4tyKv
+wZEGZDQnItvKhlQWgQUzWIfZ1eYajXNcBQNZFEg4vIMt7PPrkzlRNa1N+w9PCg7rvogh/d1gjvK
fJV5yQGoRpTV1mL2WuIm5Rpa5+c+k6vJqPq6KWRto17rTWT+NNJaxjZ5yUy9g1UwU3SApTAZ/mwi
dom4BcsohbJfsWD3KLjdyhurUpSaxG79XyjOIUor+dCpD9UKQGaGLwc/3ZSw/tceBVyPRwDG73yc
IB0KM2GBHAvzbUy/Zy0d+SrboroiegVUjadp/4mtqbQiN238v+aGG7t7riu7psyeGwrU6a2OlRP1
bWVyTvLFT3jP/MUgLca0FrPBgrL3kYdMw9Vw5Rm72qcIryWYcn4Mae0C6LJH3vxqrUenRcAD+xk2
YJNPvPIELUHxMtNZ2VMZbS0Qan0Z8bllEeEKMvHEqWPjPpRRy7UCQEz5Yw9G9g99J6V9FPv4sclr
4lY6cZgZsG4CxzlF1RqRWLYgwGt+wqi6amU1jai/XOHDq1QH8mCmPW/VhTXZqnPBjhWVj+qziPt8
tsT/9W2brf04On7BcXXHy89e59hqpdFxiFNfWv/mi/TsDUUjI3YXqHYDv3LsuoCtjvbIM12LCGTR
s7ws26U3qJX0GZ3kZF+3AMuem/XZBa8VRFJa9Nvvs1iT6s2e3A6j4eZszqBOWkHqeG9mKvaDC6e/
LNaMNgBHXiO4sPHjCV8C6TNglnft2DTQdlYvuzKhBu5KsSx+MejkUjCnjca3jpouMs5yq4Gzm0Rv
h1BNPRKpN7fiivFA+u/I37MQOPB+NNf/yoNGDv/vZat/jDMSVrm12ozhzzgAEiqsWcnFVcruR0yL
ddldVbtqoBPChu2Z/RyLfU20SbmKvXx+qNlsh2vYnPVwB5HHreMdkBTLbfHxAitHr7Cs62tx9u+Z
dduOssxcspvvyOFItTEPiRy46N6lVpCCogPgyi5Ry2Grj6ILqu9iita8FsHqc2Vz7X3fc5Tg+eTV
hx26JJvY3I8A8gZxIp+3NAyJvC6JkToffr1LuRLFf6l0jKa+JD4U8DVnalSwUanXCPD9RmvuVQ/Y
2mcm1Gv9Uf0JIl2LT8VARbFhmirGKP5EayBfYvWlm9vMfaS6pTvJcrsE2rmMZ10c7mB5YpoDa9ql
a7eoY1nl3FZmHSosSvp5lJim/LY7xMrOTLSciWLyyjnJHpafMG4yUj/PwofOO2DFbfeK5km8hYsG
Olty6G7GqkzPKlt4kak+isl4D8qOmgv+SqhafRos0PBw46HEkveMYeh/IA+K9JJFSD5tDXE8jH03
jRI10EYOLK97e9KHe/cWexzaEkFK/Hbqhftkr5rs5m08h/MgrgBietHyV1eVwPuRBFgb9+KmucJu
5iYNdMB5mGAho0EBSFnhdCJ4cW4EolULle0QRlkI8EqNu36QQ3tmqfbXIYld/7YhpJMVYUMW6E/D
W3gKfSnUu6ikYiJ4LmEc1+aGp0Ynt9Ik9ddxLeaagNAcVL2JjC0T2lK0OQlatUSQyX2naFbm4XQf
6Q8T9m9e8PoG0CJsfH/sDHsYmG1psdR9vXY8cyU9kiN/4JKhXD5At/BeILClQRsi77Araucle8bx
NMi/PZ8MYZmEvKt1+l5wCj8bA2oqmg73GeMhhMoNnOnWGWFWZztp60E0SAZDFR2DUX5hQo9jvWA+
vUIegesg9d6EzOxtOyGuzXQ10og8GinT3V9Ce9Osr0x2LbIPQKIt3L4Gq4fWliAPHNgYcLn+m87K
t4sgMJImqRM7j2t/IbFpJxIbqj9IpMuWyGKxXmJNfUNvhmCYn6BIdNdk+QEmKsVe2ZCg+Mw0XObf
ngpqq2G/+Rvn7JwofyK0D4YG8iukSdim9rsIfpl9jlp7B24nsfcadOIXCzzS3/z4OKMT0lHNcI7F
ol4RdeLnh3tpabGwj+5Zrc4113mXms78MRSTbec1tbC44nJXjkEX6Z9QSI2pso8pG/SNccTIt50h
4oxZQfI8KrxsnOlIl1rTEMb8duMJTaaKsWGGk/SPqLcW14gRXZ4E1sTp8pVo7CTfm6Le2AVBubkU
rlYDagAZ0szEXG/6Es+o1Sr8iMJDgkbro4tha41hCckt+9WlZw/8XBAQvI3tOdvWSdRi2doJBz7R
DyzaAZUc5OBecSjzWzqXrsCFeRuZGoTICBngSWrgc/auiU6P0qOj50OC/ZSXhwW1/kbnZvmAAQOS
z8A8Ey4gLj1gkJRqsoqvUerapHoDcLG4knhRG52LtnZrvUgI/fVrQS4qw9Nc26fJmHKZb/rdteUQ
4HnRS9b9JT8+iEpquMGHz7f6Z55PzC1O4crKnzm7+tri4d0YLtgEcZebCb9hlehotwmz2m860eoB
f7AFQlG+gBM8AFna1DbUoWP8sNbviee91VfRk/Z/1pCmfGAvDoFzm2uJIehIAQ9Ln+hCDIbCHrQv
glSjmKT10UKMX8LGkuW7odduhvxA5CPxqvTlEwI2KBKOz2Z6eXMmMlgfnOZOFHVwVCoEmjSeyxsI
ciHj/pUTACCeohc6U+j3J03iBFtPaLCygBgm86J4WUx+uAx3YFJYD8Gyd/cs3ZIXLWgQW88L/Xdv
w0a2XRTxQf5DfPwG43Dhp6PpMdFPBBQ43Vg4+bxCO+Ng3Ybn8Y/c9Zg/vVruN52S4/F/GX0KW6gj
eDv+CNt7gGw/TFJbIihIMywWPpJS0OzlY3zMN5SNLegkJ79TtGpeGUkvDDgvGF9bMbCiYFak7TQU
zf0BAaOqzxSOrc0SFuH3usDWLC8ZyFiPkbUSmTHPmtgD04Lr1z0l31hjxvehIOFhqpIM0Lz5hI6r
2/4RI/d//KzZTBwe+WMcktKCh79tHfOZN8nmowNdkhrelkCCwWwC8p/WICT1O0j+dJNg2fan4EN0
KmX3AbutxwC++9z5wrfOJp5YyJRMvvHi7fZk3TtuEW7S6YEVln8l3/gr7NZG2fo5AsXEsY7QdENC
iINyQNkHUiXUxoTyHg8aSHB8yzhdgRVIOmOZDoeXOiaENofpqc8gBQoPMYjWv9Vi+qA/LzZiQA0o
mmjvUwsqnJN6GFzEkqXIZAsG4UEQsyjowFfS/NKaGAcVepLHU9nc7auXFW2nXcv4YLSncIVTctR9
xLhl/iYCl6pFzoYOmntrGIRkIo4cGUXUXgmUDuo6edU1c7sQVJJ7e+QjStNzU5nP7QKcHQoDTcDO
zjbQVuiwhe9SqnLpKKsILVtnjQHAGLUcpWkEGgUKUtdmZ4iKGgzI85Q/TuiDZdScUy8CVyD6XM5/
bNSorP7rKajReeA9SKGJP8E16i6VcL+9Ep1Z9uhBBa6JFBVPoY15MCxQPjeQOsXSV7Lf/8y+6t/s
GaIw33qYJwpRG37tTd2+m//8u2veUZBQXNmwOzJkMWYrvzVZuucIHPB8JEv0X5jCsDcYsK2O9XJ3
+sGsqd4pDvFNgvdkcq0QoKG/PuQnyIaML09Cj21GTrreNmXgxiXRHPNMR9l6JxolJt2vald0UfTB
fBBGxVNjx8xVJlR+U9cPrCIRmsHHK5cFeWydoL0+WfSl0+ASWNzap2nvcya+n3c5b8OigKwoGwHP
xBpxLbUSvi3xX7uFhiSjmGOagjqE4LlysaHqHEHkSkkhkYtAzbHYWthPwFvsEqUO/SxOtVPHDpy2
UgltvK8pQfLzO4CETVPqwcSd67IZbQMd/TMAjw4LGmz6zJEaFlyEsN1pQcmP/HbwwOOUUklJ1SD8
dv4ySUzBekjSvLi9NMQ4TXjJ/nDIoSISmaO7qkcouAyiN8P+Mi6OK2wNuFMMVYkAKctFPQZWYHoH
++tndn5aHxVuuv0wQMleZHqrKqyijAjO/eFHG0ijl2aw+O1rMOBFXjunHLFSmycGwocapE0ydBl2
ugc5OJLtTOl2WTocR5xbhpojbpCYixFyFpZYRTjg8nxcpkc3e/FUWHB/Zaw8y7sfmdtzENvDzGXa
s8OJ1QwGBKxodScWEsKC5SRx1GecVAQQgNumC18L8+TiXMsvhb8dSJBIi77YHTmynzd++G6p9imD
McJbcEJbBNU2bJhG+fjvHrQ924+KvjvRCNEBQz6vK/tl3YjNMBX5Zf7PrRp0Wf+bbjeHsDCx4Nof
BYksAXHCLkuPD3cf3Wps8IzydErc6OhLqQgBEMZf63ZjOT+RthoZXQQmduU+9pSBzLPgetuc5dVy
tYuU8FxfRWTUvjjKlkWy56/HjNTO00fmjVPcxzQiAm87rFtLx2dk7afCw/lQfViEBrDZ6rBaB4JT
wuNoFjMxjjGkvIRIyLZRSdbx4wE3gZLLjk2Vwo08o85AIT7oYJlYn7c4YxwFayRd9TZIx48HwchI
aJipU8j7zi9VKT8m+GCxDIBroiY4dkuq0QATn48BtnYXreQK6VhCrwNUpudph6CvDfZP7nksrZBi
xDtkbnR56IfA+FPzi+L5yJE0S0rV+gdlb9UwIUCpV67vvu26kqo2yWrtDZcrKh6dC9/vpdF2imkL
5uZN+ubYTGd0zRjvCvxVpxWij48VWPRvxyZEwKiSPKEaPplmPy6K3hOXLgWZiUAFUZWKwd4mAUOE
Hy+UDMgZ448NGDx3VsUfysSymBX35VUhLtrvAyvUq8aKZRXwE9E+s0RPdLOSSUM+XdVBYb3Kctl+
8fybBFoQB4VbptO2hkTL4gRYtLgM6XJWdiRedyZUpmfcvJ82yoiUbrdED5s2Wz2ZdaDksJoU1SuL
8eElX42lM7AMmKcK/VBExyF9ZLw6AFT2hXA6Q5haDEZnOkiDjKOgIp0J1DaoETCzQA3zPr3KW5PJ
Q5roYpMx8gGke5z8EMHNIfdXkkaTUWPfQ+rDMr92t2e9ydMII9V4wC0T6yOqJedk2i3wKgYmxqkh
1RBSNuBhKAmAztEbZykYCJWB3BqZg1hdufs1Ouj3ds0fQpuS673IFdiV8s7O+4vwQfiRMNPG6T3P
Ukw0IAej3Z1oOn+S9z6mW2SkieIbicE18nXB5n2gJXY9bzdykEeZU+/zdpUeBHnCBLWxFQeQqzbo
5JUWFzORn/sDkkqrm9EUtJN5Zt3kGw2NV9siDK7MZ9tH9azIT4n6vSBXg2Dy6pNHgvZ7hlZMC0Bj
L54R9SC3JBUTDnc1sD9go0nXmNzqQL26vjiPgHnlIbnQ2ECGBmyhx8N6rUIuz+7vjUjNwAUUI/s/
AyqVsPL3Lljms2etvY52/DSNwaCk2i9iZwFuTamXgyPU5eEXb5O3+0Nneo1RYvv9PBjr/gDeAvN9
1Lz2buZ8lq4gVlbdiPD5tNXloWrZvBZYBvvAZ5BtVXdpxjRU3O+mqYHDUth8ZPxN8x4RG7/wLESl
ujrRRH8nrqKLIBYa0DJE6dewF8e0azuaXdG5C+Mj0XsUPOSwIjtcD/KPfpiCVcgY1TD9BtoVknA2
ZmJXE4r7CoQjOU3nAraWyocD21vGjmpJA4o6Acm5mAZv8EsUyzh8666YzXNH1AH8gyoHp76HQvom
JqbTKt5enYH31bnp2PC99IvZDHWyVh3b8loE70QR10dfl4c0Lui5KaYuwIn2sosimrlEV5F8mvKa
gkciJGCbrvDtXA7oB3W1AmWeYG2j8BATUdFkzklXkHJHuUwRVldkxExZT0As+FcqLZtil04G5OgQ
6qZxdwQd4pzTdEInvt2V2TeoIxhUUuPlW6gA6+O7uUZIoD8q/0ZOArNHWmjbQQr4h78WDsxt+Gq1
H7YUbBsUvBNaTZX8TezRyuV5WPI1kPukXmn3MBq4gZ7IPHGOe1hu9qbcJS/w6ZF2zP0Rcx+AHeqO
b1jDVLLK9MiHIaTPJVlIGROQ6sQLv5c2xTnkWJ0xwpzRO1ExSjsgWCZA7kFNxiCByRZpGYlujr8S
J6SQ3vt3I15Lx/Yq6fHpFiMTxMj3fVkG8es3doOSCAdeGKuJ5P+8Edpp8fn2yEScpy7/MvQVSotz
aihWDBPusKsvuBD1g6mXq+gAhzQLVqYN5chZN/KuIVUrj2Sh2XzlY8E3zJ20eBrIc5WFGAI4Q1QO
9BFoPq9US4cW90BY26Yu3RebQq+p8eKrg/odgCU2CsFrlJzcJPMkSOOlyp7+zVQbyfdRivBZdU6A
puvV9UgyhpH5qB2iAZFbVtJjppt+cA4C8tn2cwQJ3014SVfxvCQdBeNWjc5qWx26LfJPFMC3W6QB
cNsboVAcX8yhuh5kINNq7ZeUNgaxrGYP8h9OJRdN6dGVmFWJh09iDl8TnYULdyQMfSUbreUkWACY
G8eEbW5NTHWx+3GCUHIfkku+Oe0paoF151yoSCzqnIvB63SL7W87qKrr4J3BHjcanSp5O93WclP3
cyvRNlq8/P+XIkjJ/LbF/LkUFlLmgoEOyzuuMz8EG3HX1Q2CWJANeB4xgjT/2YxF4SxbpdavCWNp
UU7buqmX2AaDNLId/3w9hHlDHUA/PA96/eiA4VlG6yOTCrMzdd3nRx0g9P9wYbjsQVnym10/uCg4
L6iG3tpFyHmrjrOuwDUi0ye4tKjkjgxC2XwIxFYw1ECJveVQJDGDoRQw9zM6/HFtgzpKY+js3Y2D
Nm7/JeTuOQFg9h0RTH9xPJRmBONTw+3w7t6VfcSILUy0s0/m4NILFQEZvZMldp9W6xoWX1f90AhQ
aVxH1/eDwB3mp26P+xjdoU3NVH2YMc+N2DO1IE3VNAkAcMALXeBdagSp8GLoMyA+UDtOaeRAhFc6
fCecxXmeGpMz3OagbLEqLzVgOXApdGz7Wbg7iZT5P2jKyqbQTqhSM4wKy7iB6La9MsjiwbzrvzfY
zvLQ5o8decJ7m8k2xx01bACkyUYnAz0ZyTyiCXVpifVEZcGQhNZiv4x1Q9O/iIS23fnq/AMSzPIO
wLeYnkodyY+jFoT/xB2yV8b7F9xZd3MFiBk+eYcZJlpeHpC7W5ShQt5pDlU6vEiQYOespPX/hBfC
E3PvNY17pLF4rSa/aAfXzrk2wgfwxY5eOOjK5gWRRQtz37e4xGE31F5qL9JF5ThvP/QoXoJ4k/WT
TDzqazq+3UDfW9QZJzlVYE/g8ztQWuX/WqYTOWKOlg5VAHA+a4844LAwnla7zVI8GZonHcYy1sht
2cwgs7HnmyOX5bAdNUfkz/NdsaHRSUs5bNydt+EPIn4gJgffTeOabf0wQMnY+d3fpnSOumJD7mOg
YxVRC6/mDFieRu3/RBWvNpVqP+/emIDiLw3DzjiNyy0G6mIVfJrZJmbCWgsb2Bu7CRuBJ2pzTo4x
oelMsmmwExKVF+z0f/MA2vrfD66h0IBgRZdVFETOFAJ8+w5C4jsRxj2gcMf59Liicv9KEjPc5z7a
ayGY2G4IW7hYFCEHO+qFczKpT8f6KOlqc144Ytr0INLOF8+AJ4up3Didsh5F/q5n3ND+cPTJBXBU
U3dDthkTJD1nEQ25RPnYCkEI4cMTSr/GOknpEAupcKBAUjrGrB5lrhSdANZpM3JuTpmIuRqu1czf
UJYALEJTvmGx+VcxGk5FyPQuFGIQGK3COoo0/eS8VHJ0066cRHhmtaPEcHKIbqOpaa0VmIBKTpt5
QkJwOTq1D8Cid7g8Zw/s933byGhgwoMPFacILiKyOvPvkCavscsYfkmFW9zggtz29L7yUQDQbnKb
DophNrOKgLrZ79S9GkcEqnNmBoL/sN9YQiLucul9C1uoB+SMj8kG2WEeEa8U/JEi7tvk4V8a4uZ+
Mf7bagcBADIQG0UJa+eQD9HlQ4b6qdNVx3TNfCnlskfD1K93TdqE1wXNqIDKIVqQx7i+2cwMRz7d
qQxWRnjoZDc/cQeEmebjCBxw3H1/KHt2E187j2tD8wMKQHymW+69TjpFkTgcaLGaODcnoeSqq0m0
+uyABtGXLZljxvT1ZTMEpJ2m+kNQhduADOSGRAUDK/cRKcKQLFwF/gRyfebMXlV3mgQl1EPQvhcH
VguG5J5h8E0Z/iFag1HZjsMsNInRYMd/7ZjrM26cnAG2WpgTWGKmEsMM/dTHvdGiG68Cap6SYk+C
FcUHfMZpHSXYtR2G5uLVglYeRlfUu7mmQsqYL0NjRTVXL6aRUtV48UqrMXmkm//cuaZGjELv/urb
ZlWVQ1rTjttJxH5rnp82CqRh5H80T0+36sKbu44ijWXmAFoxum75GP1vnhDy/8T+5YvYa+2MuS3C
iXe+aE7xSTgtzz+aA5Pj/e6AQrXlptQb8lswga6ThBFohyzVqVnBAxSu2blapnYJSHlso7DGs7Qp
/+6vFi7CN1ivdC8H2gn0Atj4GtCvjdzxCBfrCiJx1mjIfUXcSmUjMRPqY9plrfi1kTI1xOZd64iD
9c8vOC9GbT6fERf7jvd04SzNOzvo7mFVwHe59NQzdteez2bardeaUMyfR32fcLvLuHKLCByx18g8
aM1+Azxc1N0qSJinmFrqNMj3yOmn/H25NK2mCApyN+pR5sE4iJEWngK9uwDgbmssIQTq6oTE6pgn
/jn/6XOO6+epVJrsj/oSMeGvntX21nnwmQQSYJMSGU4IFNsahDOYGywpUYZHcCvw9YFmkO9ZtVRV
t1xk0GSpCN2nsxTdzgUznZXzvCXux3fOMnFtSNALAmmQx6LuPKRsohfIT+2EYfMKXsqfhuCNPnOf
cfMg4yfp7KxVZGHtuI6wa3yh6nD73UjzkkjtRj5qdXrkO07tQZVQUmervwWKTbfYnI1GfgIVyL68
0OFQ7EbXiA8lA3ziiEJV4OCUEsly9aHk0LjIsSXMMj7pf7RvsSEvS+igNxmVF013mDflWs9Ywhc2
AO2FPVa/bfpFdwCiSPRcu1YpGc2kG28p0KoLQkBNA+JfNPl2j2IMEZ5wqZgkB/anMGbrVAGT/PRb
BVWOnbJy7B7Q6DaXs/qGVolu5HUNthm7G8G/VlOyFPIBQs08JojEvUlBUhzdl6rY9TLDqwtirB0v
8OckNbXIU0G/h8K6HMRVn4a5+ier1D6igmKCtBKzvxKdTH/7hE4Eu5qIQieZCS89qiaTG59lHCuE
kvKcPnh92OCFkiO3ieP6ELbVvY80JWE3yewh7rxVErPwmKxICyHScSWRv3ivj00sP84o8jmGaDeD
Nr18EzbqKpFlvH4paoj2uqNNJsLd7yAjSiE+/+a2wjjOlUXJnaNePaFCwv/Yc4v8MyGVJRyHoQ5a
UE/+BjbUv1Q63M0sysUrTogO0NvJbx3GE8zdFVPz0TPGb3oghEV0lSuUx3x7KUlsYYn+lOw0DZfQ
Jy4uwGJFA7vUEbiVwb82UYVQh+uPtyC1RVgrS2/URaZC35s4+4xS8FGZ6CTcgnL4uC1fR69ymvQX
VtUCrmjL6zVftIjhl8XHzVlEpn1Tfd/UuKortplLFc6qVxMn4Q3kMvu7ofzV3nf/sFUKNSHmnahl
15ahNLmjPTl3Vvn7t1+0xmhVdGf4KRauQ5LyyTbg4ShFoVfIt+MWGb7LLMlbvXpx4JFe6kS1TiCE
u/S3ei6v+43h/HSzUmHoDsoF3yQXNRjLqyRTxNOUuTMwwrO+vFuhyijjKyhED7wYS1+U55wCpYsN
E8YXnV+y/72E6E1kvhAAIMsg/jy0LQ35D56XZ2nUajTjvjBGygnEaQVa+V8CR2xgI7Tq0qFKlYCh
EkSbSprpkM8E44LbP4Ig3siGJu/UH0sdJDEWTe/lFJguHak0ELdBdDYbohkpvSBD/GBokZgbMHp9
qYa0tpeDBX5nkBDejOqK0alfW8SBdqxtDGEfVEa0hzFEZQWBOx2v8Q/IzhOyx85TXdvnMevgwKgP
a5vlOexhAchKYbxbXi+Yxa76TH3NZWiPnUQ6d2zZZMSoM7vpQDJI4pV4/GnT0+wP4nrilNpBw1Ke
AZxp9vn8U43YbyMy+IHfs+SkjMqy8ynKsW9NI8usyxbAerLe/tgtD/rm/mXJEQgEx9CvuZJkZa1P
//Wjh1HbVzPK9sY9f+Ohw08gcGP/4Pb5Azm2K4tB9Igyh2ZsiNkwksK7Zrb+bETbfJ/ksNBDMlk1
GZ20GTK/ABIUjyqG19Hs9X0NXQqwfT+0FAVWsAxuLjkNhiUO57CDwBHi+J8Y0D6B8ab884tkMDIL
w5jZ05+IyiZBTLQSQ2IgIaNJIcAqTu1LhPNR8+2g7VE/O900SEBlojr3Yeqd2+ewGNuM/xwYsIvD
WXcHaMsk/SFrrAW75iUPykXr24NGMw2Vqi5vknMfdXu8O+hT4VAyV5Z7FG38Ttoi9qwRD8xp4ma1
If5DCZVYSRUeHKky9NYCUpObODryzTD7dqFp3D2aMvEplGmlvKp2NuqjUZk6xyLGtH9B8chX/CV4
wn9JSjQISeQ5tpT925bbv7FP2XEBGLSCmvfDNQdcrpieBxqIuQGdFc6iMIWWpgRW+O/e0hbmY1pC
BkQyPtrHJtlOmKHHPSjqZ9jOKaQyKBgKooRY+OagNezYE0Tu1Yb1XCURoJdpukX+W854WYWx3moN
SmE4LEXeX79cG+AxnEDiAL++FMoqxgZQDvDW0GV35aBzgOoyPhpL2dto++G1LNGqBRprSbWMnZV6
Ud+CfwNcafZa+Q92oXnYSg0g9+akV9rZPdrdyuVOxcIfTgbVpTy896Jok5518B6I608FsQy1tUur
/0JUccwQGRkfSBtNwq4UtpnEhUQjBMPZGqSGNy0dyKHPMt0/sB/2s41tfJmfRvbjrFZjA6+JzamJ
UFdUK1YEiA1VVmyM245TUXHx2dZMXg6HdRhUW4SjvwrkWUPOwjONMF/lrNSdv/LVnEpwxbT4mUnf
jp7uqLduYAZDNbf9SpC9MvgFkMFbmTZZRjRYlxus1EDJ9AvCr/eC7NWVjmUhhC8QPDftVLKQQsrb
HNe9Q5lQcsjOdeFT+qphRduD9tmb73ZH0/1cmP654WnNKHTPTcpb8M5ZhLw4DDvhkyiKDd99gzD6
sGWOXx5UUpt0a8XOrYOUmyejVM+vv4BRvzZNBEhu9CekB88MoPL1gYP6/+CC0TrMu6UkIXYMUUyf
8fYnxwC7OFcvjbhAtsDJkytahqy6Fj4ydJI5wIgd/MdKWs+XdTMKLouCmLcs5peSOlRKXjw/yfzs
r7PjtduNnlYAgonwXzj2eauBAHKBb4atIxczwoj8fgqd7uils8wFJy6pp8+KH0F1cFCVGDsVNBrf
dCralrd3EDr5t1rfcAPowZEX0iEukDvRST9v4N+SrcOplaX7KWkX9ltlVBmtnSsa28YNUtxD6RYL
8ZOoWUEppdaxdoe77HJsVUBMOEF4cbRBwhjuvuuStZeBL8lgq4SIGTflMmYWuF8WvAwcABz5LIYM
JFfcycyZDqbEon7XNIA+DKd2Ruk5ohTafELAv+HQ8u1LqgJGE6pfiygMhuGliGM08BX5RQlRX1tn
wFXD14dQbVKt/ksc+SMA1s1Lses2ixDyRvFGFpAHK5PJPncvDiuEwOdlHynOkqzO05JNUfzBFZdX
XA9Nz6bUc9rFMfv5j5ZIBcAaiNUVy8an7xyTQqmH6f2uXyizihZBhZ/UVsV1idZ1hxjil8f6Mbwo
vah/to18QzEkOaLnZ34YH0FJ44cLanRhU9m5EGyTAApY48b1R33YbnCT0sIso2bnji2/rITbOmkS
WM+J/c6XAxsHAbbOqiheCkp0ks+owGIk/+bdr+FbgtpDoGFU3q5MQSOPoZnnEWv0ExJGi18h7mzu
ZdbsHQzZIJLRqDPB6yag/FNgY3N81ddPRB01cELS9L9S9XIo6Sb+CdPz4c+TjzVnCBs9SxRddcOF
7m7f1MAqfauDeULZS47QHAUz685t05aGHwE+G0TzoMsB3FA9EBoyNdXhRcGfbwM8F6woEj2vgWGQ
rbRQFLg9MWD4tdxiVfCgkb6xQyUEjz1lwHowpkrn/AuSOySF/ZWqNFHweKKAg1WbjLrNMn1zXaQg
w/YhByQAOAChR2N1tAkPr3V2FN4MknsC1yI48+TfqNt6DLDEl5vnesrY4fBJnipo8eKGXXB9bt7w
Tp4VP5GrEXekPYHt0W8PkhmIrUApgNERAyzLJ2260GBd9f7jnejyryIAvkKNZLbcglCuE0xueV1y
3E1KtxDgrQj/g9FHVORzDpwfVDIhQlQccn4eVm0LYsn1+d8XaIKAo4Yb4AnWnsU0h0SleSyaf4r7
ICFZRmnMm56QmfXKII7KPEutj4Mr8x1Um17w8nzAt2cGkI7OYVm90OUSFIAl9Y5ttaAJWFosWjrt
JcY4fLul2oG1j4ycLfyp8fWhAcyXCXOX2oiAysA1YckXL5FTFBHL1m6GBgF/1U/IPlo+wK0wHEWO
r8Rbd8UwETtp9mGKBjX1LlaN8h0j9tHozYIshIcms012VHe2y/fFb5vFhe12E88zTTeoKEX2lyAR
njX4FTo8cX8A5wUt4tDkd7qOD1mhKix4oHthsq6gytfi5A0Zj81Z22waBHF2rAIwMe79IUOQkhNq
eiQaoOEtEY3OPaVUnwoX6BAtZ4fr503kDgHJsP7I+J3SW4wUy5edLc8t5Zi8OnHNRTUBJeDt/cUf
dvzS2WN0C2ygVW9FxpNHA0tU9hX9q9os6vKis4H2JmDzgCnmWdGRYSBy3+ZSt4/dsSdmopLdDuW9
MbfA4s25W7l6usEaA7RXivYbv/YnfO0oIHkm0kvWC0VZoIihkxwSzZTk5YZrcB5QQw4bxcpj+eCO
H8z3jQv4QYO1gweNAr4XzYrIsWmyTxchdURdxPdPr6RLBxdQERJKe8os7hyMCPLlxvXN7FfRoIEh
vSYip3UJuFZ/niLWw/m2Vq2s7vvjqRs98rGUprYZkl9D6MJyzKTzCy+TX5ogZyqCpg+dRxDwbOSz
uVaOnCWQBYGpm7+0hLkSNhzBgyOu1gBV+pxXtphyY4wSAI38ToKpqWQohU6CaCwYIqygf/oYVctX
2jhJVL3VmXZC6BieASN9GgQu/NBJlm6764H1QK5nj9pGStXeugOBcFeCkVEO5DkZYDxpp9LLoDw2
Uzl65SVd97srD+uuYy65lLKfCufbkmLW4m6j+7bdeDTnluQEaT0sxovQ3GZ7T9t7N7hsDNxV+Sqa
iFN1BCEMMWGLYIWti/ZJH5yGB2jhgWC2vU9JJ72CUnklzNWo6UECFwhu0ktBqSjMJAX7QMMGisfB
df+8LSLQpAxgrt0tINjEgbt3XWDjIG3yzg19YCxKS6xt986eerXa+9tY4ECNDZkS7H7+PEN8ewet
JvMt/4G+8refla3vgT/iYTPeKscxmypnXBUTM4MMfboNsSnkLsiPRmPCir/Dvvq8lMhGk6Xw0Ldy
/HKrpGBwmc/MLzhW7pvsCKnMMWRiRRhyqZmsAyXMaAq5meXUKK4cmtFeq3CIy6ig7e/YSnlFr6UY
+XxJuAvcjT+lDnVwU+g2MiK/9oa5zqQG84MA+r/UKzuvjvg6r6GajImQnMXashJazQDYFFVrhZdl
gclj0EXOvaXZ8TPbZS9jOQxLnz5LPIf3oEu2y/FLzNtLATwKvm8GlxYBLTYz9R0juRnshPmrGvl8
iWhgY5I+G1EEas8Dcv3yHqIobtibbvo3LJTzABF8RyTBrSMOiyBAZ1q5n/jKpRVw/7eYSKW8ic0Q
eHacoiTDult3OWuxWE9GbqLZ3iWM1pccBtvPKb016Cxegcol55bCOhFxGtZg2FOORJ2dneJ4loiq
WyDoHhh6wuP23FsqU76jUbh09w+xJt0gjYCRRdsOqaU+3tACoF4qjcYE/32N8ffPd2SlisP2lFDk
KAD3HymrsJ3ANXETwAua5zaHQVdeKfr02Hz1PJoK4Bf+UN1wUeROgAMLDsI3A8p+2MHyarpPoaZy
b+O3qmnAIiUibqLAPNWEBRaKA3Cm51vzK23Z5fMXqvddokPK/KcjOe4vWrFXTjQY7LvUn9axrKQR
DDqd6mcu2ka0FBAfG+6WwkaEiad6QCD//n5bZ3DGTTPpPlAXWe65qcEe6nKhz9GnJPymQo8jKBsM
42Gm64ZOZN0WawvIuGAqXUmEIl36pBponfstEGcnDRaY4Qxkb2SJtlJhQ5l2PPT4Z5n6/VqoHoCx
iSiucACovtwkbmcoGgI9egqBBfAn51Dr2yGeNIWxJoFbjxYTMVSjfRbT2Jigm+68gU/WKTKJTIFO
0s4dRAajLdOAAIU1g9keVto+W8SjFo+yI6EcE6RTonT7Q1qqPOBiw5tsm6vCCP3R/ZDIft9vmbmF
iquCQ5SGieT+QHFmq8aUPKcCZIghIlK9vqaGwrnkQ9q2GMPRWuRK1X7kCVhBNWpdhEIdgycLAYdk
r2FPpQbyc/WLXd9MRFngvYLpzCNtZDlRNx+ANkpcLALBvmtFtIMWnjR+xXY8IexGTkQtaxre+m4L
pby2Xapfji4UAqbDWtuoxXPePsxlv5igixyZywFeaFhXiqTeM9Pb6S/Po92TtQHJub0BSPF8PN7O
yJ4daWVHevyBbOgEBtkuskNZ/sRd9U6+EF+W/zdP1b9m5oc2pshiNwrlQwE+ICxDBN/IBsP1eJrm
p2L5+yOfdF2UhSg1qcjN3h2vbI1iJB/jPIDfd8MLc2h1noQaQ6Hqcnpt2p3eZ0AoYMhgA1a4C8nx
Ie5HQpNBWbHhG65j6zz4UOb6YlMk5aT7tMWw2ZG3kkJKrfeMFZjdG3NsYd1pKhVfrbajn0EB6e+2
sa3dUQT0506A4STWHV/MxPBpadENQxHOg7qo8SMX3l+CvKwu9KKBh1JYM8VI7/KBCV06Gtwj7WHj
X9ZtOFhmFWD/z4T+xZck3k3M5P7XcqXVowaqUtgQngFDn/u4yB9lurbUSzYDelBMiwsdkUZ4FX+0
/x/u+pzs6//fCAc8h8Ul05obYecN4+/k85DPWGBILjit5u0CNAiMaZQJ12bGvZnHzoK3wHaOL8i9
wx+30+IcIT/ELPRZSBMotmo2RHgDcGoCSZed8ZTEMtoSt9ukeH9Klv9BJ6nW2aaFqdLFMhqMvhBp
jIgfeAu9/ePH8AEaVdk6yksZiPB0JvphM4T8GMft/TMIxHJnculnaZg7XMFfMn+tRkU+Hhmd56Vm
GKAF334ig1ymZLZHVpL76gFUs+cAXbUAxFBMVB8H/KyEkT3v/DYz0TTzCqc4lpH5xjuK4KUaoXQV
Uv5kZy9Pl3FMJzhgKJO2hR8+PqDVZ6pRusDrOxa4pN6VgrDiFgsDelkIwrk1brWQnBfEiN/h3IfF
0pkasoYf1HoKri0IcrNpHegKeBxl/77CCYyaK3GS1bd3z0AqPGVlm0fYbeKsw/hhmsWFHlQ4UXoZ
v7Ky9CGjr2jdqB/x+MtBNYB1f/eM+wCrOpJMDHUKL52UFE8fTGlFkNI6yLhbyZZ0RCn3JOWG0GhP
5penGOZkTnT9p+tL+qb1K/pJSRqnYESEITnKNyLsFpfd3WTCymqBrdhT+zbBSMJUV1pBgWM0bYVu
0xlDeLywVj4oDqNepPQRUGqGFQxoLoWLp80oFks4jrpxQ0nAbrdnbuyh/xmZmGqWr1Zo9XQkA1Vm
YP1RdUPgG7VKEenglkVOBbUWh3SHGeTee+KxjYFaSvrsTHR6HGUjYZJB211UbOapUDAJrYSU9XN/
Jt0nNcVtD1MKa6lPxUGM64lT7h6QG2UIWdP0pVwqcs/i/v5B/GU2yWpTfU02RmN/nvDzRYFQg8fw
ivCCWWciKE6SVb1xn/qXuztTGC3HE+ZSLUF0ODX8Zo2vl6WY4+oLf8ZziIW2L50PtWkynAJWDwDD
3I4cd6Xun4T2nStrCCVdGRulEWf8K8e7brD77DEgw6o64xOAmjRUsyI85ORCAW2O2hAF3OjG5sYa
WyQkDFjw/zYBkdSNRXpwFr7JbV+/XrlC6DS1Mu9OKUb7cXwfU6Rmh6V0FdlZ6ZIHK/eO41w/RJbg
CUQsbvDifYNZNMpkANSt2Sck60tg4+Za40Ptcw89IVcNdnUkaTUa7MN3nJnrceVOFQrPlxX9LEID
tbPdoY1zt2eBDU9h30eigsqGTlSDEc8jG/YQd8yNzgrmz3SbCrCv4WD9Xk3ymXmQkQy03oOlYH25
rUMTMStDNavliLEKRMBivWdcZMz4jX4TG4Ov/7rZ8woIPGmubEX65TpNrQ4UDg4MzpVSeYeIAq+6
t09rZTx6QNLDt/L3eA2Z4pp6zAe+40HBUxaoavO3scr5PbWEmKBqfWImtlZY67u0wSc7gBNzTU1j
zwvosLHCOSG0WH08IlLbshtQ4M2YSZOYjCqMuR74+DsrcbPCQyiS0M4SugVopKjfQuMI39Hjgxgo
fyfPATots97OdixmZehOTaANGWqa+uiOliM0t8NpZL3Sq2Z8G8/LN2BnK5PefZmfY1Oqh4acrTyM
TmlGu4gnNkBwFX+NNEXbXovP7JI2Skfs8QZS6lZY3Mk/x1vLs13bY03VUw7R+X4UB+AwfsdzGE5T
PxL3h9hF+PoXpjESKKiFZ8X77qOm/y+7b9k6xIgledtwQ6OqM6001lqpGDfTwJNLrdiGR7hxgToj
5gZnhl90dtfIpbZAv10HO0+9JOg+JTX9L+C7silrCSK26zqiDCIPeJvvtm2ItbJpJeL3jE5eByU1
WJOiQZqTNPXSx863X0Uy2AxbY2z2iXVs/5WEEL0vMm4Dei+j1o5mb8B/tQVnwMvCKxCoYnZijtDw
d0S/XtfDQDphnUum8cejXR5Gtybe+8zvHiyVrquSdkfL2+IWxkqbn8UKy6/onN5pkEmFhRAXrZpD
aRvAoEK9GYDv4B2O7c8FlgAaigwOSF9ywLG0SPFDOG8IKWHIooY7PKnHxWgWINXozKkgRjgjZq5t
XHZ8MNbnB9YsNIhVSyrP4Wd2Xje4Ixzv5m2xBf6fLUSLxNXibvaa+LjipJ8TkNMSGdLJJtb2cBpQ
VQzfxAqeeF73uzaUqZ+SeIiq3vKHyTH8orWQVhIjbSzTK+1GURz+DIkvzhUIwb2RXRGPppWFgXJV
P3pTfdFMbB8x1PCub2yozZtg1IFtXnGFzlBMiou5f4G+pvrT4JwGMuhjAUgxEGw+glQatsR6qGwp
C/2eSue5nxnUx1wKKUz62qq4GQl4RQUDA3QNvOO6BhPMTHUPmYpCMxDoan0wESweyvv038nrUCUb
XofFkJKuwhZRLuU6R4xIawV3/ccgGybRxXC6rRgAs/6RlkO7a8gICwwV9sdQ19DRoUlw9z3gQXdf
vBAoCFM+p268NOe1uNKlyCd5zlFScV5Y3/2dNwLgxl0xZ2pMLhJZNszOWvMYHjn45QrmCWPfIJuN
qFWkY5lcVtM2ycLruM3Gz9i2PixbWYMQtY0bEDEJt+WiEe56TkqqPCq6/ZqA/2YwgWOgBrZGdCnO
ueUupPTSLIt6bxoqwId2916ByaKl4iqKf9RFbsNIIamPzIxysTuLW44iZW+LOW+sYUZdN124Npqf
HYILAaJ7AksuV0IFrQSKm11PDZHhh/+tK+8aIpghDYnMqDVLA7Y8EHefusCrRj7CMFAeHuaYQees
RphztyLwWn4GW4930cif/e+X+z1duwJNzOaLkkHNbboYxWTWf9qxXKefaO1A+DWLQ4foR05clPDf
RARNZvBiK67Nf+5aBiXo+4940jslIBSZboJAO8NNCXnpU6MhMnK8mMM7qOrjFG4qWoJKtlTH5IK3
T+YxIexokJOjIpmkw58pp2KR1ywPBSnw2FRqAaYvEdKPJfzTE/Q+EX3Xc0ic7Lp39BMeh3Jk7WbO
O31xQU4MYTaTcra6Apitgqc13g3OfxftYz9q5xe4Q8jDVZEOqpCDM+mPcFIaFsSKA0AADq/YtePK
uBsAnzmp+pH57Ss049Tm9DNxkreaUxfb0CPBzjqUkeDUwcwotYqs0ePneV0HdlznR1pq+ejd06pE
a0Tu2U8r95jhFEmJbPzBAiTPylkTvvF2egHx+2CgorQx/7jbeUcKrBhYcFfB+ctpuWEeRSA5ggFF
D3DK98dv9xaCblGx91U900nk/qbPTyQ/L56bebzBBEYw+R+qU59LyJKLSwd29/eKwQii6RWqCBvP
log1iS2sJ9Nb+yiZfxGKeAIIiu7S0IT2ejC6bCw/RRYPRofOtkp0vsvg2jCHvFI9Tgo7esEKtLdn
DLe4NF226FQz17+sxDUoT9zUu3s/Kwn/V5NLo1KKSnf9OXPxlZLb3GwcMHaawnNw09P4faKG8+EH
k5/G5XEZ85ZXomtHw3Rzp4MB4FtrVPQGxXWtPunxB74WOi98TqxMLVQPBqYCFkMPqNbXmQ7jP66v
n+tIYxA74p2aXNAkRbwe0pGO5Cb0umCmcOwxCTmZvHRwzWclhiXJX8oC9kgoK6bElq2iZGBCA6sU
M/LdJYptMEq/kjx/nGo0/0GzjJs7F2y6v21vnQlyN6NMWIxGYcFRWHKIZdi3aXH2yiyRWVlJemQh
8ohgKVxS/pOQsDCPwCuPzSnB1WTqmjsJtB/smAnd/GQYBRwk3qDdQJsBEIZbWggc349iojp0gyC0
S014B7s4GdUceGtvD8UJCqnVvyJM0RNGwzNPfa9D1ifi/I9iEobpMAeybNO8epPU6xrny4kQWURe
SQ0ZbJHg3owsblp7JV3Psk7dsDGe0VdFdh/2T3P7zp3zMC/qCYr+9AVRy/lmkUKs6M1wbEnq9BC/
97vnVhMtjtoCG7wkm4Tp4L6Wmf7WABthygk7XlO+xXL0bnoe3ERd1wiiVmJK/I/KVChkQVCvori+
VQWcpGzmHVJ3v8t/7XgwUZpO5ta7Jl0tAkGIYObpS5draYxQCBAl2K6V+aAIDn+sqixdKNc3Gy1V
DxmCEc8VCQpoP2YsExPpQP9F3H7wPouRlt0vpvUnNZ/mE0Ol8/nueUKmcsoPwzHIMX/okG93U//d
tM5IWDXFFxOgVmuaoTFXTcoZhuMXXuAIT9tt6UTu2NpzzuXpYIqpU6hGyMYjMGP6kyZOKdyDJAhP
WtPzgJ8Q3nHD//3AUov+RAMgm6o3XWvtMTi0eqYXXQ+Wp6aLR+XcYE2nWnapF0JvWupgeD3cA05u
qd92j+6JF6JiufVLCChcAzC3U8uqDiu/clyWS6aQCm86aUCJ2vLeb+k169lqOPgPXeRNhtCnwdRt
yI+jxesuNgYXSeT/hiiGKdJ7uDyqZJK0FwczXl2lBCn44bBnbB1hNNxqVPaEtiT/qnDyT2kT4HxX
CBWG2b79iJW40ufLXItMrSwmhAWoRSZVci7lGZAI0Nl/bxfZq3hyBE7aorvp2tQTLQqgKWJheB8Z
N5pX8gDoFLNiSYgE4J8fz91sT50Seoz7wvfdh4rhPHqVwHQECDJXwsxNbAoHujmmxjM8EzNNUbmX
wCQrk6a0NIYTED5ohXkPH2FT9qRasuPid/NaOe90uufeGesuyEgDlze+eF/Y92shSw+HhWYrVAoz
LTA8IyIgpyXbirQOgkgmXh2DQyuGEzfw2b3qrdXuDjDHAdKg/FRk8tGK3a0NgTG/3+qYQZQpVX9W
eLUdTGJluaEvxVdDLryhwtmAKm3y5Hc8AXQjMuyBwSJVWRXN+nJw9shN/QfUutCQ7VxwEBZhwcvH
KAOF+EmINqvRB4Zhs8qdRe9kZ0Cf9VXZvOHqTpo0klxYERELxKH42JBrvzDEgebCZeA2wEAFUDxK
Us1FI9xLtHq8V9MNJzS4Kus0IffKfAhgb93/omwqcv/r7CTW8DjpaOgE0JHF20M9SJYxKIsl/laa
mdyywL7K+z1yRHYV43Io3UM4lmvAM7lkBnyZSqzCdkYQbqteIOMPS+dIqodxGb9cn9mdZREEgYhe
QsHtb/ymR5CyAyLIwg+oYK8nMn8F8iqG3C88HF19GLKvTH0IgeXFn6u4Ii+iKO6R3lDzOHREtsJ/
CufKnlrz53ZPq06Iwh4DzJOCFHFlvRNdWeV/SWUR+HO8qVum8z7U0tkgec0ybX4+QzpAMbGfqObC
CCQUu4J+0frEwBrgWknG0FbnULVGtHZpb8g2Z2/6QBsB+5m5Di/2bEpVW+w++eh2RBJaCcYt+Caa
6n7wT/qzUGpk4K3yJn3GJJPO/Fr8igkXrufdU67l73/sK/Hn48x03Q5L7GvKaaKkUyMgZ5cUYwR8
pqkqyi+vWlXJcyJhbA2+WbTxVph7G9w460LvYqgh5g3iG9OpSSZKTtVJ17X0Y5+uE/PZ57DU3m3E
GTrTg3hTakY44TQc2MwqhUaon/B2QJLEKGQlbm0MmLbq8vQ4Q9BX92OlA3KOew1ABe//HWcXeBZc
C7O5YUR5UTsgBrTxcGw+MmHDZq6x97LO3fftBOYHdRE3MucoYMiF46HOXp3WDuJaZ3jnPpClmXmp
vV7R7YdD+r92gFzF9w92gAok1mgSyouH4j2RnU4SEy5ZihzLW0GLQk8zrqSiE+7EgZM93ZNGfW2y
7+lffmIe5FUKDg0ydN5c7itfI3vXry9l1A4/BO+w9oDTPfsBzTDRyIj88Ig2g6h9y4WMVnFVZ7gJ
eMw+Ju6QG07+6WGOQTbRhttbIAAZis+RziW6/KgBWFZdPlpIYQOiSCwTGjVaG1cSS9lQhWb5z6C2
Be6H5edXnx6PK32Z3RkqDiyEqCbkcY16y+CvGXT80ItOe2jbZHmMTeKHoaB+uSJOAVY69QHaPlL4
1fUXp4tMMsNtKLjjG8E3kl5piMGGwRE5GgRjky6eNZ6vgX3/kuqIXOpgvTr24KYFqUZAPwMsz/j/
kGhY7X2DsTv04pLZH6JeatmoNHbdnWwWqG9XsyletOMjt7kif/rBe4sUIPi1+QmJ8Qp7GUhjlmRP
bXXA1R6qnD886o2ECmZkbPI6YWQJC64mXp2zf0nG+2a5/yQ8ckU8spIXch9h9R5hKg6oxMg1cn15
OgwCjMn3I88zXxnxsdS3/kZtoo3owRGyz2GkurCfx/1E0majIZV6pRHkkfYwM3iCF41LOAH5s1gy
Ugp+O5nkRj4XpzJEpoqVatMO8+hwGvkT8CaWj5PTtQt29TYEIaiVgf5mBVkDxriyzIT+pJZdd+DQ
4nNMmrnGGLRLuS8zOololLbqvxDJlAoImOs0ccKO0A3Dl9DbqI36yFntOP0md29RUTvk9kuqGbx2
pFM+7fcSiVz4AmqWrwbFkJDAhKv1nCph+aeS30jjWnZDP+9Ix8a3yyEvRfxCTKQxKELTPlKImpo3
zK1kV5++6hYq2/K2PcFUxPHPKUyxUCgPZGJmKVLUZi0co7ffKH3dMG4wmgu8xDrBMlPqfUqFrm2J
3hBNQnKhaWY2U2n2WHZ3jzS/Kp+pwd/aEGuYQ4ad/TYo8W3awsgkpHYvBmA11hO5KjWekXRlUp4l
QTsDDLzUub8a/hRT55HBSkef68E8VRF6bqdKJ9+6GY61TjL8222VCa7xS9C2XhG7chAkQVGBSaT8
AtgJL+Iqk4Az1fvBy2LTtQl1oQ/BhNMmS54aenunbWEMzDCsPF0zIi9vveV3RXsOPYPOKafLl4eG
lS7weoyNR/ndCwhpsW0UxZfw/GeQYo9bM9Ls1DRuW6k/Thc+Yg/LKlKOYWZV11Y3wQFI9tZ/wcJy
kzWPNSG6y4H0QTfELzaDd8AGtObdMTJt27g863cOvQ9orp88jrGrYfnSShxYceR7BnKuaTpRMmKZ
OLiW4u0BOTrYM76hZwJgChDBF0UDxJColyIfdl9UQT8BCunRkJqc3KoLkQRuRAUWOrXofT4pYnST
kVjk6ykxQQ3y7NjN2TK5wSkg2Tt5muQS0EoSkR1KH7CKf5qiWdjXVyByyY/ap8pqgoQJ3CyijEgo
XrhS2EwComLEQuj62u8zdQ40FlTOlYRCMccSKlXBugLLEuPk4Kt63NvoesKiBPwqRj/vDYte1qiU
q7djXWj3UItSGrvWF0Jod6Id5Jup7ZEAvxyEMrs816rR8qF/m0Ez7/iMwHXtYOCC6vRPwAX/T2u1
FfHS9QjXyr/B2Sk0L7drAqTSUfEzF+kQzk26h5Llc7qaj0mqIZpL0XmajByHNP1a+anY3bp+WngT
AGEFj4nZCi4+H21n/RTuQwbVH2x7QDmhuB8s5L+Q/p1OwbgMyZXtyhg/gpdjHT5iB/c8ZV9sbi4r
tR8n2e3svkrQwPXe5khtZNUHJRd3BBgioECVKGmlY/Fcs1AzYuKpCnIlfHY8cUNYqMtr3B10PZD2
O0b3gVFqp2SlEuqxa58nZRLBm7Kl64oBB/sb811Nx3FOg/d5xGJhxNwy8S1IXiuCFhBK7DY80+XA
qk3dvDCEhHZfVH+ZYninvjfrz+zoUWAXm834xP4TEbS/iJEuoYmqFzKYhZQ1qZ+tccWTew8LlUqA
jXRqRv8ODrei+gtlyRo2IgS4Wx3f6+SKqWR23TKNBMGOTvXpeeE+iATBTfg6Ab+Unwy19Lwq5LuT
gPZZm7kym4TmNMNZ0aHFFmxqQU6wbl9HDsMwocO1HHXqjhKem8aZ1+HSVMFBv2plMn2P/i+m//fi
CRtD69p5OvPBZwLSqrod7ueo+7380uLd2qXyeMvGGr09DEa2RG34Ld9NvLayYHAIx9jL5S83n4GC
P4BAnGbV0WKAT6jDKOauUyaY02yolO/ud+buqUnQyjFNdSX1O53yw0Fto2r0dYpySQ8MfbcfilaD
dNhOXa+QQ/Ew4qQKIblPidUs36zjc1y0pWeWRzPDD52nI0Fg2SkyPnYRm7OcGUwZHAO48yUn2c79
O75qm+qHaQCK7Eq1xlCbEqJj9059TpfntgMFd/dpc174XNXJ41jXcI4wTLVD95zzrh+jgBGI1AcG
z/3u9CBGXv3cG/FlpyAYmbzIvZboTNCp4Kcn6iKfjpoJ6DtWVc8Di+p6zqeje/2q+Y0wd+BwOfpX
QH6O61TI7LjzToOdwfFo6mY4xgDt4h9m5ub4IKf8Mpw1mVgapZ5/DWWMyQZEGc2C8rykVTPZNh/U
VwFi90Q/okMHbpDqNPvzA9PuqHTLXwAkAzyeQG2mH/yBYu9hKU8bTRP9loDINzl4uUM3BBMaxcrG
Mbdtw3eawoDwmqVM7MWTjd7cirTZceC9C+h06lnzy9SUrA3b5zUUHNU3cAbtST98ry1EJxxqhw5/
iKc60VDQeKJRp/Y5ybFGBEIBJJn8KePRzdQB0pGvMcXHkPlW8JxwArfiVgi5CQ4B5yvhPCpDaqv0
kZl8mtX7oxixWcqrbrLg2RMS4k3H45ZBbaIuSlzoOaqa9NsJ+ZDHomn64a9fOvNdH+qzVu6gSwYJ
BIJgTkA7udsltagvEOAKzDF+K/peI7N7AarhstQISUm/XwqNraMGUxFeIKTLUUoq/CDjdyLXv/6E
lLoBBEYGTAWFQ1SSPMqkbkf51uWOFh01EBZAIKyIXCHpfepay6aI4CPwQTzdty7VH9a6A5+2bL80
aRsbM9S2mUViSJado6yLx61DLCS1kPItQCA94YksW0NJAr7toH9BiHW7WDkxTz3WpKTDCONMPTA7
ffkvXMygPCFk16uTnegRI/6f0dTuqHKRcFIEqKRgf3lqUHmepEeZUEV/1H2I4D1EpduBW2IhPl8P
vEyzSsIVb2jnPvTzZvT/H+Xjx2MXcgYC6eTM8zvVufuGyEZqPSAVkwGc0B9cvWd0BJvDVHlWtS01
eg5Nl3/W7JI5pgzwpMb0GjjaCST43xZNQT48sEHclZzSwE1cG/jEcV4vD8BNVqmB7ZA9ckPbEDx2
Yvq/knWajf0ZVD08vChpZIbZBaUOeyXlp7is5CZYFjDZoIF5Su/KIwYCvxtH++DahZmyM3UQ6sue
e7QnEB8QLuc+PJvcqtckoqU9e8NLsoSMqXIq8qQ5Xq5tWfDVQy/vYQMnPqT+L2ezJxN6Np19XM6h
srfyAEXlP4aESgJuf5bGUkW967oSbciXRmA0lXEEYUhJhHsZlrMs4paTr+OVVgH3ZvOjNn1VQVfx
q1x9SFVrtwaEWpjyW3gybbHLDGH+BS9XyN9aoQujrc/+uuyPhIaxuoa/3mEjkYbR27agctqSmGrt
k+RclFWbQcS+kP9VrNqRcABc3xjDpkpNmva2XNZouNOcvN5tYIhhp2MuGERTQQCwwck9DwimDmm0
kFu7ZbWNBm5RJg+0tQnHIXU3ASe+2HbkiH1ZY6JXNw/cszNmdlB76I4yqKDTlV00hLJKa3gzTDVz
cpgQ4Ty0ix1OTYFGLD/CYSnoi1o7/oL8tKGbpBuNRtpdrw+D3rsm/p9xfd37KJHWWEBBDv2Y+peM
ZwJXyWls5ri+IQdahG+SeyiKNJL4u6JS51Ap/MUmu/w0Xag4N0l8YiyvjeZwQGUxhYnUxYDmNLhe
cZQNn69sq2rkHiXLn7S+xGw8OsA/A+HTmyquK/qss3SZpNuxKg/Ri+jxeOTthGoqjXCj2vM4n+Gc
sv4STWzl8bizuKPeiY/YT0lp7/5AMIo08G9kFr0kDjqREeJ+NZjMD5l2lXkgBHcbmC78CFzGjYnE
jsxiX2PBOzJrfXyUxv7jyuFOjOFb1OsdXB3YaWH3xhFrDSNqnS1e7ZbKI3QMybvGpvmrNBdj+ALe
G0goV1LRJ3FTWKFpLEPmH4YPx9cRzyD502wFAlEjXX9scrAjOZp9T4mU+LSHOfzoZwVmNTmokNAJ
jyN7eLy263HmRl47tst6QlQ1P8wb10u/degUB4l87Y4Cx5ROBPXTrzcx89pPrAcE64Eh7WbUQCMb
LQhgB22EBBmSc3XMvCLL/0HNBeP1IqwYZwfeLV5GmopJA1z1ezd+a73KOQnle119p9sDna9g2F4X
lS0ajLoNK24nMJlxy6FNrHxJr20ij+htnnByMrPlMrn3MTRlSsJybdVSLjI1r99HgJK1SWNd4xiL
AJqx6awCYVvXEQGAdQQGcSYO7Qzt8cUrq/ZQf1j4l1l2ssML/9MBOYH9zTQgqcO5pONP7KkH/Fw8
JPKwpmLPwqdOKHzxGzAta2JA6sEj/ZL64HLQ8HzPGjDd+l1skdqBJ7N+jrxpuy3Uf1O5x6HqhjWb
JgAYmtAnI39vbbXhKvPsZl5PtwgHJev6B4v7OJpI2nzEPLCSH8fl/urrbZe6E9V9SMUsSfcaQnxv
V9FnX8B9K8rH3+DFCliKdCF5AzySaHsLH/y2UumJVCb4w98vYeIYUm2w/Iipq09F8xmQqYzdq4YN
CcfPB/o3IVRVWP2tKiYN8rT32kzmQJdF0E9qOrJqUEMl0vsBVI9vWaIBxl6JKhJGn6ZMjpzr5XbI
qE9GGvF5t+XOld1GwfmMeKFRbU2OfNikkn2tUAtWLLmoVl9/oPP6KdowmStlcLyKld3xXlbxCFGR
1AWWG+PIh68JQeRVGZfAkPfLbMZyoJWFaOt/uChQsG0P1+jgVAQ1Yz1Fccq3UvRjzYD6bVbeWlgp
pCweSMxVlKZF+UccbnRCDVDBWPYUiKxIIj5bX98aVtkofQAojIi3b8SliK5JMZ8OgqBj5l57xZ/M
i3XJuWajiS/4nAUiOgUVVOIj5vIvZUtR2+4YPnpP8/c1XHCTbztcmOZfl3vDwniGHr9B3o/bkFew
zh/qgZzXtBLcrHHVw3kHhDBVQI+CNL+a5Du9cF3XiBIgPfW1VwW1Y1BdJfnnZlgj5Ffomq2+XMtO
M4S+GldCM65pywsvIc+xu6wAUVQ4WE9WsR6JU/vNKjm7MDXeubWcjXFqpNDlj0Yh6Tvk0Vri1F1d
D6eq3K6R+OXPWiSqAvNKZcoT8folsHn860wJScSbgRnEaOl4MNi2oYyO16kwHunLElxK9cWiYlrz
RIP7DxTjx3a0QbyjU0/lNVD9+sFAAH9XAdDKkDeXmFr6ZfSGoVdKTxEl2HCQzCu3FZIOm0VbYERA
dyk7RMHnAA1ZFQRnArpT1ruXQJIZn66M2WeqjqPIBwGGtTI617CxlinUKeduN6xxeiTSMvFaoPrx
mDttUlUOsJkdfLVDTGOhGoY6Car1XwaUHhlwEl2e9PlltXBfcVVho4bPv+Pl2Fa9LskjMkfsug8q
LjpRt6aLVNY85e49l0uDcPXF25dNLagwRCjNKKdjAap4/eeBRqY61j+hiHSmNmAABzPIXiai9RkB
kUyH/Jo+1inD+7AzVKn4mlS5njDZ7mfjwekoAKbPKKp/CADsbmTxuLo0m6UTrMEmr35A7FZLqP09
BX2jcZ/rWkUe3XPE00WC00nvGyl5GvLZPkuGLhDQVY+7KqVLmW2GMWA0snC6LQPJhCbNtGb2y4jZ
Xq4t7Uq2mtgRTmQ+xcm0YVR4V3Mn4pBh33jhistS1gSwdD6l4hEIP1O1kU4pNIAuSkEAeNjLyadR
P8W10w8Crn1qrOFqZvnCfTFirD0XZSKAxrOF4bNRiBCcH8M90CV9zBD1jOwNRDkk+RFBgfx9WeTQ
0yeOgKEOjNejkP+AIAngY4TOq/OdWp4L80HdiB2otlBQxKSMRozsGScBx5LYQWOXoE9fz9GuLtkT
pw/TG/jeP5nWbtTQmEz/WZAVNG8jM5x50wEkq8ne5YfT3EIR4EAggI63LjYF7vO0ynDX2XbpheKu
OeqYLiG1opss6vQj02ioXUdqA0uUkxZb5j3aOjAWYgOvmsUzTpNP2EEapKrwpjr4avtVdlh2zwbK
aVVHn05+xh4Ez31vJqOgyivX/fkLUGj621rmY2RAyl+ZZm2ZaggK2ELtmiTeTkS1jtfGQrNt8euj
2HYfhNlhq9ozF0gT4Z7ZMPXTjU9Wf23Pqs8OVk4N63VNEu3lCkxbjUQdQjP+iyyxXwGuJZNM3a2Q
i/kZIo5dOtdfNM2V59Ddb66uH7/b9cQSPzF9pzpsnNsXCP2fI+GFpYQr2ZTZx33gm9MB7ZvBtwAC
fYLmGU8N+yQkzrIXrcEFlCCJeKSy4UJIqpOOoxmSYG77qUvoJVpHIKlNPdFaEoY3DzIoX4VFMclx
xFFjXMiImu6jE0AT9h89gA40KckQFiAgzIeTfndU10ME3XsBblvBuiWE4vsnkRmne/3JlsiVtHsS
lUYn0lAGflLTZ55RGM6CS4Kl6HcXlAFu3O4JOP1wbChVBLkP3loAufmJgguo+NSA26KjFvjw0WuH
StFrk+iS9WKQAJseCcAfVe1aMkjMeyB2U6jmYYZYEy954XDHRn7C4m3IU193Y9DUwXPnXd49Y8u9
kFAoHE2ou5j3hqT4hkbJP0dDwOyJ5K4Ja9GceGnTM9ULh6ppm64dvZI/0uOCiYL6qIY7xqQPo9eh
3syyF5oIgXetmeYcrxvQT+TpCEPYmFwksF1oqhMKSclrAG2GiBSYcVTjnRhkdK47AKn2Dd49x3jF
bBua4uzXUMSFW8T6DOnvfayb7j9eMhX3eqDocbF6X36tTJUsYDtAX19XlwaSvjVK8UVGd5JiIkRl
hh+iMf1iz2gqwexcUCU97nN7DIEjrgxVx2rOcusjK0/w3jHJMRQPrJNig9Ukx7yL5DE2RCHq/Sel
lFnzu2zmr+ufZDLBnhcFEDbCh2Q8i0pIjCBuJ87loa94cGVZUPSM3omX832XPv9J2CiYa51n3avf
tOT/F3SxemUneYUcb2TEtYif9hHVmvSMmVJjhF+vDR8Pd9bEz0db5A2AyQKvvKZ35rB56WZE0FVt
NFK+jkjLMlBI9Cbe2+1rIQo5Fasg8hjXrVhkW1/rwF8INKpeuR6mTzOwMYKh8HS2ijW6GyDMm74r
762SFX1MmczEBF1ORhLJ+H18ToQCpnJmdV8OoVIO5lOvOKremfgLEihoVvVTQjyZhGjPOvCGS5k2
zkuhsRBoPpj8Y+8kJgTgSgxxjmCe5d1k/TfVJvcGw8usuL6x+GzfATb0Trgo5keBHm6FYBQ90aQO
0Ii6t7IH0GPIS+2cvjponEqvUwaOaVOiJQwRVX+kAqCY84CEFYWR5TwhxpA47hxWT1POzP23RjiI
9M2qYm7uutL8RLAjx2RrzzR/IC/ld33hiHasVuLt+e42agk9hHvMQm6F7yadrAHTQCvhTmWE1BRD
+VyPUKLWbERLu4sINZ3AMi3deGtMOdPyPDZ2TJQYlRPvy+10d1dNY9t7Qe4ipJ02/RHYRDg10KAg
C9/rqRieRcrniA/w+LLsO9pXClLdLkF4cEVZvS+6Lbvku7i89EEnueBh1KYXkURtzzyBw8KOTejL
EYheTGQpTT30Bew0nS0l1FjInkHjKoHgoyHfQFQeKx9xRdWAKmdCKk2Yz4NU5FD/UvNDGsXJKGyZ
/SC+K9RmbdKAWTAQ/zh6xL2D0TkK9gk6bd5xCE2Lp+b6bvT3+/v2XL+ktsy3tGZ4QsC5+MQ/3r10
5hQDpdrU0kHy9d6frRwtU8tFhfGTsxYNeitLfTLZnEBHSV93qAcEI9hE7bjFpGWNJx/g83uh5+0r
jsgXBSfdXZ26RFfU6SPzPXyYeDUL6kit53rvs/7Htw0860YBkkndcSiOAuYG7xwJjgR/nT4QHF57
H7Y35RNtNSGfPG77vXaxl0Q3PqRkkgxf8sQtvZX0z7LMcdiwoFBi/onbRT4RqUFaECONWqirNRld
1Sy2ATn/gAFs24o1PuIeLPLSLy995cLVn6507dVycbLG3wpTSK4IjIL4gcn7ua5t8+ngrruSwlOG
aFnxaLLii6/n5tNd0Z0fOuh06pFeeQGooei47QdoT0z4pgBr+4wc5DCPre8OKtq9OnKaGufd2O9b
CdczMUXsft/hRCP+TTwIVH66OQWYYnp/Cbap7uwUDz0CqlUwAz7+GP/iWiPj4nTlIeRVkKnArxmH
RFoqUecMS+hAjSb180U2bsQFVgL7B6CCXXZB9tbACkltKnjhdkt9k490UWeF364XhuQ9daRQ0Mqk
Labsaw7c66fQbJB3XaZHfuLad+57p0tA9iuTx/ANC74QwGbjsicijlY5g9XTUYXa/lMCaZWNTWxu
vd20j2NuOTyLXiIoF4iQYZRGKOpYcgveTWuDchFugn2evTNkhesACYAAATfkNKM4N20TSjIc9Fiy
tsGITQInTwvnbidWOiTKCmr2kmNKl/cWXMQse0zarugc5XL3Zh67fN5h+vMJB/t5VKE6J23nikzF
r5FDqtObmjgjuubuNa0OZw0ieJDXgbtjwSyDG6jYvazTXXQBVsf7KbldQkfuTJhBWYe1CG4bQaRx
RwsYrk5onb8akMaZ9s5oHW9hGoJDuLsDYazjdggOSgPzlfbrJHKzyg8WCTRE5RBrWuOYLG0U9SJl
0zICtKclw6LF3oN4ATUHsla6vUlIurLCkB1K9KC1lvun9K+LQU7MocyAFAdRGKPz+hB1KZ8vV/3v
3M8huTa+ghiqN5xPDCb34rDoSrtfMelOM6N1c08sTDE+Hs4TPZbJW+pHcTatzgopKG+Znh2/MLAc
V9Sd8Tw0qZB3Xwn0ZrMRw1en5YXJ2uK5Dzc8QGhkMcczYq3EfNIIA9Cm47nc9nJSA6sNAfznkA8u
PxBOzTgH6oVBlRnT18lt4hkau4k1YH4OIMZnbH80cISijeoVWguVcXfXfb/RSnN+MUlqZCEv7qFI
rfEqrdaIRpqwafQW8KXaMFlWn8q93xs/Dkk4leYxJIuGNP9XGKyFG6ghG3WxIlxfVjC/G6KLO2pi
qfW/RC8itV5cWwTSx/UeJBq8SlqBmWW1BMRkE7vVcsuqVrSGTw0r6nVYDvwM8UlskWuQiKaHA2WH
MJhP94TQuePkcd8cPhbv7k7MkFpJLqsMwvjNRHf3YprYgRkS2nauY5WW0cLzChRG7MfeNzQpy3yL
5DZqNW3pHBkmrEJgqbJ69DHgNYeOAEYW82poulYFtoRbn9fi5gxL1hWv95dRzgRWopV8X958/ON4
FYX1sjmDy+AkUtLgsOwmjNWet49ZrIOFvlMkE5DF+ZzvQHhYYf5F4itRT4VnfD+iRs5j0o7EdWCP
yJSD9tNOQ1nMd6Hr2/9wpaQxwE3vQ8MIKay1xAtb3v5ybLr7KGpoQ8wiq/tOCOp4iPexiP203nSt
FKhemyIZBdH4XDqUXy/fMJZA4TL/k34RoYgTIVSp8V4c4D/PqL6rPJNDZcPo3luPiPHJhB/gOYdK
j8ddEBChwvux0oa5dyGQEjRasc0R0GoZn4oICWoGQTrJQEk5SbO9pfJ8uODbKlPEJBSw0wAkNw+0
H0jax88iCcNKw2qbdMrddGeOgIrO8V061SmhI5Vas8oYJctgObMokWKLHBd3WBBxIr6C5Og7WD5B
65IKQNqjfB6WHyORgvghcWKlgk93kpsaQBJK2x9RUdJae3VXkYN67Da2uj/Hcm7x2g5Sy1pN5O3w
efg0eldpti4cLmjAk+OVOi7yTaC9KhMTOk7WMIW+haLhwF4ufHz6jQ1yQHvAfYIEDNleSyAFQ2rU
zFXkIdJasZDPYTiVljG3iQE8G+yfeJC8NmftM8z9QuHwAxHY358TDl5DQq0WnL1leeh7SP6PNcQM
ssMYoEOx7H+B0ysiHFexJR3scEOI3Dkh/pvSGw6u5YAeOa1EPav7bx8bJO+PPdiR9k3bjEVx/xUE
vRQzgL0bFs2UqOrXZpKv5S8QRCgmnCMfdD0qOhMHhG5F5KMgOO1XwxMzo9yAQ8nao4HddIcsmn5M
NXYQ+yTTbZ0fT3D4S4V0n9jPXZHQK6GEVz3Dz28mdBHxPTr9MJBg9bUHOrPfphiIXzKS9xru7Hwy
BuhCvB0jivOY7Amd+9reqb6b9JnB8P5z1X4nq8mEAgI3UTfY5Y8CVIBj2E2tvKRKaI0Ba+3VczXe
6/24Zz0u5VdU2qzu4o/5CH+RgloCehJOpIZzGmtgMIDs7HIX5ukMHTYovLzQjEE0o10BFABBZDHC
5x1cqDCdNRfOwzpSxqYyQs6z+TyrO7PX+IKcaOuIKcvmA5K6uDUlUSjSlgNSuUqWJgj5XlM23Upd
lLcFmfmHcTq1qCJlalcQgD02zFEKNUAjWKKKqkKOS3njW3N9eph38WjsonGpra140/p/lxxfJji8
vatZUXYJU26tPYPHU5tLWMiBzdcQUXrIbwIoojENKXmLxjrtpBUABJykOJD4P20A9m/uH5fzd4aP
JamRLiY4ciO+YJ93trqW1WrnSSmnecGUy69vIuYOynXgp/IAojaIVxlCP08NjAC9uggMDZWx/f+I
Om0zK8G14SKPA/bnS2/pLEtEQCHgcYXqaouSCWR5naAf3Fauz0jCLwI6R9e0unBnksTDh+DlBBWs
Sg3LZq8A//62dBoCcTRRuBdHM5XBG34tNGq2scvyELcxw0B3Cr9BezEMOV6zB5JoXW8KMTIPBH/U
SZ4gLYADd/6vJKASE9ZQqcd8QBydNpjpC436cXFm+KgJm9bXq/yiIvFQqsoXqno6us83fXIWOH54
+Gp13DJ1OCVPThc4ZGYORHr0TfJekZdEsDoyYkGWTjuOun+qRlwtaSHwdyaZasQHPU0BkCehQgB4
5HkY6cr++gXhXXEUlfTfu0pKFSyVBPhEl534RCtTYvPjQ6jxQ0l4v0y/Ucse1fM9Zk+rnBPArb/U
reZB9v7AKXtzA0BkLp8Dpy/JXVfWcn08zPvhRkQC+mmCDS3vDYPBGqSHGiwKaiN2IeJ53RYOD/+D
es+wikS6Yn8bLBJRM4kP67QcMMLVVB52qGsCI5hbZ6M6T9BSt27Ybmg3KXsUTLHRYLkYQ3EYOHBC
w4NJ/GpgaTDGz6D71u2ubG8EsGtJRt6f2xcVIzdMKzawhce6pDXoHOMwLl6/pLYtqNsBRNC0pC8G
SCdfmJlAB4ShI0xbgzNlht9rg9qlXcZv+i7AS8nB4qSdfgrCXCbe8j1iajO2r7KXGULJMapU0yuL
1UyuaeNSPNdtzHUwFvFdWYjFCDNBI1gqCH8bj7L4tAYIfVn1858apARrFHr+T3zRK1hZGe2QzRVf
ao/gwYvFCATWlKb/eu/qsj5Qv7E14sz7NLnZuq7EHexTcRBJlrDP3aTz2nWhKnOnH0hOPBxhxi6A
hPFLPksDQb4uQE3oJnolFIxZIGOqF3M42ws4JJQQVmGjFiZc59IqgDOdYUfKDjBBmw+7iHBF/V2W
bZhM7GfK/6ljqQXKMpQCif/VdFw5jRr1pISFrGvz9QUOMwNf7mlVOVkMxt6dU711DWVXUR7FhF5S
/KFuTJNvgYxgfhHBvgT820eh/ftBuiD8b8/mndfeUOrnGJmbNmXHV0qs+Yjtwp7cU386Phj/B+xs
ebN3fLnat5G0vKs8UnWknWrZ+zt7xBR2A9Or77FuI0Pt6UvDGVWeg5q+y1mI4JLS9g2sbVTIuMBM
iIVglbNjTeRv8aXZ9/DsRffnQKnW96viX13MY/euUllCFpJcQrPalMybI+QfgnwvWiTtbm4hG/gZ
07o0MEYsBZY6GfRCa0EjIwxVaa3VDOYGXJYSA+UuXKy87ErDtza4n6vp424wug+qs7q45SPh/KCs
yqeI/6e9y5A0ezneaRjeeGiIkFHsMO6DjIBBjY1QtoBRf3BRCSb9LZwb4qsfV4FO9XC4/fXEG2uw
14LwPu8gJ6Ah4UONrgHB+vT7XDXgAG2TolKzFs4FKah3OeCdi20n4E5jEUDNCXUhUET/xkuRwDr/
NkkD29Z6taKf2fSVTw3LXdtcE24Jb72f9Wmv9JBisvfelcmAPZd2QOV070YTlC9mgBbdmT3r3vmB
2qFg+BSNhDrB1PfTBH8gObHD5JEUUrmJAI5sfnRT8Ef0WN/72RR6+wwLwYzhj5G9ntnn4IVVEyBv
cBmX1JJ+JoSpFMQ5WE8XMhqQqFoirA/jo3yWdHPGDKTDxXTkXtunVmJQumpEZE+yX7ay2LPK0hVu
sz/NazpxdoF5YG6QHe97ux6SasmdobqjfVhN8/hccwPgL4vambFGRzpTMBHxSP49mKpEUR1IhGQj
J6il1yp5P5uAqwwen9vjjtYwQLoJNYC3W94J2tVl+gqhs9aqyFCVH7mWs7iUZMfQBxy/jV5jUztL
6u+MS1V0j9SBQf0THP+xPyfZMfYd9v8pHVBf/hT5NyKy8ZOk/L+GfqSYvyLj8QQYRKJXUTZmsn/4
SkOZqauocgsukwhzAkimp6UV4pRPbaI+NeGkN6ocg30CnZz9S+vxr8uyFFRo9ZpX0BF1/AH8myRn
90Pz9itJKObnZA8c7nzAz0Xxb98LJd//iKPEBzx6LJxit+epBijJf5ev09+jXghhpsnv+C9tU4S1
GQYeJyi1XzbCkQZ6xguNxgUb5+flGhdWlGqxY7bO1WUpdtFrsdC9HBVYAb6by23+83TwD+2wSrRh
1vKrLD7kR77fpT1b5wTX7eUUfJnKK9Mard8V+QEhLZ+8CJRPqD5D9afXTPeU06NSjXXdh1z46fjx
ft2fvdsC4MTWzUK8kjl+dvbLOh+FFI6XiCXsS/NsrC990zQplqz2VsGLi8+ZP6NUVS5rUFw6+UmM
kCzg5Jg/Ou3YUwLf26XrlnwYDBuV7FJQ/tAOQ3OogKdE61PW04wcct/nL+Sel3Bhmq8/rtJMROde
4HmUNk4tzq3KEFr/cuWCpufJjC1lJTBg6Dle7R9hQl9Qm2LcPRU+9OVIKaB2BcaBB/rk96HXaAMO
s9S9ger4z0a0YbpBeDTqw2k4C9fS91p5LGUggeo7EOhuNUzDtb1Z18lb50E5yqpVxV0CSIHB+ciV
EwjS5b+nNX5RA+HrJ+FKQMdvfIxbfWCHSTg46JUXMoo1L5jCV3xfez3Hs2lbxovo3NEHuR5Nxgj3
folZxd085i1eT4cgqJS0/F1gSMb8jcd5sowQIg6aodOO25OeKeujpn24faOWK2Tkv0rSVfLizsQv
dexmBoQLpj67ErzvhwR3xvZA0kfT/heAtVnhbncKMms8LM9B/nD4nUGYA1Skujt+b3rVbC7V+LR6
C1ALiQN4J2+qmlKhCC8zyFHWRrG279kV713+nb/ffZAxqp2q/tVYMQXwACdhXPzxHBk41CGVyCKy
/Lrvqvt1rHnSoRWQs0cchmJ614gJVUMqAI2/NQUxkUGfgK1zkZ2KJYvS+in8xeJTAcI21ggTYrEA
JlBdELH1ksXAfPjdI3W5D+3yPhmfYyDih1Owr4Ea/XAMl9n2jHdMRN4B/Cru1RhQq8d1bjZ3SahR
vmVJ0czKoBsLbQd4EgSMeGTiwuMEfeSma3f52GwOtBHAYpD3l20lZTOtiERTJU/iqvQ6UaR8MFk6
97ULG7xt5zeQvo+SNcSVBLH4RQ7SX44iJmsqISU66MGF1MTjeXMoRZ/DqCKLqbJJi8irOGM6Athg
daYeRqyqnPTLtnh/m11WsZ266XKfr2vAFIRPDhQkQ1gQpR7n8e7dL7G+E9uE+qj9kqvl3VTbmvq8
0Av+fRC/QY85kd8ATEKgmkgh5nxPCoucyDWbobl/YKYsPYn/Mqq+zOO/cPAxWgNDWbZOGZnFCujF
BgPSwExgIXKmN5dRXhcIv+MsWkr88pdrzTIiU/ETSHg1oQWkzrh5onFVHf9XUbTe9QMVOuFQlO4n
JAzaWlrSP9pSP8iDkw5MLqlGoNsAt1MkbfR7IbteQKEEvDyMl5vEPykpSeHZeydTe/hoWXG7AOpF
TGkPbVle+APiCA74fqLI+whmQ524xKO2fC5iX58nSwsdessw1L/N8PnO9wv/mtPklpZcx19niOOF
o1+tXWeMC/dhxgq7B5a+Ghb7kmMYJymqqj9UUOZtauE9+NzhEWF/5kdCdXVNYl8PfS0Aprqjmsc9
JATe0D2YujW0kWDwnpCYJTldqppUeekCM5GY0ZjDB8vWdctTNR8+uwYCvoXHNY4vDYyy+sO8jQZC
6ZytuxfSiu7hVThaBbk3zByxT6lgUpyElpSER7nf+xTsKb4547QY3hS/ql5wH4XYJElYdZHdwbqD
MjJ39upF7NIu4vjVVB2I2CxBeP3Qlyo6EaxVSEMXSoLJp9ObcOK3vdJkcb9NC0MuQ7Hn/FG/DP4z
fdFJo/VgJwpKv/JnXwa0ZRBp76q+PldQ6yJfYvGfxbHZDmquJo55aVxrCGOK0jdondUEtPNXIThP
N/rUiK/FVW0HEKXcner01eHTu2z7tSoGhXIg2nxl9CSk6qEIdzjbgocITQUEya4yo3JkufV55woz
H6FDQu6qm5X7opFRKQdGDCmEAlvSYL6vM03z3ulJWcHdfKCyMm7T1sduCbE7cxlWgJJLx7atESMO
oL73F6hZ2fj54G8hLcKaxA5nhuuqP48XXg8jQ6sZY2o78f5KDmBD4o22VP3KZHO24xkC3WgCCgIY
s+ihmtSVQYtx4r82co4o6c0DE4QJME3BfUdt4T9wwImr7Uwupk7LYnUEeMKzzv4uggnRbLjQ9zDU
pzfKnUCf/s0iz1cd39ROEoEBeDN1fo+dxWNTmqNnPt28aSSERFkgMMp7NATodTEyhWNEPawT8FVM
9aXHh+EfD+nysVfPPb/XqH2Scc6oeHrAxO4o1u7k8TOjBD7wPbtN5Go+TWiFlnhISxlR5GbvX/vX
DIp4lutGuoGxc9siSIzB69ZiZEvzZ0YLENTwjLqxTHqBSnU+c2/V6l4dAuyIwWV31YcbkX7iLFMm
agVCB9sIV8FU3UTir7bsDX3wNobJ8Mg1j0cL/tGPoisP1H0/8r81jQG+GKNgeXaykEbk8m9UdKwN
p/FyLqqKxldxjx6ArEdYSKJbXEUG6mJi23Uj3oCpcLLa7lTOCqRJjbUxYBba7qVqz/1vPVpm/EHa
CmwAdZKOGD5wFUw1ZqTyWjb5U5/aoty9K+uOO2IzciXgyEO740WTCCOdseUyUI4hpoPEvmq3oKEs
+74epvt8q8AmFHq9CVe7Q/Z5brVAQG4JIg1TfbwnYo8KYbPytgpJSD0bftiXGwxWBIxJaUvZWhar
bdAJ7zuamuW3nfUkctfDQiB9OzgijjSiCGzf0u1jqnOOvXO0isCWpgOWvL+nZnI/OvidUWeemcml
psSB1rFQveA88icCYGM8icgBrTjLZowGRmx9EjfaqbA1xq8HfC7dODcPGqHTFqnuXWn7DcKQzxgA
PO5rpbEPIPm90LzTdEh/f4H7ebj11Wl/cZd5dNwx/n2RnsNkk1yPtjGLBZt8EsNgqvt+azN4108W
/Pw8Fu6QlgpxFMimB7+QlimU7qiD2gKXl+wJqCmdWcI8JugQkji5wt92G3sa84LmW8ymolD2PPiQ
OsehgvEXu0APBPnZxMndEWR9qenrJdb5exOF4HVuXVf8AhBX0yw27z8gE6sYD+v1XzveakgIYDzC
LNt2nqnVlDvcWs6clI3a5KSNB3l0hCAGkJW7i+s1vaNn5CuQgU7hUNM563RcSdirwxc2i3BhTWoZ
CQ9k2J0D0NsUVnRBP41HOwcmf5MIaOD4P4XMCtiWSGPHi/FseRmtwUtDhlX/Ynd7QT8CzaNa9zQx
xOoS9dxLZ8qp21qno7up46u5v+W0jHEtFNWpldUSoHV4rZ1Kqn+Lif7PpcIF3HRbWXQUUc1/Asby
7PqIEcudi0xI39gG9Ml0bOlPc7fmQUL9xq85OLN9p2JFJLXK0+oqCyQmz8TbtS9vOiTid1zpxqr2
0rt5w4qqaqrLpbmGUVFKCYJJtGkvHy7NKMJDOw7gROb3hY1BA2s5qYaX1VbQlempMFpgsZwEQsFt
HgaW6HeLpr8JAmcLUvSth3YianRBwW5ItbHu4F+dVYJBPoFtkZknbXxdbrDhAvJ5qp+KRusqWJ4/
t9pI5Fos2SCRGSn9tZM3gqdxGFxC7kf6p6LKx+Giupm1P6IiFtsI2CxPEVVpQihgExdTkoMNreca
7+vj9HRO/mT/ESs+4sjdMcK/4kkPD5PuK9z39vLs8NG2VP3btmf0xTPmzDOCgBuk+wFYh6pvykS/
gWzGxCGPcE+HqoVN4Ex0DJNYbMgX4YuJ7xUvK4wDYebHGgYvGzCSgI4u76CzLw5Bo60KKLl2RH19
dd3iqArIqFvMxdg9lsQ1E01eP+1BiqPZeFL035ovnD4yRNddHr+qJ69MVMJq7Q/MbNOffVrr7XSK
iXTBOqgkDyqFaT56mRgpjprDfXdxlALbCgXmILAPb2nJ2QSKj9UjwvqOlNdcKc1OBC6/TKYFdXdY
Qj1jXLEX44p+0xlz5m9F1JmBGXcqGvsUud6hzxw/GoAHpoJQID77V9ctFVp6hT1rSt/Hq4DW6FTp
KfIIi1Pt44sNhHHEvOjWGwYdilmzPU/peORZjhMh+WPJKBcL7bxWWKMvz01k2+3qqltz4jWZUbMK
8q7c9lfBQRXjYbSCTfG2NoMMVnUxQUWBzodWkWKCxuyin8r2eyLOXTC6fYHH0RHtlxEGLi5nvB63
68bj44PEHqGniFHmSMc86kRuATtN559lYWhNRSuLdH8q648fWrex7Q3ZNjnOfP1InddWCGPvZ5HU
Ks20C5+OivON4vwHObsba4GGhozFxc2v7Y9GBNFljFVVoxn7MCX8rD3dYJNsyqsMRqpvp20DLNoG
FI3yeKmRJA1CCp5cfjzEd39/NU2L5bpiuCiFBSfE74xIz/G6bSTPSnQblIKN511/6t2Os52w23t7
vPzoL9CaP00/EJuqznpt9F37w60EH+rSwZlm9T+IXtXqs0mpzcdwGf7iZArzfDZg6dBCxycs77QN
PUCuGTzLTSGSmhnD0Fgwqv6yMm/BJ4ocbsV2MFnjDsabr93v8Xqg6PXAYfwKJG3z8XhY9d5rMkTo
DmqNcvOvEVSrQWUmUP9jaGYu3XjDH5U43UmsJ7a52daMf7kM4WAV6ldxyu556SLknhrYAfkUBF5I
ALIgOon/0Lrjpdlgkf4trg8wwcBnntL+DVrYePXAo01fXD1ZYQYTIbfpfPNayhex69e5aHpuEuMP
T/JCsuy8/7zmYRZNJj77lEFj+oK0IBdWBG8/FHHg2vdaPiu22AWXxbx5ktqWfzUKsk3edgiJR/Uj
ARY7Tvcg0Pqg9xWQNSFawznWjFz7D31Wb5Q+uGfX+heZfWGeETKFV1z3NYttLBbG9ySSq+vHCro/
G9cRV+KZDB/hmTCeflefKYHqmlNprI0AIatlL2LKAMJ3/wDjfUp3XA2E8XDoF+ipbDAgy2v9r6qs
vO29hUSzijxvxFXNzOlQ29upisGxv2K0CfN9d2J4FvR/cwHEFb7pEIVt5uM8Hc2wr8V3doxHhCGg
8eyiHoyNtL4btPgXLzeoVasyJyZtWXN+y9N+gVQ2US3X8m5BmvG4SWp+73rCoelYTk6ypmD6drYF
sTy74SzHcJ3xuXMrO9ys7nDH86JnxSOJRlEzIJ2v6OpHCKgRkdbZXpOUC9to3uTM18PoQwd669hZ
qO//IP+GtGt5ecE3o9TJTOc1dEl1S1qf53tO1XQ5xVcGt6ZlWcI+euY7Zb2ilZrkRsTMwFrPIh4b
OjOPwcJBdVaTcfycUUXdg42fR9VY2rToL0s+JIlD/ZgAJhaYJowCI7lRzp/Fxf+uN+NrAFIvg0hQ
VHd8zWKNw5vva8POzz5PpWz16eXKPj83c0J8C7E6v7hdKzycktSx8vMIHEGKWn8/Ucwwkjg2KCZ7
Um+9r10Bih0kbpoZaYupdFNcZRJQbB36U9KfOqyGlumSrHk5dk8sWCIM8+bLLeer8VPnoA/878/g
UWwiixmqL+7bsrOOhpp0wwRpLAmtFETHmenrNMhSJTIVdCxcOlPJvMebxf+T+ZYWYkcRfuTK0+EG
SG9ingYPxgO4ouMgJyPFLI1u/WWihnbGEuhXLDV/PHAfixfdusI5ATN4lJYARtbGytqJ1jjGvixV
gOCevKqNJdSaREORHExrw0PvIrVnDjzO0JFS2ubYEW0OLJ0KZEFMgsz8SWN0znslUFgwby09h/iR
kn4wfqFag5OvkeQAchIY75TeT6HxHMEBfOTtRqE8SnfN+teWKrVhGqtqv0I53lbknBXYIsGmrMa5
Llyp6z9IhJy6e0KJdHrYWbc3ftZWuK4tHev+bS6fIBKZGMXVza603k0qLyF16ooCm9RBz5YMjZRq
5njpNhyQm4+HevOHWt4OMDKguCYmM4yihHeinIEhchXii+UXOIWE/vqYVZUBLoA9YIsN1AOUHDP4
UBhYfQjq0p42m26hqh89NL64uSU12Jibj+yIcmuJMsR3gB2gNtc+KZhV1dMW+JWzsS+t7mDVknRW
F/9cOhm6884WMUpLve6XaZWQbg/SscYvE6ES30c9LnyEbNMPT1RdTa81WfFvZiWYti2s4aGbKosV
52DRmEhcDKfS6wSiX4+s+uy+mPJ4hCeVobGz7xb4MgroBe91lbS2wBUPoUAj0ZCO4IezHxEMa8PZ
glPmxTyanZ7h20h1mTx6rsWlPeeiXNveYhc6lUx/+6aGhXp9t3FA81tlXVGpe+zyY635duw3Zmmg
u6wxzimmBXt6UPREENk4fnVClTqBRwGN2/AT5fRWayDLKQsSbKTkxqEJfvtjsijHRX1I4p/TZPb4
+pvvqYkD4A42i0SPz2GBVSVGMqJBFACCoBTXfhw2VWIxR1f4CzQ0yijQJg35Qw5YoPF0yJFCWSlu
VSLol3hLcsg6LgasMxF1074aDnXU3vpBCX5hf0edwmlAii81KgXKGuALsRui3uN6oUIXWhkX+CLi
5lHy9GekyLWxoE3dyJ9RHDZ/wP9B9ymd2U8z7bThcVtol0RG+9qZUdUaWmwRmUmJQ6PVHsszqvt5
GLPDPo8r2Ll/L9Jg6eBJ0tdZLFf68KHNy3x+X3Ugi4TvOqsPMSB8r9M0x/5c366qgkRSJG/Y/XZV
t9wITVYX8k+2lp/UrUKlPc58cLf/RPcUrVKtyJR7laZJC7LpkbxxQQ9Xk27CRIVbqwAFpCsrCkFT
7HYwD5axjk0R6U1eJHkcAxOlda49n/xzH9kz+inYR8R5JTOttE8+xxHHb86TnX9h9HSU3/YrDDKC
n5x/sDIWig8PCy/sPYGx94n4SgV0btlO9Q5WJXlC0f1RJvgcz1cyDSf1ESB3W5WvGeFgbff2Tji0
DOj85TB0LXBrUpXiJT0fs7mvP3wihUOb9U65FWa32GIMVpE/sXX4SZgzAYd3h2wnP6ZhRlLQoBbW
y5ZTSx2U+BPtsWOWEprCLdeHDZvUphsF7M7eUcR9CZjasikt11m5/k9Swi8LkK1dKqxQIqc79Q+j
B8higmV3qWAOYR1SZcc8KOA2sLqYMaDUngtYmfP25BG40ulfMSDv2RZ9gSkP9mUwApg4GrIQ6xg9
hNFVz+h0OMHarI7zJBqW9WCUjtkyu2PH1bpsIv2Fos0wRzwrhp5McDr4GZhtV1+DlAo56rnh2XyJ
k4M3CfNLJ3qX3EnFMwSJYc60KX25CfuSDr7cjFnbgS4Kwl3g9NuQNVOMJRazZPL7I71KtuKyGRaz
lfwcedV6LVf2fxFe608Lf/qwXLO2J21J5vqHD8NNebBzJ95ppzlHSH94y/Ejpacke0PP7cZtjJd3
eEhGrLVxJ4yvRA5Y9sFCZOiyplxe5jJvpEGcSoGVFXJqE8bufuqSwxHcMdnhC5HPKOHlIOmo3Tgb
8f1y3GeYHsm5mv3InOxZFV2/EVeGhZaMH8ikV68oVCsU2rNwW2+RWMvIhMRls6XXkFQoio0PNYUD
8+rCkbUcDRAyAb/3+NCjhOTbEeFhy5PW3/RwY0n7gAztqFbSWGimJsHfN8AsI6k59UxzertsOY9Q
IhJnVeuDNc8dKW1XJcRwz7iRrjhedo0a0yZ0Pm+x1Xa4b8gK+lz62IQ5naGHVl9oY2gbhKp3B50O
0hdBTODJy+YUtJ9bJRf2XFEf51H3dCjy8gjwwRKJX8MvHGANBS45K0/IAVo4zrTM2I552j4xpNdu
MWYDODOjybH0rjfwYidjIlz3qXztPWU6XgQJ/XZYrmWwghzRnLJiZNlHT8OH/jDw2w453ETLn8IR
XHJhlOoFah0KTh8PJBbjijcHMyTThWdGqD+p0A0OHrnIJQQQTygMX2Z4INCCAd2PbM3QEw4k4fnH
FU3lvZgPpQ2+j7RDQvkH5Z10zENi0ydOn+dSE1Z5xP5W73XcWGMGq2IegXjiBYFPUlYTAcSPT7Kk
uwWIWYXnBvp0UtqP0sNfXod1Ov/kMUpWEdSh5XzAfzSltwnIWk2ZgU8Oe9PNX4vR9Lqk2+gmfISY
SLHDDNH58V8m5ltrLy6HsNe67sypJ5/4CAIZg4eRi5DtsOnhkXgmryWJ1PeNK3+rNFFQFE6mGLNY
wpfvHDXF9h0niqZuQDPlRoMNdyu50iG5KlmLuXXws0P9TQdvAwhli9FcOHuyzqwMc/MYcHkywn7m
kz41k9WTAUhfVQpvNHCkkDayqT95B7ePES7AIrFPayZYNC1pNA4lXeDy4Q3yZikapEKlifCbk5O8
dqZFu0eqRqSCUJMY5OJpkxNgl+9dpTusQIToIGmz38MAOL/jWUx58YICfXRoIXc1l+XrZl7Dknkz
I+h184hPmLPMXlbTAQyLsHyVdLlXJRod5t6iM4/AQr0pQP34EwAJQsUMJRcuWmadiYWd9crJOyFU
yJYlAJ2pQO2SQpGeyrE/pTmIFBFP4U50u9kxp/Xa4wbFaPIIr2DIks1kX5M5hgRAHST7PZK5o/wY
k4K3Oe1nTBj2NcQofHjkNrzCpRvCLh7g7ttEs+4B1BnJbTIfBXgr37Ma7RoDR+yCYYb2LTetGOuS
yTy2m3VG5RQuF3G8BvNJwUCWsmj0Cw9NWir6W0fIpn0ikT5VxQG9BH6potNLD8A11TEeBWtluXdv
Jsy4C1WPI/olCGzDmzhwxeHP5U7c3Nooi+x3RrNtOELcrLDZvbONLOPvERal+/TMjk2YwTp/1VOg
Sl9P3FJp8n/UlHBnGTmhNvk3anrcgCc5LAqMho6fV6cyLUn/eqbhT5k9L6F/OMMZm/hBH9uiuLpu
tBujuDrZAeYWGvl/QPRHpa8uw14R8JSubfXY8VCKb1hJmxlCICj3JhWKSHwZmxbslN6aw90I7pjz
8ewDHZmEqrpT8oIEOutR3izhzhtvq1cCUzWqdPV5uyjB8/2ZZJB6krsmIVO5VD/KGRENt+lL8r/j
Y0sQeLoaWe9rcSLMm3iIzH+VrFOSniLYnoDw2M2mT8Ka7SNTOF2DQuQcm7K1Bj/qV4MYXq8oF0QT
gPTYFnFSyhFNFbeeI4U4jFtOWs3GqKcgQdhbxB3FbTBXbBhvWhldy/ifIprvL/qx33ylRb9hP+co
cP4egk8YmzM74N0nKzcpoc4Or/vZ/jzRMtnkUQ6IXPFVF2CQf8GghrEnjAT7JNmxZlYJPYvBsHbY
4tueuEWg9J+Kx1mwj90BBAismkdqYvzE8MzPln+MU3CTe4KWemxSEkuQnAT/jd3Nq3XWpUjDQLjP
Gqp/8kK1eEGfDwGMckVZsnP2AGAtCEGhkXoLEkneR4UPCga6lFmwU9k0Bae6FyDI8CuxAGmOCHen
MBzrvQrMxZY3Rr20n5gQmUM1q962Wc52MjAwLZOD9/It6EFoMa2gROc8hPpWpx/1TRczhesw1s7j
tlROojUEznqX879mvC8/FEw4YXRjBTiz2toMpCgBSTFcKS8UMdG7we1dYLlpV+2niwFlBm+FMfpp
UmM+L4PG+3C0qR7i68EgkfyjiQRelz6NpvXiLoQgTosGUT9HFvD3fHMw8ETbqk8/q30byuqzlIVP
jNkkDnsPFfSgUaBkEnlK/8ZoJZlzJa3oZC6gSQVDA5FCliPbsBKEGU1eBWtNB+O+NF6uN5rDf/6F
qPV7Sb7XbvrojrcSUTZXPXzf8ClpDkDMcxqp27vrUREFBexUfx3nuR56hhZRwI/1oOgcitejSIge
3OWWOyUtCdjcmXAh3ej47UGlFni5E82zDCDG64d6d1i2RmyEBxGP+2QqQt5kcvorVkNWluflKzsq
IIPkEo/M4LQuiPBqX4za6qhDWR5S/AADqtTDyope9EfTeQ9aY5qOUw/mbYqoN1e1z0szD+D5EfI5
ZJbar62h10u1lXV0tE+CZAcarX7kltpn2vCIdTtcFyjvqQPZYXI54SUWie8pJe5fhpNJarHCmhh+
9YlfSCeLVJ4wq2qDFSnmSOpZvLtUCFWfHocccdX5JU0YkeiQL43BqsNHoZ0QQ89gCYW52SnXMife
MC+OoXD3ckmYHpuWsRP3rWg5bLq/KxN+NiR+V1FasVnueW8YOof0WU0n5wnBs574WEYPFxp4xLgH
2VkSozVlC5AJIdoKRGPSLLdZTgsuD7xhn4bVpr5Ub0IRzqIvQPaeb2+f8SE925XJE0Duo/EphkVy
YwkwXlvoUPRHM6X7slwJdYP7lTayjnEgeZTJ1/gkBXdZpo1kE5k5gk+h/gZwD+P2AiETrYul99tJ
tbR5t8GBXeT1wWgfCX4AlVzYhSLXZtGcuL7Zj3Kv5vp+tydKtSYVsrqK6LPisJK9iw9MDvoBxf3S
jBuWx3Xalfvfks/gncTVRzjIAgAfdMQ6b2jrfN28BV9T/ExcB/iFYTchDiNUNdYo351ncs1ESmey
8dcywILowXLFncHhUKr/isq4F7iX/jioa77mecIyrurxLfxt8wowiDr4RygZxJEqahMh1npXlFNC
AsMlsRFDOupQmtnJf6Kli6IS0SbvBIPtRLLh1XYHF2Nn3tzmPSlDhyNQnnilTXMyJFvv53eFK4uC
TKHdxzBMyBT4jJSqbOgN/LcCM2+ldGqnF0fMyTp9y/5J1b6Qr4ZNIFZgr69ribEeXFCscONejy6F
+pk2ldtUWpoaj23yqdx011/sEqB7poFfRpWHT3jIKNBYUr76aS1UEqYN0RBoqcEfTPtIu1jysTqX
TZDdv7ZUe+2SduDd1YtorMVkWV0r24WQtulbXnpA7mP2kI8Wx5CZ7aNSL0qX6ULcAcekHCtyv6z2
9/mxju2IIr/u4/OeQyAe8KS6uVQD4q/sIG6aLGjpl3yMX7bVPbpj1m0Jy0KyfpvKEBeIgD1TFyeY
O/QP0ZoTy+HztqNxna0k8npo7Xh3LqGAFkFtq5f2C+7hBQgJSHzOWZSzlsL56arUFqCERqTQc5LV
arHaWpqjRhf+rJT86rmL7zcGR+S/AgJ54fAnUcvP4kC3GTUk3emwJPD9JBu6rmoVDsz8cUr1hIjA
T+lY2lVT+h36oBsj2uNNcBglnsgcvMjsXP8P1XTGT4CbxBv112TI6fk2E17T0r9Lo+koVq40P8Jg
31k41oZpoZ2q3hsUZ+3bZOaUtqxCKwT01bHFaO7NsOm9oOJk0jh8f+cO8+tu4hda985sdbxOVeKt
p/kj94gwHQfOdmcsEQiccvrCXwvTsGbg6dkPBETx0tSeRpExVcrWj6wsz8KPeS2Ldg3cTK2/HFMz
C2HP8jeSypd39dV0sCaUwKvxLcMCtxQqyS4da8dhVBQe6Gny1McgVN5cqO5H/4DvZItyvELwbumx
WcFSqg3pU5PMyDZBYQ7tuHj0PP8kTSt/kk7loex9uaFkEw/G/+NUXgakxnp93nAkEvrDHEyI/juK
+fxn1v9uPYM5Q9tAVngbQ0+G/948B0kwJ+jEFOoAHnSEVIaSDJwPDzoC9vaHtbq6qBDuRt+qdx/L
JwtSzdkT9Dnkqjcm/UL0zTC59mKRRJWSGF6oB4JddNMaPZs3ZqsVZ309qa/0hZNn5fhnI/WdTJAD
oCWINCwcO0Sae7UKWXKPl1oemcKgPiunoOBaZ+spAd6gMQr5mUrxNl8EnlsFVaH8rYL1cI6E/HzR
OZo7p5O3h89omvyVXuAtCtaRo4jMhALj3TQiKB+MU7vr0Pp7upFt7BwMuITW4MR20ue6j5eYxgCB
/TGZV1s5R0+zbYugAA8+iYHAMttpmWFAMbOxVS3LI+QsFDUw6gYJqSrMSwO4S4/dgzOuXJ2i8aFx
uAbGfRunOy4mYGa/NUZfBdbHG1Cli7aJfw4e0z8v05ls8N1ggaqYMgDx338fkGioxD63eK288hBy
e0p6k4uGn5iXP9vBxq+e64oUeVHghOGVpF/HxmLGLxVH+nicJgqdzG3TXhSmWRbz/HFSGlXSHVmB
+k3yiSRRY+kM+wgYcnfl52ADDArdqYRz50Jxj6MfPwz/9hYsUVtQwgkOKtMVz7g/lWIZQ+6aIx8o
OTQtdEmilvByMOsdBZIVEBCEEQkjigKKMqCF166xLLOzgsoqmjBQtDS8fbTdzwyY9sPWWqJEg7E8
gqP+1gI97wnobMFLCDy4ksrmPHF/5HwLTrtsIYDGD2PjHr8kOiG3jCww1PBkoFfCFQneuMxCSvwC
alGX6hDg9gF4mkAh/rjvTgK2EtPHj5cNpPdmwTFXvUbZgNfZY0RnJHkpHo/JbIZpc9VkC2jlCiGK
G16aSuFez0Zi8nb7jXKzRIP5nxNI3mG2zg/ApIA5Rwy2Tcche31rBdoPXSvUFG7j+zB2n+OP+zdy
S52YhJXNLmyqQTmqwFzP7q+B0Liqa47U+TaALiCVIzc5CVvGy+CtUjyIl6RswpSMZ3qeDJ6N8eU8
JAwWd9wn51I/RfJWi22zvtEDJ8vo2OcmQBHV0zkersE/RMzeVNlsy2AepBc/TlwbmjPV4m/YiUS7
I7gf+SZJU/W1TKmjechEHY6hcz7N3kjuSLPRtLlHOI20qOq/meLC+7RWHFuh6kIPs19YRWMsasOH
TXYycEYBjKULGI6M+mdcgJI8Ur/lyra+joyCrOppUaOMLNjOApHysFhfsCrMo9RJfSbUR0eJWDvN
sDw7oXc6hXy/b5kXVZcIkoISqBUk3MQdfMlc2K3fr4rL+rvBN440l5UVz9iHGirEERQKMPVtqtzf
Ht08P2nTXFIps1v83VBzVZEtYCZWpUoJBIgQPllT+Q1Jc1JylTsubI7W6Dc6XFX7wseUtZ3Wcb+Q
plRXxeYky5jjWnzUsiCW81m8xIy1Nu+eDee9oEybRFeI28ZH9QAPpBK3LQVKEXcqZJgiwh9SpIGW
R7PXbsD1zvLhbkZ8lvc6ocWo1ew4siRl29iJCWeCvfi4i51BLnbrYXquzZ5elddYatENYrBU61he
OIn1+zCeZCHJ7QI6rGRjKLFTIJPozgz4KmuXVHOQadQSuGqt/AHFeARjQ6nAQDkGvJ800EMv8EwL
F5odZVsZeKjs2JB5QMfAXe2x1/86y+a4B7y+zkGgHt5nRlgAm728RykhA7+/H8Svkmh6TrCU19ub
w2/Z735+G3la/6HOwVJc5nDXUb9vptejpoufJUTem/C9Sol09HhWjVYHKSM4wZ6Yh0eQN+YSCJ1L
lP0F/O0NmFXgcnLdw4OHBCo/oM5spuGJIaxGrfU0RO3mAxGw4GsJ1Ew05w3UE56HsLm/jplJD0p3
wqa5aumnF4hL6hsdlcvMw1/L0EZXj7USAMOTEO5+TXPlJYpF7g9wz1couZYfY9dnJ9t0GAhkUwqL
39kAr5T5afIQ/qqyfnJfdcdft/UkVpEtC9hA86WIukmAEVk9zmmS3NrMhUcq7qFaXJI13cur1SXk
E+Vw36aL2qHsoV5f5/kZLvwZSKbygyJ45X43SQUvTnUxcXGmr0JADCb1yg7j8f4Y9zswZMzfMwEb
gNH6pg+4scJwhnmCTCjpl8SBawgc0DV9qsFSG8U/+H2/z6bawr/bAg2dibzekccKXG5x5z3PUguo
kis84gxRJi6BbdQgxkHME+rV0O0zo632fS9Jy0qK6Z7N8nuNvxFAsRkIDg5OVGHT1kStwQIBiB8g
NIrFIB8oy59HbZDllwR5xbfi+MtA/xIKQvSiNrRsgBRTAOEMOcAveTufSXedYD0Aj0OGiX9e2CCK
RIfAg8sOtIh6R764UU6HAqDrwxlXVLc39X3xZ4UqrpWYeG0xcLgntK9lJ2MWu8+aIEMsDgcd9J4o
KYfnlDXNvgvBt9noDTGgW1E/0hRICh1QUujf9uYUFe0MZOYXkmQFVEa3QH+OZ4A/U9y81fGDZwOe
UPgohHOb1h2CRyOqvhTHlYIlp6VtFS6DIEOkM4VknO1bV9Ubsxfb4LGJPc9xNcEjrmJD7M2rUIbA
mCCH/bovWVg+JeDL2ogcVQZeviCs9tc13AgG+bo/OFAWgEhhSg/cotEeHSNnsI2kRLTaQbiuMhmB
V9X1UwJITbpIkpd9ipwNAVCXpXsx6WRIcE5DaZv/N2D5IWcRVytYwknddGSI18vcXm0eYcjxwFjE
8n8grTgwzsk4spmnqdiDSxGfH7Y1IIgFtBoOZBgCFWK7bWbrCV6nc23aTrrYzRTItc9D8cCWHXV0
rvy/GvgmvuV4gg9YxS2SXhEDZfddQAgFWoucT1/jdA9bwBbEgC0ApTIbdkaGBWRT1iWrV82N4iAD
2pRClgMHAXnLlpSZvzYOEZymjI3o4iA9YZGrm2o26KnVLKejDYveyEwX5bECG95Wm1UvEQ2qGuN4
K4Ejg/Oh8EcekmUt2GH086LKThW9W3CG8lQ0/EHoBpKvRGqlinklnx3wOw/Im2vmU3iN22OnBnQv
NT5AE81k9V64EjtYKgO5a+q5XgXit3FMe8s6WDTNY+pio6+A1ahPk4RN1beXrB3YfJwyCildCEK5
8am9m48YphbKWdy0AzsaX9pT4XigVany8yQJIYi2/i0iSDgg3iynvP996mwBwdjE6lXLPMUBlq6p
FnqERz4rQBnNZA1VK34jrrvckijDIAmObxqOnaTezgEsGC48cg0DINS3pJnAUdbeidXzYKwCvkBM
XBe+gJaPmSeVvqrc4CFHDKUtPNa3sJeoTmyHIU1o7C0bb2/nUw1kxPNo0anWwMWwMJ71ycz9uSpd
WUS+3P/U7vuGHpv/ZizTJZN9xzQQuzREdaWqPS11BcvR1/csQge4eJstR3eAwk/iKuApFTVQoZZf
Suswj5pVX6o8u/URGXE+1+AwquSSzWgT0KYKdR5nhX/bZj8iRkCouXB6fFM3OUjGU5p2xMqSfvAO
A3Nq5VtxhzD0hWmiyt8o5XswcIT/bGLk9nlq8VK9Wi81ew9wBXznTC/29bYqlrJzd/ud1v3tDx17
k5/BrIXBHBEtvHYeNHYRqmAc79NWPYW7ItZAGXBMAPW9FhipvN9RL6p9MNRC2polDSE6ZE5Boz5y
QI9k7dkMInHyMTp875GKLQLEQ7W4n3Xxd0vFTU7UKNRgSXeQIz6XrYRw/+c1p++6P1n2MefRYX0J
TqQUKT3sFehYSHQNenQg/pNDeO+Uj1OHK/er/oElUD1vm+J65bPIPbAamT+8V2C7veAkdWA560Ng
7lhGyJjeHLYgn6FfJ6PcB2LV9O1feoqGYjs4k+5+9pfvMWuYDkCX8X+/fyinpnkepSvThcs3gmpb
cAWU+6mTQybel6Fsm9vRpxuXcTCL91b5NQwVF75c34EdU7hAgelZNhEX4h7xgOzVCkMAnIfjq3Nz
sI8Q419H4rTjZleApvDdwkHrWfldwFs2j/vm5UJQSTB0BUZhVZ/kwMZGP1cnGK/3r+5fCb5Rw0fv
CKRgyKCrgiuwGxXuBBpzbZOgRqL+hjlmQ+67zP0FJW6Swd002ygH2HenjmExFB6+acjuVHIKCeF2
bgNJUsyf/1UnywzYyPxNnVLN1LPQ93UqInEWrI4s1AhXH69TJ8QnR3Ukr190yhv4Rubg+dUE9nTX
L1X07vmReIUCwh6f1s0C9PH/7xo3mJQNzXwyc9uveHsPty9YJYbI3mnJrFwjBl9L43cl3UYetcOW
CoCRv5oA/qgfvxvgdGxO09WSvNc7qQu6jNesPnN9Dam2WrZD+nfmKIZ9jZXhEXEJgIQjw3MVw3eJ
H2gxrflgYUZQV8yyAd46HFcaqfuyapxwVgwpzuQ9mxIuq+t3K3lJGVqceYBEZtl0k7qk2FsXDvKv
WzcyE7hbMzOZ+wGMLoLRXZenVkHEDhM24ESRMZdIUFlb+rSSLpkXhNrGZg2qJ23bUh5Wl7wHV5UH
KXiJaBo+33z00UrLcv5+F5+b5P4vzLGMhGWTxgea1O+RaHHmIXRKkpEm7WJVT5jE8hQT2c/9pQhi
5WDn1aqlzM14LzABLbo/QahQOFw9DuteYiBRSkTRUxQkVsBApXEkYQU+QrsRkcsY0lucR/U47VF0
4tTZzLSSSMBnUrQpSUzNpbdHlTXbsXsRQdXq3Jq4zVLpWkj+OxlhCKngRUlV8pvv3yt3mWpe9ECD
Q+0xmwsOQfnkeDPESGJtoBFudQEzBn9hSl65/dbCbjzpw/ENoYucc3OTCDouCt+ppJeBBROZ4ge3
PkJI9/QpTGj0CFkI6+cjNrCdjpqUR0Wfh3VmbkHx979iE35WzsGvklVzJTalOhUArQQRH0/34q5J
Ko3Xse9s0MBQnLcJJ1H2k0+JConACO9lPC6T7UjpIJCYTlAo3vVAJz4BYv3To2az05ivOxmCXgFf
9E1AN/7Klqnm2BiXVYZe7Nqg2+LXZVQB6LXqFgtgaiSQqVJ/RbuYljWQ38xKw7aUbP+BLfBCAx77
naVqhwnGElUrGLAZJ4JKhVes4ffzeEl8dFQGiO4TgNJ8mqfCXAIw6+/d9My++X6JzsJnNd+SG84s
3H+FIMKresmmlBW/VLPDHWYYnjdpoxyS1KsnPUr4KtEx2Tt2D4k7D4H5jJFq+qGSut+8j5F/FLPH
zFLQVY0k2+smaHpWwkDRFgQ3kCSRRkzQqo7GSvBtbz0anY3//XXZ8saiB/TD//Lxdp6rK53zq+HQ
Y6CtF9nl5HCWlmtD8K8/6gA0rg5Ys4OsBATu/8z4TYe3LrxmKgo6qWdQWMMWL1Z4jOM9hE1l/l2w
26G0H+KzGjo2bQbOZqf0Ia0NurXYryDPwGpa2oEXXc8Clu+DHWHu0zaOE7ZYQNEi9tKNkeS8+Tth
3x4FSb5pI5Ts2cY5erfYCSCsPiGaw7sRAREG70iSp14fRwxs8QUuiSRliPPRqlCard6NvL0Z1vjF
CJMNm5akGOpLBsm4vK0jYTOLe6TRTp/VHfHjnalcUMC2XIqGCOg9X7NPqCh4ECM/+eWzji09+eq0
Z7JxjArgSd6Q6qQEdJ48zdrJzl2uxaKJuRAwL2c48erbX4riG6G4IeXxfpks8FrB+ST+9UAk7l8t
TshbO8xJEgAwwyXuG0BchIwldkQnSJqq8DlwUPvu+7G2l/4TCXocpXZ765j4pu/vQJZiczIxwtq/
7EqSC6jumsqC46BdyRH3L5oC7GXmRpd/qMni5kNsxKfMo+i4XFMJCVBCyZxPodl84XyFQRTM6zXp
BJl/1K7QrgFHkjzNofGyhiAWtV4rop5p4Tyxvp6k4I3SDgyrROsGH2W4oVgsWLlw99Qige9LqAZG
5byGeZnPJadIkRbsDYA7sSs9kQcyQQWGjhfkk4vN5rmXjvftrPCA+cOrzVLDbDxC+9vPPvWaNBSt
SWAZWMNwyk4h5m/2z35pdVfz+fX8mdEW4r6bjrJ9wzGUe6biiJfDFqYoMI/mLnjpyJIvJfSsxCHP
DTIfdgUNxf/wXbJcE76DpZGoGN2Qr+QBqK/IiWR60JznadimlcLVUuKro83CM8vrr2bEjlb/5yaf
Y4yNsMTEOElXow9szxZjXzdw4OHullwvzcelgrwigDOqSBjIH6hsTUVWGRMFnB01wbfnWtocj3ea
NywXxgAGmYfnsbx0eeOAZVE+gDoEevMDizoUiqEYb3nZ3CV7nQthNerAoE7WtxS8ivDpOEgRdfbC
IO5E8mkZOzcy1Dj0nyLMxwi2EDjB+jZdRUk7Fm1ZdOOMLmzFV4pQcQHoz73+bHyil6t++17gSF1G
0oIZT8HOL/HVybgqsbJl9rFd1jOKja86Bra1MIjvr2YAxprgn8geQM393pkb1jrKbeHd4B+ZFifK
/flZux2Twv2qcYaL+J8FPZdj5MxhC6dXeHV4JKx2aTS9si7oqo6RJRHIxAQj9AJJMqxoieIdZQa/
5fiU1YT4VZD2PSJW8co5H+XqqAujRisLof6ypkTudyGtN9WokaTKQw8yU2izHT0/sWRCIPZY//Ma
7I/faRxQ+GznqdHu4+dXLWsYHAWT0K+CGtlAEjUmNoPgoItQmHOb2V0mBwIYQCnFDZnwzxfOi9uU
vYwfXbSDGg/XSYqwaPZzXza2HNeQho2ytmKIqjFMr9YIYrY/5Ek5v/HPRQeyJ0VOLJweuv3yQCvC
pO2fzxxIdDC4nS/NvgGZufpDaQbXPPs4eNJ0AMp5r28pxyXOxa3sDzvOWRWcBePGddZxGkGhx6sW
yEq76++2YY/4O8dT9oA8tFpeA2mLN6ndfU2ou+aW6v4baIKO6UqoRsmtcV8a/GGV28j2LdBRMTnA
4D/04NnZP5LJQaZ94EJAL3uD6tc2pmOiwUceWY9txV3rd9ASSCdsJu6GrZUfskV7AHir3h+bA8I+
LxpLT55rGU9yZcXVi2/QsoOme6tFtisNzlVBULaW7izjyj2NEW90TDDBhgCnEKNf5O8Cj1y85VCd
491iU8PJ3NZepfRv0T6Yi7C81xO90pc2wvhuNffAKftJ3fXme7+54+EGzirzxK0z3tdL4w4l99UG
/hKqGDFMv4Qy8q2FrDPHYL3Ar0UYabvAh7+KZGRtDA66opBz2CevYiYAAUOwvnM1tVpPp7x1vPDx
XPIMPexFE0NvICSM09qOBfr44VNn7du2xaXnIg83PILf5HfTuSRsQKP8eBK8M1wGF9vq1cv1zFX5
p3uzF8ScE7zyikNDYf0M28AKJ9C+WVpXgE5cBqmofzzLhXpes+OrYL0r/GXfTPOqJs+nXKMK/wR6
Ls3SyDu+1gDmOYQxRrc2zvpkYc/cYIq7PcUNPyLSwFSyCi457RaFvRSKKDGmj/BaSewpqC9B3U5Z
2bCyAn9t7uZN73BwL78fxEYIrALLR6lthzy3y4+hwtCz6jdfApNxJDmrCaxCh1UFkn4L3/YWRcJr
SZbezepA665c7RsYcIfs1AIHDsH6prYwUxX0HStj5DBAJbXHfmh0Xq9xfjuoA0B1XtFrQ3bQsDZx
DIqD2WvsiVBfI25FeoQOM19Fant7gpB8O3yn6JQdtxqw+3am+mc7/N77guAsOuo13PpNaKmi9K6k
t5xuSNjFyl9JjquOqIw2tsWNBfDYZ1T88TVREaPW6zuLr0ZioI0ozWrCwISbTm5UsCP94ZgkZjGI
an2cUkEvm4SdLOiDsFXRD1oBu3YgZ/3IbolZm0q4ZkJvQhSxU6+wg7Ax+ECexdH2aqVe9McJgj52
sMqKbqQO7Kmq8Aj/j1c/hD1WpEibPNfokuC9LLXiOFN5DcLZOgOQetaFMjiS8SSRwqdAYnNvKiqG
RvkFOzSxSC0nlVcYB0X66u9pcc/lwj/xeaG0XIlBTD/C5wni4GRox+rAWsRiSrnXILEFSOsBGRq/
ZT0ZVEqss45TMqjaNtBgTwxomV225g+irVLHijxrrwUA6s6jFiFgEBQFKAEfIV8E/TWYs2e1uGm5
dbN47fImIPTU81eCIBvfFRiJmDbSoaElL2WICdpd1RlaE0pS7t2+IjQq63hdgwRM98mWvF6mSYfM
NmawS3DODNo4qDTZrmTRGOBS52DpIeapeOu/nyaPFzOeN24vArSABV4mYk8/TDjNdyIa229puOCQ
LiJFX24yR8JhIfHE6PNDdXRTll6VLSTcOzno7d8gNEtU43yhPF3S08dGUbB0NFf1bEX+CIO61UcM
ylQ4a9548nQW/Z8CRUuMQs55C6AFvvn9U57ZskRdDtscChIVNuPal0B6mzTzTQY1TPZRArrRy0Sa
10W5r2uYoN4tY3uXbE3fM9XEQEjMRcQez4Yh89u87MVqU4ESJoRCm5btFVdSusrAOqR/0Ci9F0rQ
NEbFDb+AOhGhWdZizrXfdfagem2O3pP/PqQFUTIYZueEQrDBkmCbDgtPfn8FdKvKp9gzadblfNsj
+ZWpjGsphhzOXZelVELj/NMIPoHZcmsW1N3Qy2uC85sryDAN5xSLfoM9wvPQS926RcEH0VSS363l
G2ehrLrdUnQ2xGCdsImwIySpunvvL3Apq8ACdwzt0FRW5hYVepzFH6fVO0GQFktaz/NWdi6s1red
DIbsaW/BA41eZuQoG+ef1XM8UZ+3tGu5c7ggDqPqi2jtd6Y+xo3uXNaIaIwco47dwfhuSk79UJXJ
Hc4JDCmg/Il7g2K6TQCbyedkSDiHjDpgISewb1+fykjLP2P3k44HPIs+kkeYmXd3L6i+OQvZz0oc
BFMLcFpmf8sBfaDDYK0s7pcka9QEMBn39L9H35UNkBzH4kKNYuk1nARjUU+sEGyr8VNGeMpmMngP
MJxGq2vEcTkn9vPVJoAl8ynRr78cCOzRVZq7/0ZmIz3xYN6MSzoBP40lvv63A+oxQz96O7JnbcXL
feS33jfaRkDXi8UhM2oKq3D+Awd+X/WeVXfuuGkl45M8VEhRsC/S1z71DPkT/v+fWbSojnUm145M
Rp8fiF25+5F3DHrxWsbc411dLwmm65dOrGA28Abh2SNtzdU5IT3Q4iS3T+GdhKPGBvZwsQo8225R
0JO+XLhDfsz0W1h2as0/2hhDcKerUiEjKlQusAKbFPkSQB/daZLPN0LLETUZOBFEkyoGGsfhI6Cm
zLw17JQ8h8PZ92NvA3FX08sLq2JfjMO9bBtfg7emsVvm91HOAGshAxrWVlR5Kl891jBpcjfURB5Q
tofXLdC11pIMmFxaRauM9yOasK9NSrF1WqZSkkuMP+MWz3jQkxfXlJMuBr43fqhNjAOO0PptL/9j
46hVBt6nK+ZF4c37Pmmdb8+48prbCLBr+JhPMllHiKdY6e0+M4lyk3YPFAJ8rnWfBiZvR9VTczJW
9S1oL/izf52yNMRjv3+eL4n7LzUnmw0f6Nego+uUPcaiX3oaud9wP0PR9MMQlM8SUBE1tmwTRE5S
0UFKGLtMerKQtzfppfk9dL1Q33FNCsT1jycGmBi+FiB+xAgGszX4OqfVJJmZRa5S6Xdhy55ajcF4
t+wTbPVvYExWi/WqbeZwhl6LcGB3gQ93pLRkA1ExNT0XNy5c2VHhvKDkYPYFf9oL0pxgfepYi3z8
3G4hpT/jEPCMDwGJ7+6yC6rN0bvGKPGFUiASr7XiUqyQ1smGuWWLp7nYsTud1Lx3eMrKqzFgVC8i
7rRUhgR0cQKCDe2STNBLoUQNTfdi7vgoUU6Ufw4Xnwvh7qmGkHrHSP+g1G2hAH8HL+bodDhxnR0Y
r1sdZDsuOc5dP9Y/0FnSOnUiG/9c4FNMO5FvnWpegip0r5EIQPoX4N1dBZ/HWJ/keI/eCj6yMl6X
nZLuGes3Jmpis99PGl4e7d1OyzYqxkxGidR+v0SgIoZId1rGY8GW4XqmJBbD6P5P/X0wEkP24FmH
/hn7ys8BxoQ4bAmqQmAWHN+jwbGg93k60EflfWeOfWNqEQeS9pXU6vxaW7CIPfGNKRdwlB4s61HZ
HOBs6geXbyl0fmVYB+Ie+4ObBXFn1MJWN74twI8e7Ev/kMZnKVZGbwPjiALKzK/T+MJcmmkoelMk
NBe1QbR49Kb1ANnFoDOOu0TiNtXi9R6VmmRqDbj52rqukM++vnsz0phRMqw91ZUU/6/7GoqM4mbS
fa8i0Kcz3bpuMuNufNiNtlvIJ9kr3ar28RMR460fnMGSuKKTPohCA2AbyzodkXaLIyUldjqlp1/R
hZ90vGUQIlc+STAAwGIh3/3A1Emnm0vICtH/3JidjCt7d2BZxrLoFRsRvg/+3rpOW4Qt9eJfHnPI
iBGSbpeP3MfGXUWFIKYs/d3oCwlwUjwKko1X1wbCvhjAWkMBzPAZilSpTewgbXQ/PzOIrP9Uppbp
O94xHVD0iGPZCtriVLpwbbYpPrzqdrhu5ndiK9h2sK1kRk3KVRVWVgZI0RVTxMeCi9ehrUPUFPOJ
VGYgXzj2BAr3+tCQwvyaQMBUjjvUqyPHU+1l/JnEzhJWe69CvrPn/8xypZ+PJ7vrhtNIN2DOTI4I
BK1tjoZ/QnWVLAgWI4nRhY8R/wCstqAlB/ucJfjMteN3G1/vWTfxSC9C/EyBgVprT9ISXR4xZzvh
JkbZuGTeI7fHMwbowdlHVAuzo740wYb7aqPjrY00AFbTnRmtAHAEozNi5rpiwqCauvEIcdZqjEWv
iFqYt20OvJ0LEltKmmNj4imPYMANiOpJBKwI0ACwX6Q1XdGuqUusN5FVvnovh4RMdsO6lFMPSRBw
f58yAe6LpiFipfM7yVYMk+NeqAzJUfDsMBrlEmAtTd+fzgi16kwrrU1Z0iVVL2YgW02CclwtLcD0
4u/oRFYpzYtp6txBNZFBFUi9zKTwVJoQz+Q0ycN48JwzesLs+mwY6CEl8ptPnkYdDQInwmmwRwUQ
wy2+wH4oB5C6jxexMu8iEHcJyo3Q8+uxE6NlJ0ovFE2rx1YpmGyUa/hAhx+2V91L7mhAfRTdO2wU
o4UM0omyyWlNjo28S1ytXUxRl4704oXyB2c9uCDgVzt/6xsM6bcOiyMrj+thAMSKiXEeG2cClzli
qDhXelU178CEDkcSE3a0yybH9u6oe8QE6pk0KWVJ+JTX1K5IAydW9q2siiylpd+fpyjM45Lkqkti
obMOkGizZSjJGCVt78Ms1wHNqFhhYI02ddu4BaOq6O02bB6ogRWdfIrUevIUMsTfwDC52mFRSqP0
nJhLLr7KqGtVopmSLbS0YfZcO4BOUQojjg3ySxJRGGmCqZxfJpCVu/fG5GMqvxScNvEAquleqeTd
joPAvShNLmsEflE3S7eCN1CAByU/xj1Sa7268/4sHBRdA0FB+2zD25t6dXFie/CLdTWu3ba9Nuef
3KoPbsYPS6Tuv4Pu7de254o4xXdnX3akRe3PKkT8cG+qE3XRMzS8jMIHX98CFdsYuKOewNohY5xw
BIPUcEgxJSnZgT88aG1n5iX8YetVUmIgW7RAeiygaHEPx3ThG02pP5WanEJv3QYBm8+Ca9vlrs9G
e/7qKdm5p1El9iN5HhTnFre/1jhg65/lY+I2cLvxB4lV8MDFXfnWGHv1XCnZnC5fhwY8CW0lrzUT
QJIxtOMWmdaTgiVepD52NQO3uIDrrAHaX+EVbaYuBFuTgT7vpfynHtiYoTnB4Nnc8Yg0HNOAETVn
JN2aXbhpGemS4EO1QfTwkyJdN/6qr8Frx2NBpy5RcO/cH1VMZzWF1uMtfM6LkeyenSqwWGpTNJ8x
7njZb4iaWr4ld+rI83hAUJa2FZqKF5/YXbIy0DyufOOPQMGax25I85tyGaMViqNdQb+64lNW4Vkn
2ZpJgcBggUALBaYQueqnGie4glJIYgZWPDaxnBsDwC0m2SE0w79tWfGVBGj0qJ07hm2IFH5n4l7F
X+SrF47r42WTHmsHFiVrtDbm2RW8rq1yOwzYPYt9qyYNYiT+fFXguNNxaWPgzmy9oDy7Px8KI5rM
fNnNv6KfA3Lx6hvijeoYMeS6fz4f2RtoEkWHrJJJzzCFEy5DW7rUzDSwfoF4mcKcgKCyILnmNNyB
TV1fQ35bx+rWvlf6RMxK29hm6yg5K0MaaDk8YonY7wJ6habHGo2hoSZ8K572CJwn8/IdiY3oS6SJ
YU/Bo0up3P91k4irtDll2AiVajPnurFLP4iwd2NbWkAun/bKwvSlrtEoucQ1lVFTfU5ElWMZSnUR
F67IjmqdFtpJeGKw149TUnVV6+Jg79K/sMRcXOU665HSi4QmSCGW5wDsi1SLUSWe860HPrmajoJ2
gviEfsgxbE0/+o88xKfktWvHaOcnQax9+XTGzgc0s3TmrHascZ4esAFhNzuoR+aDpOJb2mTf1fWl
EoAQ6pr+3YZoNOY7UUJ83CpQ6TgMiTKy59nTNFiPmDKpCm/22AsYU65Kp1io5SSChE4vn1Iw3xK7
OGcjmfcvY6LxiHeNxF9j4h9+iNw8N8lzMLj2VN8izr4mi3NCKkiG3+M91ceOWPvoGF3MJ0GiX9VQ
eM/awq0LTbKsVQTMi69bLQKeGLtfkHHjDtwuvn3gB1MvXrO/CZBoS3prX0/w/YyJ8L0yZOWdKuml
P36wZrn5r2esABMARdjer+SHzobfVO5vsUBl5F/YjQNvrhX4qVNYvCOB3Z9MQbKckfiWhGdqm+sw
uoj3dtF0PqzXOShKaTeHHWtEZHy1PqodT5/DJEU1jx+Ax1oxhIIjRjCihyY/5W1FZVZI9WKkrLGW
99sxGqZ6+9U92Z7V+wjCRS8Zzq6xci9oakSZIDsDNZVBI43/SXnRkpRuSncNXMD3LPeinPeualjv
a8Q+t3GpP2muSgXaIabv97PkOE2lCgLpzAC/V+eCP1t9ytf4urjoER+nE0gEQ8RZcPUNubUcjaA2
QtsWC1zJRfziGqvjW9K1HeMqjMKbiVdn10NOZYtBihZZHSwc4ld5iRHQNzMKAdQigAhU4AmOUJsq
rg13wI8XaErSZqJM4FUl2n7ze4tgd1JZVC7zXStJI6SEoG/QS6NWtqcWPjr0BNOyYF6tKiKTbodR
P8ZpxYgFtFujtavD5StUc4RV8F9yOJVAzReVbnUHNL5Nb/g1KUW3VlmrHin3aNV8gqxUqv14l57W
ADr8M5R695nyVpio2aRg597ntIwKgEB0wWF9D08Tas17TZ4bpiem6y6DrpmzxaWqxtuDfsCGzcW3
k7zhUOYAfVQCnU1ufgXb2BeOfETTQUUVTjADUC6K5/b8ifN+2dSv329HHy6OKBHzdsnx2Ek0Olxt
HRJGMEt0j2SpJVh3iOR+ssPA6VCEYcL1WloEODQ3lHgL+/Q4xmAa1eWc80fPtaQfPYvI7Qr0G/zr
7gABxZaOq/HuPh4cs6n+O5A3oRgvHyUk0vFHzOTn6m6yttgEGVqwqaoOK4bd3RKyPfCK7z6kQ5Rm
88qi7z23UUIlfW4G/+HP9KUIfeMFvDoFQLaZoK7XJysqaivqM0pwJ5F/g5i9tVtZFKnkf3Mt+BDQ
Xm5iBWlhBFb33uRCFH4JcitsxZI0eEJt/JHRna84f6Nj/0cI64ZwXzqZiDo0BCC7JBd0ZEdZx9Ln
I7+Xbxua5yTebLlMklUCy/uI6s6jyplPQOqYd5ioU9OzxvsTU4VKBmdomh82hPXsjfUEqF1JpF7V
0dwBpYh8wStVGFS0x+nnL7B8aEKMthx6yrmAlUy5w8IE/Wl6Sf4F2G6chBr1INZpk4tLwCD9SvnU
vXEmHwLmZ2ELQCd+c0JeW+weVdlwX71lRtSg/iXbn+9Pv97eF2IKP080JH+hpCieofLvNbT2GstR
VRW0L8rwIXp/OOPkemD1LI6YA8Ck9NEryo2HPEopKdg6GVyTVRxLdQUoU1Ui1fvF31a0wVfCRE7R
0I6BMwJCy+QTIRqGOrzGsNv3pRmxpTcCFuD6qtZHiAKY0w+ezOyp6hI6aSLVwuJKSSCSPTD8aFtN
+aipFeJFMdZyRRVPKDv3R1Qp2Snd0eL42ajR7FX2ZSTuwmgKRhn68u6wU/sQfZBEck0x26bowf9s
KtifplWJgFAYDh9cnOMHHSujjBNN7IIy0AYfex92Woc8hlpyRBmhw46oeuvY2h4UxkZDz14rl+X5
+3mblw9bwPssej0nqwG0ijchsh56QcLmDAVgVLeOxFrkJOwdlTj+nO9utBg3r6lfuRqO509lzXVd
WutuvwzFXVaxQ97qc5XII0XqKs6scTR80ECaIqgnLVJTJq6uIc4A5rVQyiyRvMqoGOiEkIODWZW1
nmYaJDObTe9SlCfsrxXde5fkYxPJnPsGvNsqAfgjsIAmjU5bMds7mMhl75CrvjIa6kRphQInIc01
MOC9XbSB5TccDdkRlVgGA+vqN1ksfpUov2p2Ao3LAQxvn1chbChN0I9mN4cPn9PDg+nXcj/4BsLN
pUxsLbBQcMSzF/uws9Esh/jaY2Wsc0rPvmtKwGMZcU5UH5Hjm7GBqL17F6CPlK07zOrwr6ajz0GU
5Tf3UJFuKQgFJ9P6pLOTmEYZ5wNA3I9Je7LghofHBZLVVjvbWesNV7rHnNwg+dkuTLn0OhFcmuCT
5bQ4iaJWFYiDW9JOcZa3HowcaiNM3+npKHorCR3UrvHXxF+IUV1bf7h/vcghPUXK+BI3KC46AHaN
e9x+QFPb9bTuMyUze1KVEnDfd4jtcIESgp0UWi4HcB/nDvVD0nWtr9bqvoGQVmUXoq0I7WB8lwFq
cDVLRHZx6kLg8+lYXZnwLh7UPb/og3O6S+Tmi+d6Mp1rEEjzzftjxbfbtlVEVH1bECFPtAg2mjBc
HT0Rikmipw+Pt+xLUeadx2IKI0PHQ5L5Y/zDVgMif+O2ssGRkhNDlyZMTHnw5xsfLlWDOb0rteN9
IBa5FysjO6ItCPkLfwqAoVMf2WsL475fgKGTebi/0VNMY0ATzpWKYRKezCknIYE8y5pv98swfmCV
a6v7voqmKWUZ7JN8j9igsFqVkw35PUM5uTGpsCYt9c4W8Ec5pT2yvlfKjkA4IiOsfTyD5/Lesd2q
uRYtNsIaZ5fhbY2opgYmpjuv3bMYjvmztRi47l5cT07p2rUCHWVd9y6Msr+8oGteBGn786RiYCzN
JCXHeyR5/yvJhe/SnF5C0PKk2dvzBiG44YWDh2V0iFjMglvHbuMzCmjh9JuTElvu+n0ZSaw5aLZq
eVIkst8I2etdtCG+2xw1yci2NaoLmCKVVfawf52dj3fbe+wFYuW/phl2IDIIglh2fA37wfRnaflo
+lUvihAo1EojkCvHQxbLBuqWVaQYduh/G0KvJtLrsWQTt1vG0AxzJS15/XM8cKFTanOtihyjb8rA
Bqp/0JEGyPabs7jKKa4snzlYoAYW8ygu4VeE5Fk8g6pMigLLqP9UlLKUQzPVhptRvADwuZ1P+/4j
qletbuE2yeEGpTUyJ2S+yx/IlwqarYd/8LEgmnjNVJjaXlRvheGuW/kNyZtkYlUKyMX6Il6DCm28
VfHtu3rBj7YlLF8/oaw/895LeLwyLV20n91snbr4kqlFRZKi0PmUwwtIOHlL0La+z96C6S/yPxel
FfjQ6JSOpRuvChliJs+p/yBrdFThMCDhcDY7UfDxRm+iDbpu0XHxonZjuzQOkUGoGGt8/MOu9cqq
VGx2534e/j5fQNkb512Jwc9ZP56ZKnY7Wi+Yo+gDb2ipqVF0MuKYqOUOsxQkMFNHImcWBYphudo5
oH+CziQ/nE42w+4sJ6mSbRfhl7t86hk1z8VhjOWMIG8I05EoPZ28xw/XbGOMf5eGoJb+Hxt50OOw
nKXlf3OEteRfqZoTz6ahQZltAG+jGh5OG5KcT0AT5a0/G10vHXPOa06g6HjczvbVxo6/tVPBx42V
oGnTpBb+ub0UmE4sd2dn3H1ZlT7eZR6sLO2+8u5KIFaaTyEiLKnXj8Wz13TSkcqXz9bdXkY90oGW
VMcYOizkXUWLUWaWfGiXPKR7iPcHf+x98p3Zj53TLI4ymy3dnEcVRsE65+23is736dHlDYWqnC6+
/xpvIXNkzZmtzlfJe3/0wgC675bYKnZopF0/nz+MPGQowyAM++D/qPaRu00G+JFQLkzOrdsv7T1T
W3V02I0JOOlc/FW955OWEBdqR8ZeLSQOyNnAMMzxiS1FV2v5Fg0fosLxl/NNPM+6vbkypzniq2zE
iWr7pD2497e7zwE3T9qEZKXyVvqDrjFVk7ANx69zN/afuJ+TLWWhEml5kFj8ZtYk5W+5hNFUVm/K
Py7SS7V1jfR73WEeotGtTCBvRj/HYo87c6YzmneH/xjQjx/2kesNu0oQ+yZgwzCCo50dfm4KqaHW
DMALFBn0viZffJC6xfChQrfdWPcQjOokzdQiWmuOwk24VLv7tOHKkzNlTI/PFnrGrJiK/b7ZekWt
pQ1kxF+5FUSTK/dPKS760UzJw829HSG4v7XCoMaNWG2ayez+XJdhKi/o4OFynsDUdVnCSrLobaGU
5dOtNWMxQUeVN2JnHtuuuTqSL8V56UmDH2TSCWzbaM0AIjc9CGor1VTNbdmSEufYviSvGs2AoIlv
a8JeokCskhgu7+9ArL/xOO8hkmSqOZDsLhKUBGHkuMqDSOG2lffqHMUofnS1O6aPXNTE5mGngLk3
rp6u+j12lY7PfcHFfUTuCca1Voq1OhhUCgrVnlDz6TUV8F2jP17QBtlQIqnrelZ9xUsBb1eG0ZQp
go2zU46p8V3SVnD4PCtQrtYTlBgCqGt+JZ0n8XXynvdRyDPJ/yTg9lF36Qbl46KrWiYW63M3+YcQ
OWBh/BqUeJh4AoV+TkL76kd9Su2jg3IRPQp25zeeRAiKDsYC4ZNWENnBK6cqm6QZXHBQs1Uzuvhw
0XXV9fn4Vu7HgY1uRTpV3GVYFJPT7NMzmL23yxQePyqqh6A2l4UN9aDp8EziwJUAoQiG6LalgQE4
xL5Ijen3idbSEC3vEhcbAUXEO29tky4+6oH29IIfGLKDEc5f4Elyq1xGa6YUFyjaYoDZl+nhLPRB
WNUNnr/SjkeBZ9LWsd/p9VuPN695QTsEGDiypOQF33lWvBKotRMMD8dig81ujX/7e2pCOM/s5K5K
X8wZ2H/VQ7DGsoBo130fEgGiJRG5R3jqloTDGzEOhMqKnPxqxBd/YJhAY282/RHGGo54YlHSc8Lb
kuLpNyn6wV2tKjB3Zra7BVasIcle6HhPn8fByqMfNE4ob42z+NELN/Q6oxMopmBr2a5bzbiZdYOp
hjc3WP/5+BbJPu5K+guGpDzIC2C5GLggD7PSeHGwZGEtqvJ7kzCI+mXcEtsiELfLS25zPWRw/8wS
39ZiYsgRNSZw5gGeocfb5qW00yL8J50/Hl+JDl4gFnmzdyHqJC/nJwULC6nZJlvXYcWatWH5X+tJ
0YsxJi2d9wlAvb3muY4UTpuz0dP7C3gXTY+WRgAaZAEHlvBPLe5Zh17xvVuwD0/25cjzzzUcEYIZ
nAjllzyGVEPobBaR/rXGuTgsy5BuQtpdlHVOkiFBTJOsiBAJ0p2C+yxz0GYLefsD60lzR10vBfD1
L8egG/d2AZs6NaoDgr/QzOXlA3ophZFWc3aqhsik7UbB3sMU2zQFZevotG7GO6p6MSpFP+WDHR0D
R3rJyO8jRn2vZDxSjmeLYEiJy/yeTR6JOHLNP19KeZkXPQZo8rQQZstiwErRvv6pYVZAQpTskyFF
/qhnVnlo876wcazv7q9F74BskkL3WhbDKmBxK9FUuGjOyRyjD6eBjFB7ctcJMJsgYfl/1+kLnZZO
dxxoyFMyKb4y82qcf2yP0ATataiokmBCrt48W/F0oNsMOQniBR4GCb+GGSTzPRyJvVlMzEKbD9TU
8UDcbthLu+q1yqd20Q8RrYNVflzWoKbaEPugMYkfIzP6QOZ8U1U5DH33xrWsN7S6TXeQ/CApWm2H
G0804pFzztm+3LC5NSAWCmoLbI+nUq3hYuQWvXKeDvXjOdc9uyjjF1fcBAynLNKjffvJ+MCXZbEn
BUcn3mlgrb6xiosNWgXtu13ZQMlbcuP2EK9YlLLa/OABF+rxEUHGscM/MvBoPh+giv0W+eHx1qXI
jFX8LExxmxybg+VjHuPuZRlyPT2i2pywfmu2fNmoGTuKy/vKvrzDyZToy94SbVVQrhNEjClr4sJ3
N9ix0c2ivykI3ElZruvqWeIFr3d612qdYVtSakhGHvcA8QpyVeeUun1yjMlDzuM7fH0Kjj7H1eFJ
fbFJisOeiqcB3bzTU+ParpfFdlC2Uvmp+WpaUMRykeyFfiacavmLD7pzdMcoX5cSutmp25ARwK3V
51eCzgHT9fIgnyAtUlqo40FLlrMG1MozDMSdRVdkZJ/Tfd1XA8tY5v++g4Uunh4sxRGRf2MOqvgd
7G+UlJznsowIjQdCshKSPml/5TwcRHOZ1yb5OzRihY5wqcmw5PPjor66W+klBKJRGfdObDyiflS1
Hi1H+Ja+lHFwZqmzn7r5m6nuZxL3kzmcPRwC9oWU3MxkrPUzMVBlsLgNJVVOP2+p8mX/eQPBj7MB
2xeRdPI3geAp4nIstJQ56LbvdbHlvnbmK0QOdAdJ1/de4InEWl9KOZELDZ7zJSEIk3MS/A9JHchC
Hn6FVyHxbSENyhXaF8XdE5zK3pVFc4bCTdjOQwePI65bZRABShLoj6KKI7SjrZgBekjUiHYjRw4a
06rUroWVsaqmZUoBAPB53skzVavmtB/eLsQzzxKKAvg+NH/j+qL0zh9PaFgVderCHAbXuqVRlsfg
ehkIIKFzrvU5VrA/4CGTGjuJvFwSbbzbKiNJ0SHu2xsKXrxFF/SqcLqSwKwOM7xFr53s7HCQxANb
DSCnCLYrd/NXTsS0RqdzvQzvBJAVWd7lr/xaIjLDq0jwJD+KQnZTDo4vTvhlBB1O6qfDyI/89Zga
ZAqzxjwoPwP40Hs3v34UBVu9iEMS3nTelNmcKqYDAUqH03cs3HOQDaiuydagxL3bizyo4/s2X8tF
+XfKZnu7SFhA1y2CGC1qmGuzsL2A0Fz+HqqdOY6dmz1STsx4as7PvFGWtYWwELM4S6pVlbEhx4IQ
TFS75VWQkXnBlgW9LgRFwbcU4iOgsPqf+WMiCvsM60DDfZzReXoX7KUOoExSydEpOLUffYB/KubQ
+QzlSUx/didGAvvAtIuA0oId08HZQy/ktJ7FwVUks0u7i4SIy1z4XolzzgzcfUXLo9BYIciyzLry
GrcPnNW+VIkFp6Utr6SAwu5gN+zh/v2TwN9cma1D3WKDkop7peWhSA9vGE/vg3EpkOBn86weeRmp
mXIGU7pjtWuqaGpqV5QLlVmezGpyJN9ZIFzNlxEUg9HvxysJ3yU40eo4AhgeMtilUco25RzW00tR
COg49TNSHkRTBvWZW96ENi3//HEG3QfR5IgPQTXKBx+kgnPEjdPl3lTelqBLbsEvOtxxJJ7ygzBh
R/ItvcyqpIDEx+c26YUci+WL/k6/U2zL32tmC2MmPqwkBJB82WfjX+M+0OF4G0D5E7fZ4SW1Zg5v
7leCzSukZGWb8wLl3G7G9L2eQhZYDn1JbdRWJd/VVC7+9nm4D7uOuCKca5vkXigafoEeWxtqlOCV
1IXyaGYoPu+acUw8eRX///TQCKnXhyEalJh9/iMARYFFc+e1VPWOBHAJfzBqQ5BTm1BETQ2WPnN6
wZKeuNASM9Py0mgTbR9DjNroepyHgGHgetJcLmbvRnZ1WRinNZkmD8VlDfSMt750urSsAie2uSsm
94lguGwTq5pgqElGlij8rKz/iSX7qtWZpE4KSw5BJTaktWM+Z3QgxsaO86s7h8CKntvRZBD4YUKa
AcNchAQ2qdLsLYo7dzr4y5unukBhtCj6lpq7HMdx4BdSewk+7KFa/j0jKtU6ZOPhSY47IEo96TIv
3wI1/0I7Ug8yc2ea+3j2nvlmPTzEuRBjLOM+aSU7GGIF1ncR6d+0oGIkBq0NE3UcYPVT+dFwHGku
ncy+wLzsyHTdBq/dFp+KsXMkrmPEPRD4vGK0uewrvcMLKQDTtZfH3+DYWlEfupdAaHcU1C5q7Kd2
iGvhfvmH1lJjcXuJ56DlQLmZjcVFGMhuLdMawlowA9lzyEwCUaNT7mHTlHR/0M/2srojXet007iW
Uk4061+2VWdjcSBCjXTbcl3u9dH+EdNk6DMR5JWbLX9PZo5q0EcL1ongDxSqhx978APzZFXYjZUa
1Mi2iPar2iKjFTV39jSCVKB0PuEFkp57LmUoGiEz2V2GJ6k6ztrG716L28KHuOCvKXL58wBmWY8D
OfwYJRg4poaXMVMPOcfzI1zEi7AUANfwdxA3b4ybmbfGNQKQ2hQm4lfvmx1B01FO6D0Ft9Al5uT8
NmuV3GzwEpSkVTxJeoHo/mxeXyc4L69sLcX3wWf9x9bqVadulPqUTz+zFmSFKTfIhcqLrqsEipM6
9GmKW/EtVWGbxhv+edWh7RgPeUus4u4AJhyitXFQGBK2mLtnFLqL+mTf+fRB45EQf9JwHFsNda5K
aKRS5IZOia5h/ZQE556E2zxbZMiI7XAVjcZF4qlnxyesmni9tbryiYlvUWQ23hp82MgxX9CDtBuQ
+FJ0C98pp+BlO7DqIYA+XrsBztHd8IDNiY1nHX7426nE7kfNx+8SB3mYU3VS3zdy1iOC7EM0hvKC
TqRVgkqW7csPwAWUfPb47uwM3P77gYykP4kiDnBOIzzXxrwWrOr0GM9t0vQ7T4mT2j1cw1KAMj99
v6EGi570I6ypbX3RAEhDFqTPrKNWpDjTgNnge143mBoOz9TZwUhmLf355xl+23/1vRyXrOpryCyj
wNzcG9lQoukK+qgRJdYJKdTNhvk4leLfX5b/JY6nWETtj4NlY4gR3MOsbdjP6/FQZus1EglM3Dem
kzuImHKjlsscG8BoxryNoekEq/x6tMN+gsYhD/BmlgtIhIIsV7Zzwt3Mknqgx3TAAszt5rNzYBfF
udlbgQ+RdYAfG+LDa0pzhPcYz6BbNkI4EfWuNj2iCa8y1RPi9cWwpXYazpF6rJnz2LecGH9Mjkuh
nHedBk+RWrSs45ZnkNWfOJiTCvyPtg10rEufK8miRsxhdLm8MVO3Z5yilMM+DIOg1nIAe/5Q/bvw
EP3CtW/QONlq9t1LTlaO44dk0+H/rOWJQPGU4J33JPSnNy9geKuDYCPtGu+aJnkNJ3uyi036dTvT
uB2LY8xXdJwnOWBtQq5OzZxiGRI9etSoHGjE51zIJWPTxdc+SVLI0Q9Fj6fRKbZV/BJNnIYvSgdO
PLfATD+0zSA9iGTnRst4kFYr+JED0n0mbQo6e6sWG1BXGqR47C3+KzlhxE0MyVD9MDByVs3m6WZb
Ik+htBBU+0TKcMMr+VISp5W0FdOGsK9+eeisdlqbKhiV9z/DjnObmPgmRMSAvHu0fBkB+rpuc0Hr
Hz3cbFwVo5gJdMu+xVbPeuQqRAlxvLisFTZcVXjiFd9euTs9VjoAlfaup8Grh2hWCkbJzXWE4l+6
y+UbX+LPRypSx4yXTLejAhtMzXpQ+w06QnbbsqRaKggE+KS6ImrJkYwVKUKDX+LoyN25w3Fu5Jvj
lUEAbMlJdJ821XPcI2wer96qPFpCqjClYd2jgawWwA0UCvfK9gcva4JeYrDl+s8MZL4OZmIsX686
s+CV5uRUJTAbpDhC+V8dMJWsIC/v2fSnJRCrCoAANQ21opF+qOWUyicHBgBbOVeyRUUxhIFOq+MU
L3pJaxQ2kOatZTQcDrFk9birmvFfon82TlZn6QpITbae+uRCXiEmoprWZWdZsh2EQg7iHuq7bk76
51cSq7IkhvYqNgTCYjCvN7bGXgZvX5OCdBaUnQ9EXvW+fO0L+zPka7XFWBKUO607WT1oTHYjrLqN
fNUx/GXsSp5Z6bAwQbIIloiNWk3SGiPNcCYn2jXx+f55jbZTUZO7slzzRw1IFn1ow24pudcqlVjv
rX/Ahl9H/0XPUGHShD8mH4PRB//CVGX6pLSU7Lv6d3CEtlVLU1RuL9f6e446feDZQjVVvY9deu49
qBJ0AoRlw1Pn+3Gvmhu/CGZoouFv30bqdeRgDvjeYuO0jJ7PWubx71h3niC56+k3EKfh1ZjM5ySD
bZw32Ej+SPObKVBKvm//+Pc51ImOX+7b1mjhhvuOzqm6W0dAVYDe/3oDltOOVA25uIS4R4AlNBi3
3I5UhgmU3CR52NHADWLrC8jbvsdw0ybXun7iVX9WSIEeAF5c3Jfe30aPfLu5Ekl2UojrIg0gnGD+
gNDFfEwsULs6sitt4aSO9acn8eJeJbqxNs9xzvkbwd2VXG8YnavI9S4vDmxr15DJ71p3ltuh85Wn
gsvkHEBPs7q2Ho9MKVX1bofsEvClcTPS7F2QiUVayReku0PoLxjOl+g+WbSctMvZMkOXyoCxUF/3
9V6ubOR4iKG3B+DEUZzNEofau3Qj6lTTgg78FLPvR9JHXVq9zWVAdqDHPdR+hpUhcDyuAGKuWjUP
VzBe23hyrNjyPfFMupEn/tOLHUjHLZMClutXMqEhaI/6ZGcS6wY6Qe7v7UOzQukGWuAG54E2I9Yd
YONaDuv6KuUovce+Pwe3kWbD34PBKBAEFtvZHlUDsoTtJCNAbQiF5uE120+J1pSRpP9Pwi+Rs0kg
F9p1ujSXHzpr5KFmnbcI3f9n4LPbUhU4cAfXpfxkQxT7nSZ9S8zf9QSEfnfMrD3qzX3Sd+/+wE/7
u9mfLQdRnpiRfOWj6SpnLJrTcTBW+rdtL24qi/v2oUjGx008kZzR6+XvkJChUdgODlFCCOiTGrnT
KBFzuTIhyiLQT8FTI7wK9J8nXt2xdE7tCRwNRvzDQPDn5CSPzBZ7LdnxOEfBx4eBKwxui7CQf/tV
EgGjZcNwziOjiFxi/yU/6ZK8Pt+X5QKYVwoX8tpQLBAIGFFbQILFs8/F4MEnzVKXCDDlyXOQZPuF
+pGcmZKFtSWU5p8Ydx/Hep6tuvPU99luxTFNArHnVvGc7QzFUT+bS4VYG2tjeQBolAkB8jqRy1DX
3VxPLbNxJ8fVyYQ8+W8s969T6+ys5y4O1V5aXUuHsgbo1eibUlBOOikYt3Ees9UQb50Pm688r63T
DFJIc4qvbP2e0XIr5mzYOStXwzAwgVU83Q08GiMf5HzxWc8lXDYUSLZvxJRg2y5wu/Sw4ybFZmpJ
fDfXQ7J7WBgsQMo4mEG4O2/oRU2buSHNH3gRAj835/xFN5XoNqGtvppYSDfz0e9Wr2ThREb8MtkH
2rgyDmMqlJ4SW6WN7KznHGJ7PboZLOsWQLxkdPdr6XuvrmEbtkkP1VVuzEsceS+FHqV8yD2WDIas
DlPjeuVf6C0SKNjIuEyY6TO7U5u4aHa/9rzAlGmAaQGu2/U5KWUDqcVgq9pYgrXqE+IsI3xdBJWe
yzRYcYJGmQd+k5V/ggUfCYlmF7gis2X1PMvTzfgMJaPu1QdiWMsmSUv9buDtaD8uUshIl8+h+vOS
N+K9dlhurgzpZ4hLhSMa0NFN/y+7/51Vl0t7abvkL8q3x9lqOUv8bwH20TFrMwAqtW3hzsHm/E08
bqjXgjAEwvGEuoNKx6l/sHYgfYX0uyBvGtfVpT4WDTO1/Qmvgd3R3SpIILYRpHUiPOXJHsdngONW
3aNjhoBbRy0BQEWCr2SF1a/Jr8vYnYC+91Kj4AuoGmOZz/pj6LCCjVDN1/BuyLUAapJcfTb7Y5zb
d27Pd4ZlaZq1QpsXAWRU1REPkpKjIPaM0EJDUbq3bOC6bTVWyOkAXb+tUB80Qixz7NT5wi3iVvNJ
G9uC9BfZNotqiiPKc3GWpkzubbjGBW1DF+GXSG9pJoMHTFHO4kQBJG23uvNGKUGMuvnUOayyYIQX
roqOWT1Fua1oFsjO64tDn1vLydbTOHMG3OHjqFgTZSPBtkScrw5Fnim/6k9Rr2gCIZalwDlq2MQv
JsTQRT2gA2yj+qvxMU7+X0PJ/OnAk/BEHU6qJmXuk11tRnUcPKyr2fr/XI8wYUCs85IbqCzkTdN6
gPHB3UjFju6xwoQGGekvd0KSWOhRVdVl0MP+133oMJQhcK7nYzpp8u6+D9Vf25MFU2KoKZ4D5Mfg
P135VWxqrjyv8eJVvbQua/BX2VoaAPDBcQKHHFlDXeYOnjT1P/j/taIGNaP3mU/N6t+MPyhDrbil
2kH9eaLW8Fz1082+5tf5aBQaE5umwcTufxha0lGSUGyTAjynCbMFLncxMiMf8ggNlgP26ivy/14b
aas7VrvSnOVsTSuWpzpLkATOny9iP8eMNvVLuv0li3TOEegsz5fQSQp2dD59Jsx04cJPcyQLjXQZ
lTkglEHVInPv9xKxFMwbXWPjAVoSkee320KHGfjrvorJR+6qLy1PeycciwoBWFkR6MmaYw8kyOAU
pvISwk1tsQUmF7hdaJiQA3F0RiArDSDaDADJ2+D4shOkwzJRuDjlb9uZSf3TUAsDQBLRLlEGLFtX
yfP0EvRdZ9gRgzIxVOQHiTgj20Qihlq7Z/z2dogf97xIPoJzm5WY9kG384mdq6Tp/MMC1H1k00z+
OV9/neHzLoTfQvXqR7g1JBNvymJXM4n2W4NVpwR19bLO389QGHuY6X05HkTWxuOdYbstUcCOo/z3
cz2FzCqWHjcxpDewn3bTKr2Hcq6ZaaGHUSEUvbgjda9kjyVxETI1VueTiMo6kBe5USgS6Jj/mhMw
BOoc57OFFgAP4tbary6BfBs992YuD0D7lYaAdYxvR8mHkb3yf0TpeIfjEqzDgXRhFwcJoUVr0PwT
+3FjPKQjcm3zrBw+e4xatYaQyB2SU6f2I6mQeTlpgMjwa/+IW1755nK8ME/LJkbEqlDT5GGKQF8M
uu8coygQeh8CLwGOMKlF/WU5GOfv8R9k4d/Gn9FzGfVveCZzY1quAWq9f18k1v/3NuFBlnKwVVmX
gSrPk6LoqLpB5PwG9gsU+l+rUi9QViU15mFu75oiLi5FKMjP0JfRghK7qN2eZxBbtNm4/ZsdJ1/A
WEgGAXKW5L3UsV9LykffJ95hSDEpYZiUsCwUfCTDA0XNnTkD4cloJLVEcnpSGMtwNetuDinh/WTO
c0OwQcDZRGfOoubU6Kkx2Cv0h5vN2Kv4FGTew0Jkmmi6NQFbla1Gcc9wnW5PzPj7y3OkhWgjs+xd
KbOKouNHbPOSbu9PMYeRgz+kYVJqeTiRmPJOtPuqlxcyap7BpyELiLsjGrmmrWmykbC5WC60+OLa
1XsDpByLLeCTqihmJVqyYoviCeslbazCBEaKxrKT9DWiDd2kOOe/WapaSZ40WoXwaYzXHVe0uYVd
VBeoQ8eNAEMtAeWgpKnqDHA32mv5hoxvjkKtTZW3ZDPxNVRTiP91gw6wroPl68k0TMeVDi6wUCe4
efuS5DzjUB+XjVN2HN3sWUoZOL//cpl8QVBLeSgpwQLIipowCee2LY4GgIpY38pxTeR+67l4DaIM
jF3nDLVc3OVN/aMbJv4waaXzkTK0ANK3HBMvT+83lBajKuhbCnW3qk3f1wExJzCU9zp+mRDNoESx
k6I4BPzcOLktAqulyN2EgINjPz7N8ol1shW+35fNlGc3l/QvRTBrdvmtROg7B8vB6lNfir0FNF8m
xu2LdBjTHezQDJaPM8gVnq213rFnMUjSZs53lnfqY3ZJiklQSTjP++fMgwCaQFyKWR6NdoCOVOOV
tTSaEeGgwo1HAgKqc5EEWl+1xCRHKtai/baY0s9nmJ6x/Edp9hwLfOyDciEvchMDzfI4K5ngakgJ
2EUluK3RmPQUc3akU2i/2ki51ZkwrdlZuC91rrLEAz90kN4zgsdryUgUgAl5MeZIDtc1ocfbnV2k
uyyB9d/vmdjdvYajYKKBa0nX7k68Umn5aMHjbfmObOYxhRTRmVy/Br8fFZKHJQQ1sqs0t79dCzql
hjnQ2D7qvCCcJ4iC4GbttJMhagVFEUfHtuptfBDCZyXJNLCba2E/ojxdL6YPLZzwlF9Udv+lIIu3
eAU3eQ2XNMi2zNcb4TeaqLgBMC9eQHit6R46ncNXEmHnh9UkGlHz9SrkTKWqFv6CC+2OLJ5w6fNS
4IdXvVasH2caGG+mW7Q6a73HicJImVcXkzqRpMWY2/Ataf8xdcXDkXWPzkbEU7vtTvrQSURmmDbT
cnAwNJH3Q97ZxEuUX+6WzvOwcHGhmiXWJZOE53512dnZvD91GTKV70xuyeyYPt0h86Wzv7RYe95w
NFJqFDYt7FcbaNmC+NUr8sh0aCBN7hoUPr2L+q5kcGDHQPopHm9M8KgsvOUnyPrdBMEf3geC46iP
pgjisTOcJLXp9TelQ3wygKcRWNye/iNoUhLKVrNmaB0zsg0dVKqv+hi6GvCoVyus5LxqgP+9E1xY
toM/Lgz28CU9nY0e4qv9xJhjco2VxSJCM5+5TZ8pgYYaxrc4/qwFgu55dDfUSmzUcFFnIzaJz7dg
50bC0Nw1CCRGf0J/6Ivry7WUAqazBMWGVYGSjigxZJ22Za5j2r1DF/DQZWrcA5xX3DGs+GXWm6B5
6FkkXawJvRBHUu1fnKJMcxCsG1F0QnVlWVME4Ojf57ZGrfeQGO/glBbF7m4R1YDbNxf4Es7f1987
pLvR29qJ0TT2bSR+RuHMpNyo9yWUCI5yeANOH1T2g0YFKnTv0qxLVslLlwe42Dj3GbCUsefVTSt9
9+OSiS+cym9kFOamhtaW1L8Vpork7X100+H7vswD/EeLZ7bIIRNc70gzL/zsRRSlcKqGcYul1vd/
XejD3ng8+MgxtvJp92CeIt925bzhC8IMifVcAg131Jdf6FlBZjYARugKRs8W4KVAt4k+gZqRnCDJ
YtAAbl3euCb7bRtFT2HDFzNzfz60IGOOLPIimVjPnFOCHmH6s8mTHE94TquHONtnOr3ggQNLWU9D
YyMkfdwwH9lD4wxcCQG6Add6OtRpyAeympvI2PUkx2UAWLR4FjANPBNwuMhtYn1wxpf/+GkrVIOI
lXwCP6WDb8XNWRSredJgKw8ws/WwwwSHYVhaQn/gB975q9jq8nnLxiSbVPlshgsRcF6WTzMAICHW
qFeKKvvBeFaht4N/uSD8ZkLP0tjqd/WsZhm/wcn4mWPlwP/RJfaCMC203Z4O1wsKKr7gSHkzjpDw
YdAheF7KXNCybIz9wDOKrCHbb5xnIUGLvEPZRSWoGrpSde0Ojw2X3u6w/NDSs64irwkUtN6I+qKU
QG5psDvoes/WL2bHbY/6sqtrhcqvM5WBzPQGB/ksWRpea0dTLy6mOdmSoA7E960IZhyUqcIJ4wy6
E60euNEe/+jRSk9T79rzJYxOptbk9NQM62XlUXQgC5jQv+7CqgtYgib1eoToEOWaWVzkQpzKFz3H
QTOIJVwjephAReuNgzYc1ViIOx+LntXTcRrX0oDW2eavarb/Mb1Uf6cEfvrUaVBLTNtNlJL1viLH
2lTBjeli04XkQw8NnKU10tZid3h14rSG9iIX2xNySh820arigrmsl0/bxBvZdkiUQH0+Mq5e1Sf+
NLmnu/kWXpTCqPbIrw128ZqqDr1WUBFkVec2TSZ2/4hyRT6lxZn/iyh/q8fN8xU8FUkqTnh3mxE+
JpCvL2YtxJBvvHfOX4sBDVFSPpVkEt5Ir0yDT9aZ0jvdXuhUN0JUd1QUtOCFFHtbkqVuaByKU8wi
B0B/s5WOH4SOcGcIw0+Td/H3ZAovpGD9VBs4DbfyOMM+2UhdXDeeGgRjKCd0YXIPBBZBAsnduiEa
decdXctIV+NkrfAvcKe7wzGVVuIfQrNJPkhSw48rWgwQTyuAE6z3iuIshZWSmBoHX3fthDqysobp
DehFbX3XOl9h5BB5S+vmCf28H4aM4BC8WOs4g4wxlFzBwG5TBdhDFnL7WiUKzjn0XfJtgQEEsTOH
bl80cwXderMiB5/Y5CAHgXZjlHpu/iX0UeK+G+GKZHOTlx6WhxNgzwQF+1JZEAbT9vQtB3WNZtIc
WhcZh9LrV44lVhoKts74uoGoWx9ox1Vzt0JrNaUkNHNE1O0NzLGwnP/4Vanm0T/XahPeUQ1RG62u
xkHByrZAgBfPgzW3Fdgb//brSTzRC8ff3ac2x4z9E9DqZA1yC98IJmEPyRb4qGYhA9oVTOVA+yTB
HVHthfXnpjPbyTYBKPTyUWs2Y3BBXgjR+FwP/3kofrWBs+AsM/W4JkQG7V/QghSF7G5D4LSEopY+
/wpwtzkvcwAJ16M1c5VLCOOfeVUQvsv4bJRgukvJSkSIIBKIVgMkd6Lr+tPNrB5avk4bV1/mhV7J
zIktvBCJc5cNw25vygvCZyXShCZWBCkzvKM8jc81lEw9ITxpaDGvCZcjCW0khKSfMFwUqtAjPxjD
/IzcyJUSjTfXmjJgZ6ToNZ3UyJJk+6by9Xhtj32Ei9EQufNE7M3c8R3vaYmI7dFlajkrtMykm/Ts
RuAol5Iqa/TW/nFKu6LRLBzvjgawo1tZ48fhAIqg+eXeL8tOJQGjMA4swjZQYYDxDHKBI9TNkVwE
ZUI+6i370GqHQNtsMx893qSKp79PkIsyON3HPtpMI7j92mDJAB9A60Vi7mrpRHwVkC6JFNVNIrGs
0FpetUNM1asfrzsV7Zr7mHOGGKnfEfOqe16+7pdP2qnsX/4EcjZHtozjVBop0aWkP9ULscwGtgny
VGtTkYGeKtOhVAk5miJAWBNYRozQofqedVm0Tsu+bEIKRYjVdl96jT33koSPJr94KV3fymaoBgON
JT1YCf1GontJI42Z7ddxHeWj31A206pdlxMW/Xo9/n73QGP8Q7T/NnM5vjHS72IqtIzW8HVZCi3q
b9fgBUP2kRSPu9Sn+vC1Cc4s0g7VFMnHR6MneWI4ZQHrdiLPVXkqzWWLdEG+b6UWDBajWzEASB7m
TQlbaMR+4jZcr6QHAG1RG12hYOlZJY31XxDoUc08efbsbhsVqapXlXoF3b5it5cdOULLhQO4+qbj
keRXVRO65f9FySIKNl+t19rObNMejsioEW9GW70bjhHUkmRzAPOSMQfSBndrFw0esgi75KBI/iYC
gyUFanF0rG1NbTPih5O2fs5TZikxKMDAlA9gztwuNo7tkgxyxIIqyzgypnQ83BLwmAuUwHe2o47N
yAMdA3VHEtywPj4jcS5K1jJX3ayYEqQj0F0W4lqfIQT7s6ajU/mZJXJ4B1ljH6/kJ+IxyRV0ClC4
xuPms971PIk58yBKDfntlnrya4R45d2hI2EM726wBeHpw5BgAm2lyC70Gil89bZD/ywGZyCKYVEG
/DUFoDobZn/DIWXOTBmqMmIHcYGDXVk01PziT6WyONYKrc/saCS6VX6wCvldU8sppIKBVy3wKme/
xLv1/SWfcxUNkyiB/+ndTwfcUtWkRAjtahgDTXKaWr8NaTrrSXid8wFowbgG5fHpe21Bv3fk29yh
tspfs+jW1bAWtwOdcA9jfYY30e1PJ7JEv8SdNF13DzOBFM5qIpLTJhcRPVdDRqBse1noLKzB245O
D8jpt1E3pd8Nvvkkw3gdRizK9mB3aJwoRNLg6fDLNxijDr26zziLUkbeMblFsQVMZsyn4drQNJZh
Ez3/LZnF5xWuXW/PDvPbEOs3SegKJcvMGPtZFEThdT8/2kVFa2Z9H/iHZHgCKuRh2gmHvAJvQxKW
Y38h8ZzuzUq+JKMlYFcziz9c6Z0LM7QElcsTux7CkNrpKUClEebJmsaxjLI3f3QWYjcKsdddLfSn
ZgwnSymn6egG56n8Qyj+dIkOzxiiDQJbfbEHBWteJh56obq3aE1X0QVvZQ1x859StFLSoTBMNcoN
Dt+T30ZEpUSpsdeWu3+1o0pafge1LrYicYDrMdy2Fnvr3uePBnVzdkB1UW0o9tO9IGf4n8+77kIb
z4EzyognW5TmN+VLwInWtLWwaD1aNrvhfQJgdltiBhm/Km78yeLzO8RGZzrKGKDOo4SRpjDRTshr
pA342px3UzB/GjjLch8b2bKd85AOzrlW27+NN03jdF25XQB1WfndDJAuRrKJFMhw/J9rqp9KNrbn
BbTWNBhHygixdT8w7NDeEI6DtRofmhhkRkMbjgj/0+a6jET11Hw3uOz2WsKpIVYD1KnsJO9dU2Wy
2CYpF06oX6CFFfH78CxeQEzn2JVKCWx1f8U11RiQx/T7mbgb+AS9Ynujq0EyKxyw0HLRC0lagrlV
iUrLkk0cRJkt6kSAaxKNbW9Nnf91lqteGAkC5fmWBkLfchBDtTmy+qdjG7avl+4XrA3cdXVLAL08
zhvmKZKI3ADLrtogTbYUVxFTrdq/xMo8b8uivCMLkPCp6iQ7pvr18qi7y5zpToefRsAbyognFjOK
FGngwT0/qxabljZh76wL38ej+37Bic4yUZOlwumqlcVkCLfLs1jtrVzFzKSAi1iPHxdQtIfkxtx5
hSAquaJTuQPR87ngKp8xOQYbzmHVBAi/kJ2Pi3ujK5e1rYmK9DGMzbLIICX9M0R29Eolubz/LzcW
akWI19+SyskZ68aM35A4MyIu2u8tj7ooKBOQ+WL2/3SnfYpnUbqMmCQgbAuayXDYHBBrjwcHPf6Z
YVpE/N8j6orkkDKmea5cVrgx08ld31gnaTY8ojZyAMjgySTPgeg/TqC+D2kKyYOBrYb0Vg3rN4aN
q15B+94Eo+FL0xYWBzvgG27B0Sw7ULrlWe0tFtW61NZP+xJvom9/dUk/tN68MxS4xWjDtrFR9u4u
d3SKYYEoCRCF9+PNpF1T7lwsn7mc3/DnEd/q69VMiYb9crlWtWV/MP/XZas5r6t6LVLm0uCmmuyw
d5VOGmPRC7eXHkjAOORk4ZwC//PH3JhiZU98Q28Jko/Lpce1K4oGpk9WlSp0+TTxZh1f35H9AjQs
HNU7BfKEiWk5Ar3K0niFOtd4rBsCeYWWRGoNO7QOCwhZ01QU+U4R1ZKVyHmiXchLdK+2BSkSUbWm
qiPvKyi7hukhfc/nRfmSwZsCNp/iFyLYJHh2TgKrerxEy8I7g5LzBq+tzY/ZLFOxTttre9ASTbjs
7ikltMx3zYiPdKt1TaA+KE2dztEmmNhRWZgncm5ZUUXWvy8t3Gg+4aS3FGZpzEvuOcWn7ysl6mMa
ouOV6EvOXw61hpfh4OO8kA5UOfaoK4Ue8v9i1vUal9Oxt6Q5jXtRHLZkZbT9kxsOWhXBT/yKxhyl
f556HmP3Lm0Da2x8PyQX0+N6Dmm+T7wpiunHeA5L8AfPJacryYS2JXXRt/UH0r12v1Zl/z9vMFiC
gfj5e+n3Ra8nWabBS/cMGRNlLrtLAEVuKU2kDsgxmnfqYCnQnq/O8eUHA/fN/GZuQNqgr1XfdfNJ
6ZO/772Uced95gGJ0Wm7mufuKWcg/zbCtMnzf7wBILmcv7azvFiLYwUeNjBlVdYE31+d6lzKWcRb
qdiHHRUdmEzUTGPF1qZ7ysOGRhwHbp5rRdnmz/hZO3zKULw0sAPm5IEBFaBDshxnLmy9RhGinNJc
ebrYGRcT3ecssVUNOJZk5nLkstZcNlzvBJJsxUxuSEeB2QTwMtT+h2A31h+/y9jVP38rReDms3M+
2mO86KiAdSip5On7xFkqUQmZb5T9mWEkk373jXyGHd1UIntBKNDJJ5w3+WxT4nocUZ+LV+vj2IK2
5p6QSgn6BQYOqtLO38RwaRF9B0lQYmqC4nKXrfIWzViCtRc2vUmLmBJTYCO1d9o97j3hA4Me8+Zn
DGi5WWTcu8Is6Z7O7TpQMl/zYX7RZHwmv174XkDCsl7WdN250HzXVU3IQM9kpxQJM11gjKxfRrv6
hsQAg20EucjyLAp9DLaSjVWw0G6Y/hr1abOcbjHE3gJ1yITuuz/iVZiyWsHwx8nWNnXqfzf7gpbz
DVBIPl80C4PvA67tdnYFm0C4+VF3f0oY4zIAZNGTNR4CzaYX/3TOexMGi5kq/TByWt8yYcktFSNA
lsen4+IdET2aXAEr20HwJNFE0rZJpUEgu9bWryWWkEd7jUPoXkWjxIg8dlBFg/kZYJXE8O02uXp3
+q6gDBZoAggQ2pKxynRbPyrYAOkj3vILrDthhhytBSAahl9VscouKno9vYiuAJjp5pwrZdsXJuNn
Rt8qC2BQp2T6m34JdufwP1kkHk063ZYy4H4PC7Pxw9YCqlFzebUh7T0uhVbTUSco/CvRyWlmb4cw
qtBeOnIs7+zsn7HCm9vzeiuF9C3A+lcVD2ppcG+7rfNiHFvXeTYIdeays0TdplYsNJyjGb836T0q
8WfAoHA+xdSYvkgv0mmrq363p3IxHYQxFm8xwQRo9E4tRHqe0KbogFpvvEvQSpyWxnGojgYF0YYX
nAdqyxpKvg/GW4ryTpGF2sQLSczHEeNoNCT48EMChtBPU7DClmGesRf4WbTFRuTXuwB/JAaX/mQK
o5EuH2RCehBdrpAbkm2riXPPOsX/fNbHd5VQHi68ItXrbUvNX3fSM5bF920p7a+03Gl3j193K6VQ
ATf6bhoGAz+cWsNi9ZL9hE+pN17K8df5qymj1orQpTWv2VJRCDx6e0P7QKDYPMhBjO/6hL8FF38t
ZLWBkZabzgckeximewQhDOByVkEeqkkAaNL8FesmR5hqrIERNJ3wHdsnfgSVgKHhkE+HJabUZIWd
elNEXqA5OhZVEcQyby2mT3F831Iz3NO9ya/ywNpoxCcz25CVGShtHAjmY3/q+u481fHlfnZTeTZQ
9ROclv9mbX7MIzfI2KQLh/ayzeWv/fRO92SZlURrV6uyNd2JT9wt6gbj27ph+miAtFeIOiQ3Ood1
ZTGbR3btyfv3AMLvaewiMwYfTZ76XqOsBd5/e6zgrQc//9E+gpZ/oJ0wVRvmN1tZyhLlVf9pV8H8
79jzqHzmmEdItYFzXOLmDd9Om6k6GHloMoXUPh2cvYt30R3fXtozulpUC+LqKTuZNCyYRGprcIRp
6n3Wfjv7f9QsBwahiPlTUz3nxkBsYkBmMoPVl4yS1r8D/jEPIe4cUTTuWJSNNQAgz6nI+xVGO/9Z
jj5bwUg4rNvJ79bQUZfDnClC6gQ2Kvf0X8/f7RBowyciRxtRO4UqjSEiprZqP+hN7Pd6LBcd7E9L
u0chq5/1+/YDg/R5ETAx3AwM+5ztFIWBhe+0/cuJkTW3J0onJ6wVxX2rMgfp38XAQOm4Nz0ALAap
hOY/iyD+Rjj7j1WUob1NxUxv5AbrmjmxAQPL4vyNdpchYD8QDOAoxQ8uaydeXdfQP4ICKRhlQgrR
BIP4IH5cKnQ3gFp0f+BxerSlvaQz3bcbVvNWG18Nzfwu+bg1hI8cGe+CSAlTVeSpyRwlSS6c3sgt
PS6BMgZ2yi3SI9HttBniNMaSMSESN4t/xuZKW2Empb/b3rSL4oq4mKmAWl1VTbILGc+JXETEgA9j
vlgSkZ9uqSu7XU8jg8T9wT5LzI1E6MN5L8FlcgSWKgENxjmvxTZc+0gU9ulvtSNMfYgXUkeoyDwQ
YDCBGPCcD7q1HOnLFbdPFvLx3jO+EeOBHZOUUiRCqZh70XOJ3j3qJ2kT1xCyT9BQBO8zD/Q0eZTB
kpOdTSdYLvuKHUNh5Kt5Y7T6fg5EWDck94lAlZaQKPieZmY1o0PUUhwpLkMlfxwHktlWtdH5TTdA
mTfbLeyZV0+nbcZ0FW0djoybwulaNb9pD/3i4VS32M+7v2fp6u5lWdUSOFuJn58tDTy7U8hcMYGK
la0RBKH+8tZxoHw82eucYaT4vS5075vmqA2QIdDlD8bAV0Ses4i2ZyMkClug1A6u7pRRCm6vle3p
/AsNMpOd1Vc49Eav5Ln3wtptzapxPbPphoqNE1FSJ8ZDtvu0kKD17CiW4ukp7JMgqE+kDgFAwsQ4
Jal9/l13/SQaLb0ggSsKYLgk4YxjHzPoNZbStWXHHsV/bwkBjo5NIPyhzI8ICPNPXAW/G1VIU1co
Ih8fvDLKM9Ii0+VdIYDKqFyOFfUaNS2MkOan0rbN8F4A3mJ/NLejQrrbPkkxgvvZUfQ075yK69En
ygI1/pciNoiRzXYk69l+6i9T8ygB2PLdN5jPdmWtRClVvDVu0X850V5yW0/OFRLyh6H7/qbAWJ8X
UeFqUIWxwLofqHyDA1WQxLuvUEgJLjUIlWFEA4u0lPyJw0Ey9rvVL6//DCbGFT4eU97p/Y4sMF00
4MXMuWMWe2OrUSnwtQPPM1Jb3Plg4MOUk0xNugyS+wfPr8IEp4VUGtpf7Fl0E4v1GYJqvjJ8LWY1
y6HEZOgpZrKWkuBSnrJ9KICfwWYohRhz/wERQTNTXbHZM+yyMc+Uf3Ohf9Z4g6JuDJa7C7shWQve
1fytOXfm54KcZ4enaUkU4uffye5G3Lv5LYftwtmnW3j/ePUTrTOlbKR4WzuqmIUVW2sOxnWOApbL
VUokM7o1mXOE+Ee6Dqfsp0nb6QNy6qaiSGDnLbNblaj1N09Y8EX5LDH+QRfOmfKQRGqgOdHNKo9l
LrqHrSS3wpW/3HN5N2P6RLb+j+82QOUM9bYXyxEYvCf5chaN06jBczDWkPNO0oC8k8VxYPla/O+6
KIgAfD2eBpr03pQ5DfrJFxTdYvVmEeMSoqtcubQCQP7MHa0kncRXuv/5f5kE3jTshh0KaQ+hgx/Y
91Gy9IGsPc0at3Kl5F2YHR8mcrSnlm9F7kSuxItl0b8rs1T+4j71uS9m2/vIHEWVaWqoavutrWUH
1DGXqonfSzaiOJmbsBiGa8YFzNJRIABZvYlUx6Y1LhZXxkA18xEIWpxrCXiVnJLUVyupF7p9VFQr
T3KY98OOqYOYOhzQdwycNuxEWoY5tL7qYDjfUj4A/OaADKZ7ucbsHsfCV622mYzGS1PtNXC1BZvt
dtoUMUl0i9pVJx9g3mirAm/hmRSOb1jhlOWhmC68jQPkjuFed+YzALPyToEfhtHDk0dh4rMr8lvK
S3VC3/j6MK4WR/UDG7P7BmwfbFSBzLkZMaMlB9I3yNQ0YNr9ILubKmgKmQg+KFt7Ish2SxfK6UwU
JekftHhjmCypUC8AMIQpHenf82OfE76VYjbHPp0X2TzLMJyRMSmLrxVeoor/Qcim0JkI1Wi9IlCX
OHlirflf/pHPYzyYFAsVVk5i5Fvb5/dukgpCyfaDXN7/IXRZ/C1iD4HSPny2kf9uV++LQWIy0LWz
ObNz2zgdPhozO/grUtnzcXIxQjcTaiql46xAH2IGZXjiS/1sGpHY39MYOgWbajuMIt1MlCiqcaw8
0Uza1Xdrq9/PRn8kEDMO2kufsIS1bTCPdlmK43FNRIGz8EMUtq+5uZ8RwI4lILDx9y1aD8xirsEh
1HO02iRehgTlVqB1V8pDaI5tEmeN1IvSEk+KS3Talg22o6OxNbKhRCtxhip7oWPAOQTLcW9NLaC4
XVZtIKl4z1WjznrHAGDMH0jqpu2k1fSyfJ51frU0AGojfvHLvXxJfvhcjCRdt/niYRMjGZ/sHkdH
PBw1swbQ5LX85Hruupzv/LYvU3ZKS6xrdMUxYpNDf8dP3aNt8Ge6i1mm+n2/+G6BY1tNxhDZ9yKG
oq9W42ohkBzb+T1fKuaRk4IfvdwofJadOe58ueJLwV6cO5cWA0iho2/ie9IUwXz0G/tM++8ttpVd
fM3vnbmOZ2xFpo1oXXLhjb9E/7i79EJ0OAp2En8S2Px30Uj8w7oGY+OcTEcS9bCv/izEUCBQtUHm
FpwCBxn/YybfV9VsqqoyxacGbjhtO+8NIvYUj396gBMD0V1ZJ/Xz30Sm5/yxzKlmK2WK1oHtbJOr
m9jYPKeWaCnLpTx6QKLwLp0wXC1dOWyId8UjdXnPXTIJ75hMPZhFehq1oCEjF0inDdjy5oNoLo6i
2MVedCykjSgJvVyJ3zb+BI6nyQnvTOv/+p2/Ggh50Z+nYgqelQo4Vjkk9TO/LbzXbrLRsvkfq2XW
ZcxbhE7SZsxmeaGe9d8JHiPLlwWWNhMWNz3Eb5N8L/cS9Al0kBORIpvQEMdpcSMDUwy6UyfWe1rK
taaU/WRT5QfASbs6K5YAROgyX19nmGBPrB/KsvZBMx8MbA3tPZ0QwjltLmz9MA+7CmcEyHKeyveY
o6qgygZsgYfpHSu7e7WNwUqNLDs/Y5WJu1xSryvvl7uJHcoDXJEGG+1KnOdo+buC1RNGqcO58Vw1
EjIAjiAmo94IGCOexTQKaB9vDseTbcAtn/qjp+vojN2H5CTs7hce1gF2WHzSF7PchtBfzl98r+ds
rVRBgw4CwtUhErH/JgPeiYeWcGiSbERzv93O0MINizrXIoGuE57kXopaailE9Ges97++e82vhg80
aFiJqNGV2gOj8bIaEzVIAiFquFYK5dNRyG5097XrLFA5w04mRdfTLSgbFqT3dnRlqGQ1SLd5tFbX
zbQ7QIpymgKXwoVZibwiIud8cZoV3FEtCVMKbpv4Yps2lR94TnYZTsn0b12u029NCxjcVUsEhO7o
AD+oSmhY6pBnbet1JxvH4WQsIDhhQs4KZEZ8MB75eum0IM477j74AcDGxjKXiME86vYMaCyJad2h
0Q3n8z56XwLKSP5hGO+jOcv8SzPUEuZKFup/BVFjRT9IQYUSWQIEmKWyJ5II1jHKeldZe+iFHIL8
OqdOYo+hLQPvIUiewy+F2FBZDNXHJes6rIgIfZ8UdBTrlLzcMTQUBvA8Fdl2PnJfQYDLUH+IZ6Qw
sa17ehFcaMxMkPYN0gv3GuU2DwsdTv0jyKfcJPcIOnM4uqcZu2PIKlBlIB/Mr/PXENcEi/QawrO5
EvrteGHzVhglC69XD8uf+omf6VzKGuKndT/tJzNus3gQZFgZ8Pb3DPw0nYKeOm/3j6xD5xmtZE23
Zr1R3VBskhkLkFsCj5cnUFcaDTITAFLclxOBCc8ob/QEomo8gKplLHFk2XzAtcsUt3dGbXm1Ludo
SjpgN2OcekgZ7U2m+G8Efay81PNeeKoitYo7Qj3W/kNCVKJnFARaPaW9ipl2xdgv8/04TbC2XgWk
+/W4zqMUvN1a7VmuwG4lJDzj/NZFl1lSDi/e6WVHLerPTh9PLhz9XmAMru3yl3ilKgj22mi5OWlU
hFg6FfwbvUr47adqn/brL9OpInjaVzRlUa7/Qdys2UM8wsPfgfBFWZ/tbV2jKng3xN+CuAPiIdxp
KyMFdgIiY9Y/XTdn5Xl3v/vbJRL63WJc750YBxb5LY4E0+U92oercaa4uVmEggQcms/LynMXMzzG
kre55CkIt9AQz+8znXdCY7/HNxXN9hOhvmkHZLaks0yDDT8+NFsmhEgZYkizNKVCWirGvAEcsgv5
X4SmaSWGnSH2wj4zS3UvHphIMrAqXA4MDtYj35onnBcxtSkwBU/P7I17WHMCo9OB5xsKwrtYZunK
VloKGPWkctzk1NB/W59DwXNFYaFe1dPIAyg1Q1BjCqh4DEYKe7+betadyo6hkExEkSbcG7p6abj9
/w/3z7eaWnt7cFaJDHRSTI8SwQbYEMKWit5W41d9mHPgZjNGjEHuvGq/sluNzYvErUh1Fu9GBKhC
GHmIbAdH4lQWJQTNTXUzYtNYcMQzA7YOL5bEpcUaIr/vB4YgGlcX4ksVdP47ycawfJjoaXNaqYob
JUXYzv5mCL6TDZasWFwd2Pfwmwt+Oc2h4AURmXrrwgQt07NcvSTi4LfgaB8a4nubPH7a09ubqtcl
pf5C6K7ylSHcVuVFhcrNoNpeWfTg44MPgVvNBptudwmzw8YKaEUO7vwVjFUqZJVkanE8OTtYox5T
N5le7KXiZm6chyZB0eZTlw6CxYVWPdscqsNOlm59Xu2rzHlI5xVnLzBIpg0StFH9BU4XI2g0bYOc
T5viYvPuXQGW+1eMvlyU7lqYaFGpqWeSy0nbaCpIR+LgW6OnH6FCrd8Ewx79UowFxp9mzRHltfaB
Z9lxHt2OEMY1PAeiZxcDu1+oFkzD2H917gu6aqHgjfwKiEWlSDVCPRH1FVuDnt0cPElTQh9Efd3C
HMXSY8XzxiJHFsEy4s8vGSJIoKj1hPeuGRm6ff0QhhGSD2+iIPhR2+BFdX2olG86eTS+RIDCc0X1
9ex+98Ir86hGqnyfDL33j+0bjrQ1TXFj3uKIegNRlprnQLx9vDD8OYvmq/84sIfcawETJEc9/U40
+fN8dZitqYGmlvfOc7JWcABWCDpHfe5SwbhlcOecWP67wnwhJ8HoljPWqXspWGhzkKJNDZTmQNeK
wNU1gXngIQdZH7I0v+2J+8eFdrrmhbYERw6jDUCgJYPbXOnrurJa8rjBcMge2npV2CB5ZybjVFfD
i06/hIS3o4odePgnH/tWrgQb6l4pwL+nyJjpTaOiMSFpzBq3Y5FVhjBRaeWqJypA3HWbrIQ2zPss
/URWlsv9BTFI//wmlaBUTc3RrzmMjEONCzYwPG5KRYcK+T/4pS9XMg8qq7Kydk1l+AoibvKeg/3F
HV9+Cgpz6JzYqxvCvc8Qa6P0T2cncdh9i/AQ/i1pqDv6tZ3+AZFEFoLS1XVZg/RYKdt9o/13Wrwk
tKO6MyYfyT+gFDFOAHP5ppwoQS86Ks6YxH8FeMhg1QtjuGmTQsHxEvhC1TC+D1wSb5+5GiC6uANd
vwsd3xCLD5xB1xHjmOdtozHOJ8xgiQCMayjSX1KnBWp0G07+6S4T3THJyl7vvZ6J4IMMhQrHkRoW
ZceuxdScLaz2TUvdNGdFDsVBAE8Phapxr7hQREOr+ge7TUyJDCyqfevdH45dOLkcX4Ldd7/3/DCE
lkoKm1C0YZrLdwoze5F7l0tdapT7SAIkIyiUnmbTjjiPqffDjBZ/ZncgsM2ZFVByxlo4U9LkEU1g
CLGwmrMKTi6Op8MzvWCqalyjzsfTk0Yt3bqG3uk4vNMqx2SmMit/gRtWbAfKLF5vmUZF1Glkohb2
H+WCBmEnemmf/LMV2paFkcoiHCu1YfcWaw+WQzI57atwLbctnwqfo+/uLATTQ5R4zuPAb3a2o0PX
Y25+WFl0SELn9Fjkg30X/rDPhECOj/ktX+Mnb53bdU1wXxey7ph8IzjoWQovTFSd9HSu2Rl9ZEh5
voI6Sr2ZxvR3Ftoc5cfQhT4cxyUSykvuto72TR7WoqzKcxnwkDtN+y6LkFCZpNa9dJ5WJeuZHrCS
GpvMpISiYD/EADKjvmujIX/kw221MGnoe9B0nr/s1Km20ZNbxQeo46MLGCaXg6ZysYRF+iBK/Twz
14zI6HU73FSSFJxYk6RgLXL+rRyI5SmkECAUMnekURTlQJHnOii/553CVga7JQEX2+PHQVwk75kR
toZM6GOKiDMVozVJveK6ZavStlUFbMUOu70YelC+Vo9Rl39On06D+ycn0QgEUXvogtiy9VD1ElK7
SfGtPfayMfL4d+aAf0tuPxiOBpTi71p+z1PUCwXORsEx4Ur77ACw4mg7wYPvF7hlRtjeUPBaJMPA
pcAdJ8CM1TD1wD0EwOCFAR4vpHHQOqfoTTUXMxx6k+YvImdNUnh1q5WA4xxtr2CWQwG/5khYc5lY
2S5XN1QrCCr+WPjOvm9815utYy9KrPnoIbAW1StYGAUnJagsyn+mrqobQnmrKG34pQq9l/zsmBom
wWuhQtPvl4BazyvF6zsnWvxPiJn/MnqlCQPS/VUPWwVFzil9hAl+ILcaYHd160YJI4vhySymRUKo
aGaYdhjzYKZ5nwlnHQ4Qs1k8aREOjmCHxAj3SVf0ZsR6OzdtFplNVHC37iqzxrCTKOsOtLEU82e4
rPUHq4QfQvAxa5YHbE4IxDiiRed8ylwn8FoJBU5IJMhhsXfJlFUNW73dcGWncJPgiH6VCqO8H/ci
bJvNIu1/QlEr17IseOD07ZxQZ0IKzjmasVMmSyyAJnu+8Vvem6wFliT3isBpzYF+DqfGZwUFuADG
+nqBLyqoioN2cMvgtGyE+nd+xMHePiMc4n9V677gMGR0S+n180LKZBmBoEeBO8XZkSTuU5q3hZpP
WR2tlc6X2FnL50FaABxefuaU1rGFsI99/TgndnTm1IntnPQzOOkcbFLrAe3cO/FmADqiIDZu9GPL
KGwxTDcjMXw4z1oX9sewEcf/boSxoHybSwHgzt7UUFynKrSoO1i/Fun4yoqpKQPyoBgwj2r7Kq+5
VFZcMvGcZoSp3d7fM8wF4xdP9en7OfYTfBcJ2Cv6UVA4Ow348RliStK0xZ/bJz4Jrm110pB26eaM
EaQfB9qC2oT9CuWEj15djcFVNZTZIAamCusH+gXO8sso1v20sIRH/pDg5SzjUty0/syz149E3NAT
wKyLZBg489VJCA4J3Jj8Bh0xQiLanLYNfBbuEQ6wnysnB0se9PFzfhYYScG4abXl6rVihJlcX15u
nlsNVv7vHxBCX6J3dA58wsZk5+mYiVEaiwlzOYvu+lDvsiMahFv7DZ2DPwWcJnlrA+fXdH4AO+dr
0wnW31nuKpkSG4lFYFCJyD3qgHmT9x+K+/ceLPbaztGfOw2lXV4DISpm5t3ZaSnn81H3KTVNzRce
VavW04htnh2hKNN8aJdnhyVur4b5IvS/rP2b2vDBWbypMzvxvO8FtPFK3VcWWF7ozbJzElT/rk3o
9nPgdu/HcIucvddgGrjfVen3SdX8AGliZYSwncc6qaHimPyJph96keYcVhbIICLW3xHwvXPm+Pd8
LUrnP4FqN2zsWZHDibqU3Sprw9LlEznTeq+8UrAXxpdoT00woUnOhxSLTVVeadZ6LoZlPiIPheht
qLmuX/0MoTGorvyj5EEvA3Bfh8sXrWOTdFQD8KLdL0opqlim5zB9FUQgYOPJaAhmS2h772Mey3ph
7VoS/M9fsi7izxM2/wJp1QWNC9GKL/2qvV6lyWYNvAHz/fFGl0q/8qmB66oMc8l8BnBR1JBsWwXO
SKRjywcWl36IL83F9kLBLhHhtt2tgjWLlkm3+7BN7gDW++cUlYn7ZwwWCZ7XoPbOiSaopWRmAfS8
CYo5LrJt7vVQsTxtB4Llo0e6Rqa72ylaSLqqE5jy5Xil0y1fGH2bM/DHMiefo9IbAOCrCayFFw/t
VVITtmKV4i0UyemhMQjR5YDvb/ATLQre/U0n0rsQKSvapN4tv9ccu6XPCwIueeSN8b0wgb7qyV6K
88KKFouMeDB0BNHLMrMsTzOzCnARGpeSg9Eiz+yA6Jn+QE2SexaRZwszFXWhWdWAmKcfeGM5aYB8
S+vJh5RlaotW/79rcbAE6pITJ7wLJ4Xg/uBGxxlD0LUZ4GMD12HEZZ98y0iOD3hDiw0eRCUCVnOk
+o7xhMchYrwUsztBEgf+cFKThNlHaI0rshGJJ0a+2DVBJMwLHEecKtkdCNRJZnNtKx5Dct9my6mb
UCmVV108u8XHhvymF610Nro3EXnyvdrujZck/zOme9mFwVvk+Uf5bRJlpFJRX9k8uDcRooi16Nhq
sAI0xprZQnP0dwdG7WLwd+QN2vhE6r3oPs2s2OX8odzmql1jqMHkDipQQ6OjGJyLsxNo62m8mSUI
D3XF1DyhvqYNjfxLcmYmzfzV/ZuHc6o+vFlYR/67b9yKwDKJf2tudABbhNg6+AIgf5sMmy9sjI7E
9V83kHejUPQN3ckJmJQZ3dxpum7yX8d4mMhWWQc+awZSQf0BjhUN3d5g5vrctliZ8Z7fw0U1V6/m
CRwL1SfqD5uDjmSC2TpvsWsYPlGoviv4c0jwybyaKt2qPgsdKrJ9Q5RW7ABk8EEasKfggwvwUZc7
NDwm61TWgEU2o0dtk7OaoP+tuxxMoQXi5zK07DAKMnZloXBFv6wq8dpSRwmxKT+bW5PuKoN6In9p
CFn3lvS3KYzWP1gGwxePKfmLo8chmv/Um+BHgJSqeH+3Awxu9Qfay0CKhqvpaB7EAoLEbyhmFQIg
5fzhiBBzsAvFmolim9WW7Lq4c3eORwryUBg93j0olcSox1mQIuxcT2Rm2TgtAB9qMqckqq0cKE3F
linCH36B5RSmu2+qCT4Si4nwVOygyHSkQ5s4Y8IFeWZiM9sQlazjGzoX3A1iX9YvY/KOSBVuXYX8
d4K02A2xp1zyzIOp+Ej612lokSfwEl5SL7uV4AHhJkFNOtgRsNSrl4GLGoDdddb8ELyY4DsAMfip
bVr1YsMHCNSyLN9laoJR/7RZ8kXf6RfJOVn0fCyYk+q4+2OqSNS+ew5xxDNFysRv9bx0oM5rV2oJ
cTVSAv0djcRM7+kYfVIoHHU+g/IN8V76Qqoj84RDXUg0GMmM9By46E5lPmZnTyP4VDlWeGpmpDyj
Gacgd5LNq/DuUyFOMcY4w7HbV4n/8wyca5l4B34KG+R6nvKj2Qf7N2duD0JffDjXiHKiO2eD3Kvl
6Wkgwy/L/zJnC5J+nIWpOvWaWZx6T77waYTZiBxssa+KJKhvNrKepIihvVheC+xK+QRvIGjzvfo9
NipCZbz0rDgCzgnAeF9/2TOudwKGlGH0LDdWxMH38asOaKXwP5kiuleQUxFYp61yPRMEYUmZyg5T
nV7MM4W4l5hqRYC+hEhC1lreyHzaFKsTrdGJInn1PoSPpd5eJnD2AoMzWWi8WD5ItYsdzbwOgPIO
hBsMooXf8tkxR9Qg65dkeYP4BZseM/fmlkAMTQgvfqss4zL2n1cL/s+81kW+5PQTBXgKjLlDcXQR
UEinSb80GqLJEN+dDmTMAjk3nsOqTcGfvOPPTI2HJTeFpj9T0r6N/JFHpjQR+RxKBhKqTTqfeha7
aQvAAUsyr9ynxxJkXnKEPlCAnrGyE5EK6x7PQOerP0igz5to+H5+fJ5nOQrNyS7s+TEO2E+CiE+d
nkxgFTFi+zysMIzVQi8SmElC940KPOOJb80T8rtpir3K631UqapejvTLQ+roPQtnrNKJDKGk5lSU
u6owC6Pylt3p3GwgSIjW+Kz46hJPlPa71TWtfy7E2We+hAu7Jq9bMcsidhj6oM2FaxDMXQakBHTS
pbhkuS0ZXVxktjLw3NTrQcrNghOj1YwEt8jxvlIQPxRFCIVGLHbnN2hgO+6IdEkJp7pcytD57Wt1
kgJei2AxsxV45CY+cD5P2BNWTmge8iaXpq2ZigACiRYOaxbf9gtLTGmlsxBYvYVWQ5jrsl8DXJk/
VAN+KeuSbvV5kcZ2rz22XPIXZUOlE5cTyMFgcCXhoTIU6N5Bmm0dyrg0iDsgfAPiamibrob5L76t
3JXp4Cga7R6J9FNchBDRPwiPoaNNSj93sRngrgMRN++iXhGMGQ+7gNGYH9xdAnbVIQybOfSWPp9/
GXUKLZlPnwk2xs1jy+E+iJbJKK2akbJYOPCvW6PqXQO9u/t5PgXivIcuFGR8RnOKMUUatgV7KgsD
Ks+JyifyfsDmobSJdQH0I1g7jj/LGMrz3qwa1M3Oa2Wnj58+r6CoNeRmgtRqeNFCx6msWz00R46u
hI/eXxp5L5VKAm9t4IZNcV9v9HKq7k5obupJqbdI+0LXNleyowQLxwqgvWlkzFn/bqG/94kX2Jey
KO3ouYAABEAyUc+u0pvExNG+Gvp3RbM5CEbl3tGRyrLKY8jQ73nWOa/kTbxhW2yZk6wt7QTevDT6
TRsFXORjY4T5QR2b4XGVe2V6k6RnIZ+mtKdSpVZI0N5GLlGc5O5YFoVrCpImVoMi9qmLN3K8UKA4
VyP2iCx6oBtdsnyhOLxHHFhxw0X8F0wbfN13ksVK15LumiucwhwGVv5/vx9SEcjXgsIMa5jpd08D
u1paHRXUA+dCT8iWjGWaQcmV0Pswl8uORPgWrlsyyPUKcbQ43xl9mb/eZb0jLiBHjxlqZOh3VjQg
ax1F8fJCk5inRlPrIvFWRf/uzEqDeibkhsgY6zsqRkueKuF5QAJVLhgprhdDRptcWpuX//A32CO6
OB+DfwfKRXfEe+AA0lbSNp1zJzg3nxXgIwDHhHYAdJZiyQSGlHjYU22RluWKm7vRIA6lUua8gyp1
gObtasgPmNXr6Ak9bgsQBk+m5COf3tXCtOU4TV8AtKnHVWzlA5cTNMmhCGLJcyGCfYT3Gc3URVGL
awRo9a92S2Xh11rzzF+R+/yp/eyQqSNcB2dG0KhoCll1Oh4usQ0qMOjSFonmDUR51gbdg1c8VaQq
vn7edmpA29agdrhiZ0j+jtLUAPuUgqBd6nb+VIzgs044LJ1xte5hMxU0FkVGstfZ+6Qq2/7MDouH
tckXPqh3qy7wJRggplsWVhemct8+RJBkuUYo5NKbaXRjGnV0EKGaqSDBvThg53Z8CfG7QfZYgDOm
rBdpzh+4m0UkrhfR+kNXNzXcEJOItb11FvDOxl4rLopJlc3Is3KBLcPBHchl3c0PGkreHxAuUfWU
Y1hbJoXGua+H1evFrcgBrcXCYtlIQdyF/lvU/AZH+9E7pHMMZz5mSY1YpX4M8LgO4eP9nLk9777c
tETezgVN8vBk3fmjUw4UNPVXb+FNbnKFwHCGDEBflYPt0/gzJFhL2nB5pvzWzmFEqFO2ZTPVtNGz
dakTX9Zau0VC2hsp8I8o4Z79LHi11uBzd1OQ48UWys6cBXC+Q6YxkYmB0+nuJSmGAo2r5q/ObGC5
4aDWYSYSFZaV7LfG5C7/LhEzHkM9ZW9Ucb7kg5SEduxsM2aVgcoy2t1NeCPLpq4jPEKvex4CSkkP
qwlrA0gT0ERJrn1UO71bYX++ss8VGelR7eaG49dtGpLSO9mR5s0rQmzmNgrPF7ivHJNPp1yK65b+
Dv+Re4UmbgIwloZIwIEB/m4PY2qu2XvrQpZos4c/GGHCPOmRrBg5MvLGxhOYkirec+jOR4OEgbB8
TtWJq1QpqPn/XhcZ5cudEto5YsfqDK2m8/zu2ZHKhB8msR+QCx1nNX2m4LWIVy/PgPdWgcxUIU/m
B6U632NM2CyHj70+yy8OAJFWLLSk/crmbzofMvBNIYkQnHeHb4X+Wzc81I7sONQd7jN+DqxJZKkV
G2EeFX9+ZLOkTNCZgcflNQ6GWXnokypVt+4Zt0CuSPNtzGEhty+/Lp4luEdO516ZCUFktD6IPLFy
gzbrN7l8QaHcOB4ilYGoRclQSJLi9815Bh4xJLOLJmTVi5LkvydxSSDmlrfr9eT83rXsxwSf58+7
VG5tJDmfsfoag5uUQl7ozte0rc5/c69YoGzKbhwEsuj/D5J0jRj4Ef0i6OUS1uTjdFoutOf9u0Dh
SCOmHXEMtzlx8Q6xkBJwu+/ArOxAA9BzPTxLL6yz6fWqhjz7fv00BO2W43Z7AFEKlhxxZCzCMur7
9cGjrmf5ifUdXAFose+Y8aAhhwXC/p9L5A0MAitxZRGZ1XfJupiJWoSItrJcsPLMXDJyLlygPKp4
ovJz4R3v2WXQoI8RkWTHNB2ebZY9hUXkEXuZr/er5U9WNHSVU4BUlk5BRaqoafg/mvEY2JnD6Wt0
Mlzn3hmQPMziOsVTJkX0NS91xS5FHULLWikjWN2ryCTBv4APx2dn1nmzCRSFIVzoGonTOAnMpyl9
A2crHHJ4YyziFr3B+0j5YoJb0gT9w26yJdX+Pfbaffgl4KsY3pYKTV22NtKOshzOc+3HOZwEw+hR
FOcVeqPJOguFPiflP7V7NXvihASr+B/l+cLKe2qSo65swSVNrwAynZPNqMoVFJeAVi48S/Z2+87O
Hretc0KyOMxkI1vSEIt/dpeTITserggpIo1XFn6GGXt2ffiCeTr9w0neDWdYr/E8SU+sCqClTvHt
F54D2jrqQElaoOMFREdgg3h+oxBKKhLqj53BjW4JcEDQEUJrn91niCgc0obWXY4sx6y1XuJCcwjc
zcH5/uv8hOuHU2QmLHk/VkCJyzP/Ia4sUpIxRGw7ecBUv4SfXDsOPNzj80OuLal87x/QaFlFcYMk
8ddLtKn5Z1s3i+g3S3s3ulRYE6pvXvIJfRy91UcUD77QxN1v4f2Z9M0scnMwjGji9axhs/rNWBCH
0axjZN0+41Z4HYCeZDnSm9cRC+sXUrMxp4hKF32+N1C4vBuNMaqTKYS6J00HN0T63GYc7khNHyCD
XTHWVM/XCrW4BLVydWDkiVTTa6YM7b0RfXpuYxI6Qiro3JnaughdurvS4fJ1xk6AM+zPH3D13CHg
gIaFqNtFpN6vcZ09mx6IjpGkkJjyifzXVVz3Z5wkoXjxvS4KmlFZAsVk7/9N5D8eoWU6OTPgsYw3
E/DzOCx4s+nnyJRY3ki0wvmiG+2TZNWhgTHWWx4BqUKeimDnJIKgLf3FxdeomL576QNrE4fcCD9/
72xVVQ0zVGdBsFOza/Bayem9z9K6C2fAydcGT3BT/bmwoubmYfLybHeljymSSjWtWXTbXLS6DiR5
Cm6DJ6v6puqOodq9g7qTDMHydOdNZ5MH3W8RHcVd/YLtQ0O/FTy2JcBs8G84UUvAGF7RhQIgWa9i
hw+BHYFqsa/LU8OWO8mud5ssR3wIr6/8GmcStuYaByFCpTX5pvFiz++wP5QKwSgZK9TLzFO5QfBX
HqXNIB63Vej4hez5T4PZNWlPPpDz0wz3LVqyBGn87VeO9BWwoVHd0wDhqeWk1FmpOM987GFzGo/W
pSJ7gVnL07b2IkOjVKJMSD0KsQxVPdG7YkvIWvsoCGEBacelKhdk7fyEnygh6arOUL6FupVLwp/Q
hn/JuHdTIW3HGObQFQiDgaLb/XSD57SZ8C9Uz+5X3BUnhDNL9WKAK7zjFoJjrbBLZOXyjVdJ7ACU
MGTd2AyrdptQkphOvbAYtZItuIBTmBaTr3sKDRW6P9YgWr5GPNFVLi3VMbAgeG4yeJI6tCYaNQ7K
MWEkZh3vPvchTgCw5hKOP4eu8pVYFIFZKyBcb+dF/ADZBu4yxXC75dpGmusK0U3ufEjSUvJLmmnZ
0xpX9XsedOSMLuopOX5TUpiIn2qPmfnK4npmlC4r+qMx1+0zZyRE3r+r64mFtJ4Ep88BZqj645W9
DNTJtVJ34Nr4fsh7rQthcb2yf/n/vkm0pGZFU1saQeOwG2MgwRf/V/eKzFo3/+NmHtSu61YqA05b
13ND6Bv+aoKlGf2vmkdRWZaO4/Viw/OOONMGBNvrdiOjIiocmXxrVT4Lb63USbHfAd7EohgClsMo
mb21zDIPvmWCUBUvpwUudPFYlIewUybJxgWJfOngIZlbddJyDq3PUK1nwvrov+/HgSAmpqf+nmfC
Ln1UBF+So+xGPasBNMLs1/xqxP+4+dT7V+sQf/urYFAJtk0QaqvujobnwfNwej87hpJq86+yMAGu
kS3sM2hFwaC52050Iv57OxiLD8LZ54WcsTdJBfquTZerMD0kHxVdTWGuH9UrvFEALv9GYCiLBSXP
79ZAbdVbUisiP6NJhI09ZcIpJH1lNkzQdIzuYfE7wQT645m/XsldvSz+TqZ5kZfTUDWm0+rkXN4w
Rn1YvnNm3cB3VwQ63dE9FZFchV8obMexee8gL17q2UQ9rAqeZ7gtaULQlE4ZhkmkArGz2h6dHtKE
s35GDpkybSywKCb3IhwP+Be9G6i3IuJbyS5RW7oNSpHs/dxGZRFnoS5nH3bcselNwIPmP8ApuREG
sq6T9Cm0xwQyot0aDajsd0W+h+tjySNgdAcBQtDstY54FJPLMUZjkW2565KlS39wpCYDrpjemlJe
EItmrkkxxebJpmWFVpXycxeOfVIs/8eCdzy+zkXS7L4gOOLL28h6Vy01yf6+WWN68r4x3GkdAeev
65X1HAS5P0qZ9O0+tJBTD+In3HjLfT1DEX02EfUKrGbIyw3fDI+fRwFpqgz1BMDZK76J7Tis1muz
9HkrtpQYH4awAh3Q6Ru1VWD1A34L027Ma65NF+grF/stcma/SA9JqOPTh1MWwJRsVLoUTO23apeD
w9zgArPrFSIi13Ls/6Sy2E4EF/UR+3cdVRl7DTGEvn797Vc9hdpEVRckhhFYgRsx8C5IHU2QSi1U
s6rcbeGNnM0i35Gx68YNOm5oEcQ+kdURJF4qhyiSKjPr7wsPq25MVQ+KwHg1RjaXWO3QSbnrYavy
qYR2eZpTZYL+diElsgCAi2A1pcIc8Sa94ibVZvvXOSOWSP45s9m68bmFSqpiFPg1MDd6MG2FlPg8
PTGuxVmxp3Vq2+bc3iIWcPuyrLrdlTcOqQ80SbGjVxiA6KoYc2DDxosjopR3nxhnXPDvYH6kSYxs
tzvWKLgUlfXUf5OyaZx4Ugm76F9J7sHliZI1OBGRFyUWEDmA+dR00NEsammjPsm0+dBirtCkZhXg
5Rx85/Tq65g1MLtuRejad6zenFR8DxqTQ0U+ir0CjGTfF9ZkoW6ysO/r2FikcstOEOFBZTQIHUIw
ELy7yryghOdC9gFaK/6r8DqC95hzEsopWkHGpZp0bRF9xhNy+Tpovdnuf21BL9OPcWss1v+/3CFL
81f20Epo6C+kWKhsgXZ3juNESa9TBKvmdJrCTsD8JpE3J20Dw6bUHKwVei/x0OhfKzY0QJe7UVOf
eNI8rvBziSjJn4JNDb84gv8Vf56cHITVC2E12hZu0rin7rab86FBXF2WQy+6rVAwDx+BxXi37n+5
/I1g8Z+RvOBFC1Hq3bwr5dNhq+qBOdPoNkhYtYk6SVaJu9YnBhOPT2DraaWVARuIjq2wt5O06hiy
1nK/6tQvYNJJcoZ73jbxc3yS4Fhr+uf6AqO3nMhk/xS2jZUvsl+9KwBTJ1y36hqB/cAK0i7Nxcwt
mesk8utoGZhLEXIl+ucgDhdLmm32muqPaUqKBy6y9X+OQP+5VaUPOhhRI1Sy2HDayNB4SEnj9YMC
AtbhtdeYPSKiIAOjgO3ecXg/5TrLKHW6UVVsa1Yg3uUzXVLGBQ0sDRzdVQeOb5ZAX8kExGkGWhLb
maWOhhD6LRSZgxqfIqiJ4iLQcVeeJFAEF65ezNwR68XcszkgYXjCqDbPeakGd8DMkhiaHFj6A8/e
4HXvLAfKJigZrgAdu8iNDf7RlwGWw1fdH3OGUiUkFdEYxlYbNTHav7IZRI6t2ZZ+NyUefcNOqUYp
kjnJy3vSzKkLQ6t5Q9l4kkz/sJqkyTOupSsl6Xg0I1P12RJOv21d2rDGNmY/xW55zOv2FqjX5eJJ
uvXgeI0ZQOIPbb0UL6gXYNaHMYFaqKyjzUNJjQ5NMfEupHrTZB2hExphwXi6o4rypg2irvTOsaQR
x73WTdIp6JY+a20dbJgJV+qH2KOLhNbFUgosuQiR+zZFPzYLpojwHPRjCHhsAlvnSLRr7Oiqcntb
ciLI9EVlADW6HHfiXCPknvgPg6lkUk4OGvXESXl96pyr9ssBOAvea0i9wZb/2FtHqKJqNQC3rP+Q
tfo5YcKCv2H6Qjbarld0WJinw3dXK/DU7flVCeR+rNZ8QctVNBEhbgQ2Z5KiQEZQ4bdGMcZUuR3K
j4LDGX3H3LBDjEW6pGiVsCDFvJDSCAUoF09KoJ20vizhD+gziL2xovfT3Ew1M7w3RRxeDj5cb1/s
m+jb6uZpWWztSTIzCNvURFuZPvuaw4LwtGLNv09GwU9k2Y1jchQeYOsdnrxqILsRyL4UPQ/mVvLx
AEGgrjjWto4d/ybFUEhPK+D0icrMYkteDjULb+uWcOmjOSVHHsHcuNcznos+7JOAZSsO25mJXwhY
GGg6DYAtTS0MGr0drnXOYaDDsF0Hu3dKZduFNMEKtxx/tbSM2Jd8xMm8tpJ10pUtqDtCUznbu7iv
UyNPkWNH6m3XbelR6hl3LyXVvTT4Eb2r4oghlQPI9VGz3EzknhYfGvFQ2zxmF+iHLvp2dLQ3vl6P
c/w1DZaNqhC8NAkuc4lgXQN0b2gIfl+zKxjC+5S6qKg4q2kCuDep/YGo+60FjPGGohfb7T6hVTKE
59NM6v9X0rhwGFsTNwsXMAiYbXHVdtp8PrvNfgLChxVfj33OdFcHFVdf5NRq+6w4zkCbhthEmpc5
dVp2dJLI4++xZh2uYb/KYjE0VMuxPhdWJcSf+zub+hL6T/kP7SdO7HYt/oZEKq/hGEFDro3RuDXk
LGU5jM3ctijhD6HQHw4/L83b3PH2gci2aaPsgTi7kRnruuRiTDSQ74I1pfZh8LYkyeNkLJP0ojwG
Wmkv6JSlkvPJBvOOAcSljbMUe6/fZGwcFodIK7RlwNZuRtvWwv3BPSwl4JxcpVfMaOn6LHBtkHD6
GA2jmVACbe1x26pzefTnSoGmzcrzeeLL6ipnRyK8e49vZlFVFBCkAZb2FV6VULdsSULBy7WM7IJ3
UvhNmfHN0UVFr+xkBUSx3citWOTwVUUvbnq01Iu5npyAB95v1t5DyKSTTOTQU+EDwN4X4JL23vTo
6HY7tEClIG5Y0KATRv1x8PlK/CDUM6NL7kg7kodUzr/MAAvGbKgd84NOR25QQAMMk2/wpY4Xskma
cl2nulADxHWA0YcjsZJpAgSKqLh9yEgmuwFl2D2CcuXMoJw4r5CrVQD4J7pMxsa71o+cXIDqL/EQ
Rach1cnXekVfPiwIV6//nUYennPWHNP2WJXcjY78ttfY2HMRudMmKSEnpOT58eT5dbyW2w6X3kxr
nJgmTT9Nw6nFfotuMlFiHe306dCOKRlrZkOj3zUTlDlrt2kbJ597VtNcqDZHLTP5OlgxcRKVEzev
YMN9FMzmEC/Ymv6+SflzhHrIUIqYWOGWKNcSr+fpsACWGC0DKFg3FYz4MAHthOCVMaGYGV2JfcBg
vX0qjD48bGwXdbo+9v8p/xcA8jkw6lHPPf+u++a70plduTamw7m//tdl8tF9j5urrCmJBvZfYLkm
ym+gZzu5CO3Yw6suBUx8Cvr2GwwhG/9j1OXgiXMjbowuLY/BWZecrk0pEmydx1X+YO0cXvcuPzfX
WUMF9Unqa9Mb/GX9WloCUGnuZpyymk92YJpOisCXEcooRQW3QzM8lAtB9DuFE0FHL+1TWuOre0uj
Lapgmnm7LNRLzYk0Nk34ACGHILnEfHUUBFbnZh78S/U1LE80okpBsOqvaaaMCFFueV6TcAKRKm/r
7srC5YsVySZXKNcIZfWxXO5Q5toWseXxqwhT8RL41zV84uP0ReaxZ59GYBFPq/sHBwJ59ANOEfor
xA5PH7adl7ZV9klPgjHmcws81HWx3vO+GJ2s4/WYh1p6x2HJT6ErdzRJJel0r6PYX8+zpB6dEwob
3tLsQjWP75lAeOdlsxvA64ivsNdKUYjx6rYiS29NSmWGGT07rkVSL672DxxAaRM3Q0nvHpkXvjXl
8ivp3wpSVoRTz/zCpWDVOykd7KLLts0tJFr4qGxk0mqUocLk4XWAniffPpl2eitOLS6VkHSBewSp
CFBklloIi0i/C8RTGyX3UoYD+CkK2I0gLo6hrV1jU/cQBLkHK/sHrcm5rfUyU8K6RyimknI7e+Lg
S1zFWtiS4C4ZtpeIYD7IMBtrTtSOe1VGj6AibF8PmFiq33wPp3nhaXGCDWKkIX9v88dY5Gb9kK8o
tJhKZ4I2Ync6KO+o02nXZsggwquHgJOoG8kfsMW3OPMHqGtBqn0xK/xrvk9+nxgRSBnLQ5onzesj
g0dtsEg86n3x+T78K2X2DX6VnPQ35JQKiOAWXdb7/ifTg8sCbuqyP1JKlBIFc8jHW3Lw92ugm7ib
/J8FRJse7zTvXz+556Oh2i42XLNW/i2UyR54f/SxbEOtTpFNZeJvcH1aeYjVqCgLZh4v2uicJ8Iy
XFZpFiDVs/Qfw+LksYiTfKZ+dDrmWzDo3ImUHuF2fTjjYHFgj5dSiQ0edg44Umn74llwpQq/mW5A
Bs0Bc9Y0yIH4dQnu10qifXjgznBoPqJPWrlgklGpEl3AcXu5Z28G4i3qVzIAUFBIfkPy9swYffdl
LLyKHSD2W5uxDfvC5CQpsUzZr/io4csPENOonj1NZThAyrNmh6Cmkmu7FydGhKkCuaT9fHQoLsa8
7wcaSEt1NL7VxECS3tksIC9fRM2dfpMMeW1lvZQo0HgTt0sSEmEDSF0atoN48P95+HWd6F8Y3hoe
nCiJI84u+6PtVVxZ83lfhTpiHSWR+vkA6PCiAGlkc1/rL+n0YB2qDJLmlWTDeUZghReUqO8aP6ku
O7gRzTcDpHSXGxmGfJgohwH+hbIjkL+nsNjO/QuUVSVQ0qXi5eWF5nciiyKNdDQTx02E72u1UASv
JOb8b9+iv67ysQjg8mBmjqIyqZC9TLJcBq1d3IosGw5C/o1XuMEZ624s71TihIG7/78fuvR5XkqX
wcYxKYGirJUXALu9gMRqiGiXhagv+D5SIuIG1aHJALctWeBJCxGkgwcyRXqj9Tjsaik+WRfl6qLG
Tt2AZBXGFM2k+wratQwUkDWsMW+KoRFimEsQENP/LeRRa0VRparQ+BGTuLD2dsZmzIg/ypybCCiw
QHp2/e479R9Eyv4HSt5AQKNh8VDslQU7EoZGEULjobQ2KR0UhfTchsKJWwViUpoEb/OyNv1SGLQd
21gSurlnxFv0xPt4tdRrwBudGZ47QBqIyt64cyY2mpSaj2lOVhjLGVx+bwBtUo/oyoprGypdSEfS
suj+68NJyrRnCL8I7Eo2SnSCXeOk5M8qx0Y8Mssy39Ny4/aPM5MuxQUunIjlO2nDPMMc8XIDAsEP
MhL1ENwqwlpRXTxsdxvdo99Qi50n2MQhHjsXik9WAi8rJkiJI6qo3nayQ5xlLo+YjbqJk1gH/y75
6BaRNcvULnGDsxBUOIxJQ5ICERaCJm2xRNQpCMKkXb9HplxnNjoc/Q+Wa6zKyglh8vtEH2El0RUt
PrJi6JzqQsRuX5az8/o8yTajm9yQs3eHtMpqcmZeE0o6MtV4H8vNumn6boZkANC6ALkGd5cY0BDK
pOCbZ5Yd4MuD1oWEu0WwXrQwOnufv50j5GoOoHgJ2mRepnYpIIiHg7uQXv2bFic0uRVzfliZw1Ql
B2iV11xgPP1TZ4mohLnpFFVdrnmSjF4VWBmoZKtMWNdGWLE9j/iWgE0sh7TFb9ZMAsfJwPbjNfnh
Cu92ZAzKCsODk/29DvmgyduiNW0HQKof14LaJ7iTGMnnA6ZWM0fR56S50h5W6iMvAbSrBttlxXqJ
jUQKt5HkdbZ8YsNw/qFhPy2x9/JmcRxvRiS7pWyXvA9NGIoKmIqNJXa6JvU+2TNmwRU+vNjVo5LQ
CmKWoJEhCqjtTcbUPrQgIGfS9sA1yftVCqjCRZjKZEjg2fDcmj8uCl3xenxbYqRPZ3RUKQP8AdXC
YlCWRrYIBbSwbh/PcgKUmGAOmgi2tEwEhS2tAmMLFS45iPaASZItBCD0wwX34cHSAAhn1B30GJbg
VuD3vWQOH6kK6cgCpb0mxw+8kBA9HIOa9BDBHVUChkBmvNDpj8kGAMCGD2f1Sbi6vfXl10lLLjeZ
1pxjx3+/dvfl4zRQqrg9ffXKuZvp8COSrxIBjMIaH7LrS/4MySzfuUZ8aaMW6nAn1OigfD/yDUfE
i+boEDBGJc2molBs1r4f1wFyTeegnbkPwH9VZr3cImARHSLzkNtWE5k0eXu6rk8MRiv+ToAHS9Sd
epw5iLRUjEkduNBfxk33G/sR7zN/skClyTjVZsqp+7XLygo4RqlPRnRKTkYDM8aJVDaxDokqTDKs
DIyQ1X0IsQgUzrypANhKkQHrtvmV5ftCbrj6TSuUicQGPGhIHzxU+qUFpKmH6hQR0fXOqzL+ldKd
TL2ERp4JM+B7bKHbEVKjRJDZp0WPDQXz0bgOK6SCuNLEYb2LVXaYP+1GbXhFDYrGAaNA09Ebj8hm
cgiCo9XqHnp2fzSAM8cRCFHJ1H2vzQPXOsFFT5RQC9wGalMXPvZ3QqbOHVQ1DPnqZ7dvl69coE2D
LeZMvqCrFnR4v7TwaMUhlPj6ECkV4rjH4GAW/6EYQTBXF3ZfHTVKMdf07CHonL1dQHDrSIJ9nsLH
iU/qsGoMLJfsd68iTHkITAhx3M+dNO51F2/ydJnSewQMtU8Z+19GPpvfaiww+AdHbgVmnRFKbajY
Fmpf5Sr8EjyrueLF+b7S1CMNbptm5ATADG2hWapAqIgfz6LPUniE568jpIPlwWep2NbH+s1g+s63
KysuSBT/s/ITf0OiQvUuRxFHtrKs1cY74GsB8hqcWYihLLjOYDNokdpQsPu/V4cBiBXDIlriPHm9
xEC+BRSvbXy3VZ0UKLZT3QbhpQZ2Cr/FLIOlh6CMzf6lEanS3oxYBIcuOmwyBpctb1KrU9EmmaDw
8u9DbDvVFfLXrKOPYt1n41LrJU8HH1y070eEUstWyJJQv0JSFU8JnIRmAw1izaDhs6+et+t7tqap
/neEuacnDaTtiKid0ysFJFpU1ueWpOhyL/NorWCrL7EbqYJ6Csum0UVNkT5miVNsjY8HSnnUwNOn
s0zmtzCcOIxq+c7JTUIDmd/+dAgwBNy9wx7rgqBgceA+xg2r6xZI5WHtzo++DJVGVwTp6anLkEDX
7y6pmgLYs3L70JC9Wt07bjMskwoOc4CwH3AMQ8Q1xcTjKOpYwq8ACnkLHaheJbIVZE4JgxclZNl8
lJ/579W8FYknXMAVBhm2DRWrYTM6bsbzl0M9nQMtV+5mcqCVo/GiI3dQX+ocYMCwVfQWzQPrs5T4
yKpNlPiHKJiJ9t9IeMeercHKciAArRxS4jgMw4pl93TOaAqch2ms2Guxz+8tJCivzPPr4hwlv2IB
v5E5v3TVHR8pL9SQatoHJacA1aPmtmnHN0Ak7kIG88qYR7zZUoDnzb8GJ8XXvFzSibXFgM0Yy1Oi
iWq5tpLDORwYzXtjSQXdHHOp+7gQHRLRwqNCR+sqsHY/91waN+0fyVCsIfYwt80Aaj3ZefvUxlHY
3oc8NUSNCKkxSBMUjZ4OmHEJpryt2NbpaLkRm8hXfrsQoVH/9j70ZE+LTLSWx8K+oSpe4Kn16bwg
aQW9lLScj/7svb/5T0RXIP7LwLAIN9BgNza8UYJGKw+nWaniokbMdxVjOLkM8DFGke16irSyQQDR
4FvCp09muyiLjDzqLVxOCXqFweCQ5kqkDboPGmtbwkIRZZDvZy9gjhrcq/GxWPk9p8jpqzNPfbVe
grBfXyjm0Lg2iOfigpRFlL6OGdkMiY/Z2dNmxdeIPJfQTR5tNbziAZ3/Y5rkfjTdi3rRaPCzEfNH
wlVgHfY4MJ/Sn8xlPHbNr1Okss2QVjHfMwy23KpxNx9OMEjPWfrNkSUFwhl9/JOhSQIwlszMKMgw
153REkhKrpK9jQ3+5EDAsKcnkYiL9jTdF9JaleiZaN+OCRkQC0BjPo6EQ4MblbDiIgwMbN1UXNtn
bBKIi7Jxv4ANAjLTdNHqeorZHYvRJpY3v3R5KV0OS3qvO+lyzVeQ4Os8Mlo+HcTf6KD8ANUT+Ya+
WTA5MESXFLtPvrCdGRwHGhQdt3FgzbOJIcSNRlTOs+/T9PsP67QGb53x1p6PnLVF00qc9hbfY/yS
9c+INhjtKyxwN2+rMkBHO4HDeP6AR0BJPJ5DM3y4dUu/xElEgGKuEQf9Z/VHgWDeLa9ZY4lonaf7
Bh2BrdPxGfqHIi0VChC02oTgF1FgaVsrj1gbAWF5RUQtsrvbSRzJkAysnC+f2o8H58x49R69J/By
hDlsqmGztiUtAKgcSAdUVh3oelYjF5wYwVcinUfv5lQvHU/C5LmCarVmut5Wc0+UMgZswPTDtpwn
/aTFquUWgnyp551GRRNU8h2zMmJFKdugNrT+avqU0V/K95mY+5lrVfQsGLv0Kzt3SxrVXqVST3/U
vF+e6CnxhE7aZ54nE5VSl2f5NBUxpyEyQf6vEFW32UEGSvCjIXHv5KWRQWhWjv2LXbDq1L4SSWhV
W4tNjudVVUE2V0VNaBMe8cKPKVkUr1+FDRtEtZABio9L8wi2J1bFmKg537NXKeZKkzTw/B2Y+r7z
NyVMRSBA3nrzFcOvnDhOgLe0+jcASylw95sInE/FkDoKGaK7OW/gXDjNdIIK3qBu6m3wvUJuNGiu
wAzdJP5cAKwUav3ZmVrPbGfk15EEZCGtSArweztGR67RiZNZ4xenndh5cHsqvFgEQ2n/rWGyMbDQ
7Ul09jgkvjHs2YakcLBrDYzVaY4fqEqCpV5lsm5g9RmuARRhdKDoNZW7yQ02b2ChO7NUtX8dgzPd
gCZ7b/8GJSZmxlgg2W/MXUONriIkQ3aT0MY+PlygvCuxUxh63CK0GflH8ubgNRusgwzfsC7JE4cv
Dh46WClw/IjziKRCGlUOlSvNsx+4G/8As+tMYsTU9CCU/itJAjXySXevcEtv6ez/l++Sfrc8KDPw
wout++KW05vXUKtSTfbc0E+MhDnFhgmoJVOfV6kCreGJleeotvl+cn4NuNt8g2XYsbQEXNQSCZ4e
O6M5Ynuo6BHUOcbbJQr3xxK0njiiu7Bw5msdE+yCQrrTRNikMjxx3QqqRnGR39Y18S0m/utuIudA
7r5BbYs0Pdf3kJBm0ZSn8OKDxkPjx3KOdMAgvinKC5hkgPHAHjfBSO/VAF1uhZ+mx/Zvj/AkUNgY
0PFA3S3dHcZxRYwAinEl8G6rK26GciPF49iqeTvhWQbAITBXgozq2HxPTP+hVWIk8YFgGj2BE1Zp
J2K5CR0OdyTQnY7fnGOVZIQlbR+kjpHZURV4JRrkci+EjoJrDgQKRVMZyoWzvRt3gRVBHyThDzzS
Lf2bLQ/V4X2+E4j48tGDnmWHjmvhyzWocrJSGg8VBY4DlNMgi3F61X5CD9dA/RIuUE6p9YHs808I
OdsI+rXK3WreMnB4sHIWt6QZoB5PMnbFGVI3i0irvYEY6NyR/9I71gpxgy2JnCIi+Y8nCp+IIbAg
Bi3ZZVfpX0JOmKZxDzJMuqhLjZ+Bazsq16Xb7SdSLX51PPCXhF+cb+XVOahmxQX/QMj7l8Loz0sB
y8FOFymGym6ecfxdvTGUkuxG2Bvu27ZYCJEG+86u2vbpcfken4DzWyo5gFQ4zbKoCiTkYGz1OlCr
PqEoR+2zGIzOCsTiA4wMdGMf/zyPVLyqJGyRR4wBAqPQe5n6z5LtG6pbYC36SKXKwNE+Hc5Bstvg
HdNntOhO8ru02FBBTwR5PNOf+52GOjqVA+Cm6yY8AkcCpU+Ob/LnGzCK7br6aV9c/7CAckPuRmYO
pmxTcOTiLQV9KsxRnkRkoLPnM/wPbtPxYTjG/4yQ7RPyt+QRPDs/NVIXXBzWEntLQOZFxCfzjcnt
oLiRKEQcJ3itUqNCFH9IhZ3+8LF4L0PmsM+oUZiUqq7sodBWM+kLURYyf1FXpCI2WZN0Dr6JwIUs
K5Y2iqfj0PN0SyO8g5JB+p7j+3v8P69BxLg8hQiwAnmzqw5sLaTV9mIEIyd9zMb+1y2fjs1f/M7B
CEks7Rsm/U2ui4U4qFHG6RC7d+TxzFJA/eLz94lkgPzpxhEPMyawDCtP45VRCfMp5AkTpihLZ/fA
jzoD7SSxePHKmZPh5aOIhvray3Sb3D5RAsoZkUKhewz4AbPnPjV5Bx5k8FFcCfX/bu3w+CNg9j1F
fWUYHPppqZ9Hkc/k79MBSnxQRmoNeBT3LYdtVh88klVQEZdnH5AJnhJj5NjzKqjgsA47FsXm9v5z
mev+NepUl4ZPyGK9iFE/bZ78eDy2THQI7XViUyssGsLv+7PAW3kepMEXiSbx0ph/L97AHz5nBM4C
4znsV7droj4VDNwXwGYZgH/SoucL0JGWw+TcBvW0/KUmGAsTajnh77ZqPXKlX3whZuRCKNvw3MZm
GOLFhWHAmPz2wQyHMLr4WvsnKbHKPYvGR4G9DKZ8AQ7IDbi+/IubwUdEjVrEZAklqg6295ojoWTC
A9atwdPwVdQH9P0COkhkgy6IpgnUn3fJoZs7dEm/IKxecihSG192dhpmOOASSVcJwinP9wW5DD9z
UCAkjLZS+opIdqU5EZnNC26OPjADURtnVU2bgPkj3QDU11AXrBgeaKS4Gnev/xVHlWBj0iH1zXYp
+/UKZtzUTymN/o+3q6KrTQTYDmumk6Q3QzDDky8Ik4NR4YTKvwgJoAGDyaou9izJoUfOO0Lv97Qj
BKFM2rsGrhwTxT7hzEZRgKjbunvHgQqSHFYEQhRG3ZjIQlFzd8QYlL0dYfjKE847pNfv10ZwPxu3
6HbByQyE+proycCgqTD8agVPTUXidOu5uXxtiLkzFYjtC10/iTOadV9dDI1CVXp4s8ha8nwpwVRC
q6vUVv6jF1DVIzNyyx7OMYBKD+zkaFDGTvr5GMYIaFkrbYX0d6XbFKoA5Kat9eKy3ZNSBComb1zv
nHUTqi4rEWfjzBRUjQ94fnbBMziDQwQ5RXqOLoi5LMVHUa62xkIZMyeKhBYR9iru7bzp/FswrWUx
mAsTBK/Pr7XNQqLci9v9YHX5Q8U+hGIHMfZ8VDT6Xvt3rF6X1CkV23Fjdczkres9cJeBlv9qElgk
64QG8XB8bLyetvOgAbSAT/L7s6W7ekbtfI4kx28dRpmMJfK3jSx2LxL+hvTLt4HKuvwlMMPsn/Nv
fBiRs4BeE8+swBsLcx6w3VhcKcf2g2xSWZqybEWgRkoEpWqqdlF36T/fRCG0IQreLdo42ft/zqpy
jrjlijAIXuL95HHuoISxm0kwZCKd8KbYjcrd62raWOjfxFNcqpgIPfn8ADOGeRdkKIV7ciaK4FMP
1RGE3GRQ1JORfnqqGjkih2TiH7Ey7GWJdwf61bYVtDJfi2mQBr/bgysfokbpWDdHi0lJfdpnJGCm
6vJYcKw6YsnCs/yapGWr6V0q8MZRpf4NEaskVmnSN9FWhB1AwT2mOBxaci39cgxYBvm3AHxQXZZY
iEsUrFuf7bg4YXvUcBFIwj0TeCWPpdrO5cV566ad63fXA1lpXq7Hh6yYIYPSXs9Z72nc0EUzTPyS
y6LEpvB+ABJAQ4OQgDAC8bjIhP7tqWtGfPtPdeMd9Cr0oYJa/ODnCWjxYHpSNgN4EZcvkomvsFjg
LPRxpuzcODYHQF0T+9pyk7NAby1jN6OUWiQUwPow4Hzbmn6vOqA9eQ061XILOHGMu93fEW36j2wW
2snVOK4aoDdNo8bYgZ39s+OUt0IzDmD/pwOenF+g+fg13Sl4XripNsSfQvgq61yJVrMkljQZQuXO
6Jd6RcrUICNAwaXBSG4dE8a4NXwLlahgrB5z2V3f9WD2OEpQ1/qoS9axVIWLoIO6KnDszhPRkSwR
VRWsbzLq29Ybbrp2TOzog8DGUqHLGbydxgfFgkTTBZDw8DbcUL331J/8oqyCivxow006wW/Vbkle
boJsORsvxa9XGyH+IjvBAsuuzhaXh2/r/ZJrc2/XZ1LkbvM8X2yjvYLkB80Y6Jf3GgEtLqLs5jsc
eUKLeI8FTeEUdI6EAh5o8sNo9+KF2uViWO3eWuCp7Q3pMybjRb88DuWZ6mhA/T0drwIDpl0PI7XY
81s9fs2cRPRgQLisZgRxYcKD3r3SSfIhggu1U/mCdUZmCSRDBbwm90RMfOd7T1yl4KQ1muMxh5Ow
VLPJs9uiPU3D11rGOBUDUnhyMIrqAAt0AgMTHXF9X6dO0A5nVRhk3ldcyuaN+va13d005xA05v3y
2whGDeENeql0GYGMBfBY4P+jkwX45vP2KVxFujxihpWsSZuv1tanKOOPTHSF40C+qsn8WLShabf3
BENcGuSMhcQwA2KBskqViLOpqzffquNE8m+Rz3G192iWHqM809fy0BjDDFjP8WkcRktoQ1eewJft
7ANFpK+5HIz6xCVhKtWCzTqzqYH3SJToyTsDi7VLwoWuPQ53I5NKSMfK/Ultd+rvA4FY2sOcIlVL
ZlgsdR9I9E7AdAM7v/t6vZ4VY1jmYR+/Nyu/GyibwKsWE/54MRl6DWVCj3YGb2FLlKYYeWBR/9IW
2YYsLb7j1/6K7QYN4LezIEc7WtaPsIQ0X7t4Ht0yd+y+VZa3K2UFW8gRfglfCkRQ1eZjN2ftFDyT
LOqCwWUhVMi7TwTuAVyvJ0nckr8vPV63mbMCfPE+IHIetmKq1DW6MGyuXdWAU0fwE9/PHbk1dc2f
ZLAdGoWRcYGVh57usOKVvmEFMtl3BKedSSyb5dZVpdEe1eHbOMx2/w8zrXP6FhUYBhnU3iPSJ6GS
w/7EsWxxuXFazA7JdfDvsOiiEoMy+jadCA7uAgscxDPzz7/ZunfifZIVZ5sb5T3cuDwhDfMZihUE
DkM1KtzGy92ZDmsgByXXBI4jxRTGfmCrgMBAVSm+FmQDV0wPGvYD667XpOWFzHr+O3zIS6DXdKFC
vda99QFe68Ft3/pslsHSBAMWsu1RD+yLme2eoUamu91qBl0Hnyks3koyMccc0DjeXhfuy4cq/WVs
3Fk0TopdUkDpMfr/13Hu8yGlQm9Ard/+ek1NJBPH+/0CGRb52BUCn19Wq7FWvtXyx/rf4TfHh867
efOrKdb7mRQFNaoOq+S6/VPKkIrwivBQmeXg3OkaFlR10RF+XViSXZVNuzYfaimnx0U8FAeFpWQB
nB/gIkj5RPQ+kgotytbcP0MK6TpFIH7w1avXvM1VbgVkAIdpnCYoF+PgXkL8cA3CYJJkLnp6jJPn
fZjxlUAa7GwovdyA+GETBdTazpXOVP3/vkF2CRLfR4eTOcXaCxbN6btCblyc/SKYutWGDlALeNfx
Ov6VIm9JVvEkQ3Nf2B2IQ2vTilzK7JEx4ztvm3keGMhP4DmlRsXp6FMy0qs3KMkcpqy2ae7e+U9C
jJJGzJxQFYUlxwsVwK+i2AzIi10nJW7NKC3sNDpsPDVSaRnIpdH+/sj8WAvDEJ6Cu9291VeJC7Xk
oCzoQNe0rjv17lnfW2P9rnYNsHFm/uZDsYwUbw7XF1yV6CzBFlnj4RfIydqqJTHf4abBWDeQsViu
YhaAOADh/r6jfr1/u1Sqi/Be2tTLMq2bPZBKTe9BqQziAp7GZJUM3pISrmCChbJMe10VfFnAxHaM
stQze7CDhBl2S0zxVybZF3b2pODl1UvtGd5IZNaLkPvR57fNr30NgeT2pA+EdfCvmLpeDiONO3sD
92ZSpAEY0upGzNP71AAx+AQJPPUjdQjbvgG56xHXjoAo3qMjxe9kqjOSXwl2TS4HjpLioPCI2w6I
8gk26nk0CK1oHGysZch7KA5fBDKykQT0HKZ5m6Kf1Nw+sbeXA3pcAhzWm0ZHXHAavkzRpWAOrr+p
hRjtgrexwT2cH/r3q1jxC+w3whCpImSKUehUUOYY4tjmFrP8/hE+rKVm67wZ8sV1zDr2GPGrM4LW
jFucvPn/AjHHFLxZezs9MtXI+ivyyn/K+FEs1u35jOeFG8+HnMiV8yIBwYCXQM0/iGospnOqGxe9
tvMTuk/If7dS4DS2jmyM8csRE6XYRGC8WvLkAAUO+a2wRMkuEFTOKUHBfxxUM4R4uB32dOfv9UeA
KDzR+CtKRBrPqDS9JtZZEBwevf6oDojHyKVSZQzFV67YLwcRK92WlZJEc5nMULk+QiF7t54zdFpd
8xrjdVE5DmHMI+LJz9DT5dvw0AmXuWrooUqmJV0P+fwS6Xrgh7oradfmdASfaERG6DS/Y1epACZ4
XNFpNvzL8ft8D8480Ing85qVC2e3LjjQZTNwKLTL4yxx3ZIxAqSE0lDlF518QVGppe4hF/CdY1zZ
0u2+szcqcyp/fDk7IoSZUb7uuDUniw/k9iIxvxWDlpwCOaPWzD0tOf1AOQhfyEjMNkMws3gi3ffY
i0hMWazMIGbPHG5xbZ3suLg4DRTSmrR2AHRtUXi3z50Wt3GGlAyAPqa7uGTgCeElUaF72294PCko
qyz0DY8NIcYuzByUW0phKNx0NVUYm0ozSRYFYn1ceLA4zMg4hD1zRQkw4YxwEhzjq9jbvqRiUij4
TxJZ5Lip9RompvFBko62ZfBqD2QWqydSOh3zU1rXQTm4bD4HIm6WkGrF1njKaclYrFDw4VcuqYsb
/ItWUK5UuLhOj8bQSN59IY2nFTcYw7KQjwtFJRqMizgUQd51ckMp3UIk0hlstcymZ2Eq7mMwQBC9
lpBNh5KddxUSnD6H51oR41132FCZqBI93Bg5gsysncjPyrrvalQOBQoXh03nn6gsXEQZjkSRuJdn
u2ltRUXTaNhty9ikd1kDLVH949YwRD+VFDAD2suceaC8RC78Ygeb7LAq0svbPTTzYscJRcxNjHpl
bk+fHGglIKMbiGSohWDl6hLlKczVqdB8asp9j9Ljk/W6jAK41UA6aohP3/QQRB9d7ids35QFsxta
MTVNMYW2x1YmV+Ln0J4FL7csKnbaLlOF+7w1iY/Au632lqhSNmr5AmdC4B+ZxExIVSzex+x+Pa/I
QmSpskTDNGlMfh+zCGnfFAkq65G5oa6hawVrZy6YK6XPbl4FvadDKg2zfq2hoFMj7sMOTTbTBNiK
krBR3RrevSrwYNdPbHpHSKQDl9wcopaFvN24dVuum8ScJpzYHxLB7zwuLSLxm4bOZvQcd2kye3fV
dqA3Zch1v/Qq44g4Y2lJtEJuv2lQHFlqHrMYvtJ/FSoqZsKyJnt9+43M4Yy6WWdjdIrQY0lYI+Ge
QkYq/F0NeMVnCuMByWx097VEAplaFA2o0Ajcgvg7uVd12TfAIN4zgWv44TR52dW1pOY7teD0CEnp
PKsjopczQBcXJGqaLOUHwwpTBKBvmJdlP8CYwDm/QqR3FVJjvgS7SfZa8TJHAp69qZVMNNI2YDbW
E+B/s3igN3Z1r6z+vjwWCXQyES8SF8Mid26EsqR2TtUOQm8MDhIQb19iNuw1Y/3FVEA/vxwvFU+n
w1RLNRyZYoYRIyL/kUrTBQ2UygDq5l56jSbUhOLqEbAKXV3pIFFEOxazxzdEO+MeA1pZgBKjoM2Z
2DKF+Hj35lpiKeQwcZsK6GVesS71ifAWHh9U6tcMqooybS1hHwatF0m7VJuAWpy40YlYBzayXyV5
WKM63Jgm6Slk4aoBY5dD1AH+8B3RJwMi1oNYiiRzyRhzdZut1m5FIlJd9oJdJnhNh8KRtjw17qBV
esgRHiUU9n0q6/lwxFpxbkmu8/IYh20OTwji0myHBqNORdioaznd/XHlIsuLUFzvdROeClphlEK/
QTAKKOTNeFXI8yGzm/d8PwmBZ/ItjqpmLUkkStZYrVlKOiNWPzNCqBuykiq8jOMUmDdyYuMxrcu2
FpFH08DVeroGTSsc3ZwUQKpFOjWWZu9pzLctEMfH8dpqX5YpL1IymbHilpvj3SXQyDF5rqL3dRPp
x4Y7/gtaV5efrVt8fbYa7tma7P+rSCLvDjHyGivuoXUC6tRaPNnzx4VgJTYr/aT2Mm9PhB1AIwny
SMVDUU0A3pgJ9aSZddHfrrvdu9vqU11Y70KQpQio++JDFVGs2RPKC/lcv3lyoNtpmYZbrXCzQc5q
CPJcHn3pKAdcB5klEhSIeZWezoGiyEY9ZS92Z6F0Jg5XXapdXELYuoUiii/fPmu8Xqx+ikEvQgcW
htNSaUWJtVdJDDrPsxmxLC0G4iz2dIWgXL9f4lTNQZoL9WP+QKrIPdYTkXNZu6qyzDvlkv9q3esd
vYU1bx48lcfy72oSwVSu5d+8sUseivTWJHjYnHIoWwHfgqJxRf1qmzTsS/mjgD2digdw4CUniJJZ
c5FqIobPCQHr0lQ6hGu8FnHaT68o5iBQ5erfXhogk//BTyf1D/94Y7eLbCgVeHCeo4Y51MVFhyhN
DtEXFAr6oyok12JFfYMdRNDcuHz1AQ5xMe1xcLY/2UuEi4g2MPhIguWoiDlCO5UIYQTgEJ49mBFP
hjdlWZssFn6ArcuI72eniRr7L45j5crt32CynLPBDE4c64u3tVDtnlxKGNXK/Gzq7s/frsXYL63e
FBXk3P5z8OuQRSay8LFG4P5o7ImjMAdS0w/unZuxgZHRthcL7rX3SMvOscCExwLLWb3gd/LAs2+2
avIsT3dzARnJj1KMkJupW0tltkUjO8J4HLOvu9zxG3sWSzEEQb1EDZcNMyik0f/PfvGcn/iMe0pT
+nhtWJxldf/eZaix1ljXAUwlOP8bOFmmglS79B8ojy+qBtsRemgd2wPs1FztXYGTDclgW4R1/ENA
pqb15TQP74Es2qYAizc945LSuMQV+Zt9hxYo5huNcpIhaSewd670fR4whAMAzn2IZlE5xrLscQ3C
+rhJNqRlaaMmz6fH1a59uUV6KeqsmfpKAyb0ZemVA8C/KC2it7yGVvqNIhY4/xW13uyWhhixRRlT
DQClv6sh0FtrnJ189SQGS4EUaecKYqYXnOXHoNnsjntxyPymzFRN6gNhuccPVZln349/YVVgqUl0
0U6pZtS3STiYTQbEfunbL9Hcmn7IPIItht1mIVLyEIsT9WBpqcinKdzGEFVEpEP3P2DwJ4/Txj8C
DZp6n8oHHuvlDbE/POE0Z2K0XiB1S8lsqKrNL53F+z9eIYaiF38hyH7sdwc0Pqe4629D49ZZJ/In
D8MejpwtLllVMnYoFgYxoDwtKV5Ie97DF83QFxkHTCK6Hs/SUm+lTlYgGroHKj2WW44dFdA7/gbx
PtCt5DD4Fy/tDKnqVwbRDSgTWka9fsFKNKd8W/jSPqts/tUxA+ZXnDAZVYP1xEaRH/AZZDLSo4DS
1sxGsKht3jfIjPFQIpKIj2vva1pWqvYEcVJOShYpk/Z9i8hq74bWQPeA4FO3KzOPyGfRitJzqo0v
EXOwRf83fo6D+IQwja/hSBdj9Dpdaxs9V+u+SP9baW5gmK1i7WhFmQZ6bd0J5s0k7BskJu/PEqrq
BRUcx3njgB4roKfyjKgbqL3kmj/GKVDhcXoEPbivN8XPMbMwzT2FjIiYfLa0vKS5vfyzQTcI840X
RFUjirDbzlChM0bFsA5HuV+/ignOGbtp6a/MEf8u+1VWoKHyFm41TO2U00FqMbECFzQD8v55hkhn
u7+giOpFdvPqTNl70S+zzgB2GS/JbBTD7eBPVvImaUOC4+Yb0rfoSPqIjMC6fNhK4mv9p8Mf878d
LHcui0hX8C9NWq+lfqND4IZW5uQwztJ0S2sVRaGXvqAL2G48tvehPbLzpv22qZRekw0sekYWOB1A
7vJR6rx464uTHScgoE5MlE94C+8pSO4qEjttd8pZeVGUwljhQ32/UF+/HatbHEwOApgUNjoDYBD3
yzmVaQmZSlV9f0AzfzYGmDhg4m5XBUzmNSvKnJ6ZKTRnObawOPcfLkIPKFJ9qT12ps8h+0mFtgk/
ohD/+z8P7MOBrL3qCrrrKmcg6WYnDA7YczajASCJT+I6DEVZ6K6EixSu1mqSS0iwvCGjEKs8cRey
69EUEwbtSxCiXiIHsxVksMRdV+H1OHHuKcMpnKXgfX/LpLa8DM6vqGggkMQD2vwWCJJaUltEL3dj
PO/gLidzDkChuRbriqfhLDioJbit9R/RP2pXa0UqUWDzop4h6KeYvFd1ig9amt/slCZzxAVZEZzY
ONlIXgkle+mqc/IllffKHL6DHDgMsSO08rYqjlhJJazVDXAcRxyltSFEydG2kL8iRQvxWlcoswIP
pdaVYXJ1z7T1jVirm268sni8Y1nIL7ueeD8C8pYxz6hqDRC56GDLkM4SAJAPP2eF9qMvi4vP+nyv
c8eVVqvtFaygkjYYK+XUxDDBb8QbEChMf//v2+xScV81Bq7U/10vZlAh4ttjRcJrZfIywTCt09O8
/J/kWIQJ8GhFRh+oMMGj7+8tHq+BV4TGtmcl7Sr4q/aYoySdJSTJQGFCOUl8Gy1I6DHuR7YGgNmt
lJsJnflPaNHvlGihBTLom+SZXj/Z/e7G4LZk5vq1CK5Xi4T1yJTN6d8vRUjCxuvWYnJj9ENBBWkp
JuC+cqT3Akz4x4JcPYeOsbsGKc8qGY5ug9Pbnja3uY1P8/7u1YYfbijQbZIF1Vt0zcsBSMelU3MW
FMzfmA5WZD3RmQ+xSHDVh+scD78yqnbDXPEW2NSRVIEktG7+RZoVqp77VLUmAP9aHV8o49wkQ/Nl
/+FRxYpkiFu1GAcKq982PR5LXlfk3SqIXoiICq9oLRVU7Wiu1USYRA2oO69G3vWkzdhysoeJuy+i
AlBmAfS7ozZBJkFY87M2Ubn2e91ZccAjkJd/LIsu7ItMG/huS/8d2HAwMdgXhVfsZDdlF3aQf7EO
ofd86wmwhgbfhbQY7SA2KaTxMb1sLLMT78EYEQ2dJjaXe6cGB77LowrIYZskLavA7rYqH1xBEPKT
5JHszYZM5wnsHZxs/McWrKh92DD9L93/SW7aWNbwkGF9YwXbAf0Wz0jcZJ6eUTP0OC+XNs3SmWKj
3PpAG5rTrCmvGWbrbFeKbr25f011JcjAOSj021662ttlYzQSyqKGGCpHTrq1KsyFW1y+RCbrnk+f
K6/qcto996fuRfa1Ri7ZVJVgxol6sw1VtU5fzajyyJp4oNaUmDUFJr5KvwyOMiow1sfG6wTFcBwP
zZRKXUgCFNitktT/Rm2xHrwBMEPcJOaOFxKa9ghPTsQzgHtT5tggJLRo6IqLk6aZmlkuMjJ8b7ti
+uTVK47fDk/ulAFyXGWtVZ4p9+0s318UCcGv0WH9SWpxhAaslFI17b42vtrirKNxT7a20YaYzwtg
BWWxmDVYSweR+M5/ylsWEFSCKdiJdvagr/wRjPy5Yi+X18T00q9UGT49jKX7x2A2xO3wN4CbDt4+
VuEGr2pdHzaHg4Pnvjp2WZjRDodR7ZghK2Lbedcm5ltvI2Pb76KKDpqdlh6nscyLRcyBiUkwiSFg
LqFEusRHA5J2AukVJE5m9zDU2QLVey+JYBCvGZvyNsW9E8kRCFlvcVWfeSdRvTkKYcYN3FNsn50x
nLLY1nfCV7IRLjnzrWYgaCAjUALVLO3ePAyMxSqV5tao9WTBmW6BuaeI1lJR66VlDxP8WSc/LDM3
sqVz7AM/LaPj5PYiGhAVEoq6pggW3kSU516w/7VbtvcDLFuHe1s4ggdbyjN2agOiXjLL4mz4F+2Q
UZzspAk/FfmFNEIzXOBrnFy1MAo9rzjE3eTqtVVJSSvEbo7iI/vw8BkR9u+nyNXF3b6yIWbpQJz1
6ueFYZGMsTVSdTPAz/xbHc/nRcv8Fmj/OTyuZY8Mv/GVX57jVI+e9PX/3lvTFWG/OzjLjZLM5+Fg
drC10KvWzpwZ3U1uuu+bWzB1SJrfZqCYpzynZRj3FsoxXc40UoZ2aWxSZq4cFbykLXlMNGBsy/bJ
qbqCB0DMTXlssCsgvhhN4dsGfXOcSQK3+BEfG4NSqJnPNYPCp3XiUcPZ5IzzNhvNXYLIBlBXUV4M
LfYPpFVJH3TgPcTARJt60ibvYgz2D38yBEFSYK6Fuc/85qyssxVUMY6wddTVLyDMb2fxxi99uXC/
DDd5bSeGFzFG1ocu/s9kimabMhQ6OdAX3pxy0npkt5+Rg+k2RpqjMTy8VNR0CvlrGbeMC44hrzcL
zG2VdLuaNMTm/WdCYpBRR6awJ0j/+kHuxblZarPVw22BaDMI1Sk2t0WI443c59QlKyPuTIociT2z
8xoIhq025V2pbFb15PkEWHi2fu37326ps8NBPjIZ22LAzyIe84BQPG5im+VIxms9zEtppPWlb+SV
IsJ1QrYHIljOdZIeLGAHGqoGvHOD15eLl8OlUb0brkn0LGYFu9a7vs/HHD7BUVZN6+4R5YmyK4sH
UJodrntcZTPqClTiV/C1wGuVkqvSmXTqIMP6oFalgkP/+bYyo3rU3DSjlPP+rCYNZrCk5mKjqygZ
nmhEuwnLJ1nEjWtfAMd0UIAZup+sKuRqSoQchPsOIje+oMrVX93xzIvJASP/LQ6JjX+a7TfYmG4R
L+HQd+HYolf1HhDlW8SE2et7VcncnKA+jbnh9JTmpSxjC9M7+RkW7gwN3/6FFLsqT6o26pKGGbdK
VWFXn3mXyThJRL5dZUWL3gwKzrYBP/C/Jj+IsIQEqlvb+Jv3O3CjXMv/kIDO2wVRZb+U9fFYZ8Uy
2ZbX7QQaC8dI49GzG0xT/gASXlLmRdeS66A6wIcE+01fNiTDDYNIxuuiZbVVEt54LHm5H5BcNIgo
sdWeQpY892YtM3sr+PGSTc1ofkQSgOV+uHqqugk8JYV5igZ1+RWsIByJ7IGZGsykRIHKabsC8L1f
E6YuGvDOqzdVu7z6ICL/HuzZ35H2r5mYdC1UVbdnDi2Ub2lS1eg56ykmzW5AUKLfc3bDyQesLvTc
JJaLSddQ094HjIEXMXy/RxwyL0R7XTHKp1eQMZS6l2H3mV6mPF3P7Mq9LyqpZR1zTXXpdMynjP3F
IiZ9oQHWbRg6WY9Q2cM8Px4rbNu3ffMVD75QqjSoE5SlFc02V1mQHks3AfYB2f5EexWLfTtYxirs
Y7YrQEAjzQ3iUOyebrwWpua1/0DWej0tS4VeYSpbaNRP+JMY/s6F2WCFPbOc2z01qXuPWnH1YPtS
sbCnoE5MhQhgNqokneJWRZOS5+Tpnq+sUWQ2yI1noAFw65Wqtf5MzEdSb2RehkqvCJun3TPjM8ee
YygtQ3jndhNTd63Jd0QFSJzatYn8VmXIM4ZyhFAercGF4jg057Y/YRhQES2Jz0pBuS+LWwACw5Sf
a1kSdAgPVxFcLkEgpYZJhk7x1tC7TknIGnZdpKZ0xvn0aG9KC+uncMi1qGe+OLyABo2Dam0Oz7gq
h01bvai5j5mTuYz8udRs6NAvCsszUCMAxwVv+TVs+Z+VgFYRYMRJ83ohQQTEVDG2WmLi3TiVYOwD
2I4Wb3JcQGD2gSLxQafbq5Bu2Y7Qij8cxc04MVddQJARvAnuXJsF0wpDwAI0q6o66cLuVBy0DYU4
UDsgdXTd53pw2yv8k3uIQxplqf6nJfDUS3xDJM8T+W+SSxpapz7UrsBCxjBhtx+FKvMM6d0zaL7R
mOMyNRluvNhv4552fJZP2iKIW8fLnGNNrKbZ46om8SZwtuppnvX6CvjkdnfyKrOlvxMZ27PH8mkk
PIJDFXljqCcZIM1DiS1bh7AL8ph7jMpUa9+BhKmZ7YCjFPpyyhWVWiHwPR9cm7dHM8LwExTaZpuR
nTYgFhIbkTfCzvh2U3dOOj/bSVcX3kjqJTFRQIxbIwwhH2xDDDecWsns/ZzS84FECm1fq5+5nRt+
FmziVnOt+rJs2+iu9YhaEDsyWoQjv31lsTEn6gqpSFNTxdOvDVw0JiGCfMR268+xm2JYNWCbZIi8
j8w6TPLzFnhjJIHx/beSrFBxQ92Gnqx0U2V9gHcT3yKFKkQu9U6VVDCkNX5kU5AdLG0jFuns26Y1
yfGS2VCsOUkSx0UaZKxJrIiZ9nOGzW5XIKciHlCAsRjv8Te59Zy8pQ8n2Hq04BtFXCeGcI7VpKzY
WCXhtzZ6QZrxQWNH3cUAbM/+bctTQRRxQXnCGbEISqWpVBUWPcTEJGChP7I+UZuLLkm3hxtMwc6b
ehEZzGh4CR8VpRLyGBWKon4SF3wP9spWn9FDjwR5F9SSfTutPfyvxjdIvnMaVCpHd0iDmyi6XhSt
vsaUp6nopCVM4wjjJMaw+Fvd5lSwdTDD8z/jE7X8r1GAtoVWTYsCQMF2u5SKKkXDl0wgf339jrfp
xtFwXMU3rqZCqNgccO2BRW9bDuFXKAONI2p16jsPzelDhUpoXF6T9agZY7rNU5mfCkMLsvAXIcxg
qMKslQQDob9x48EJsOS3fnC4yPiyvBEEBMottm4ITPaJvli3+lc50aMX8jiAHR6VA/vSdn2GsPDS
1G1ttgWlSWhvjGxssuKU/SpRHVmTg6PSDZ16P6vLbKg1XRVK+Q5zLETHaaZIK8g3ho3t6FwJJL8j
GhQox/n56axBqS+aR/tmDwLgbq8jlMyigcx3AR08aroBj9S9T1qwo0KhIXA2aEn4YlU4V9/z8p6h
kzYgutFmvjibMneQz8orBL7bPHmh7WUWXIKvBOzI+LWr9Qpx6SiEIekMd2mfrNL15qdsaOgwdYTI
7ou8gsVroRNkvWejSS7PL0kmup1T3mjRMbtHnl9w4MTzP2iujVYSdFGSp6d+sBm4tj+WsXj+Dari
kZaBQyPHJ0HxAdYdhF7DeyHP1NT5cFkSmcoBb9/L6SwmXfug4r8GMwNif92CW79UFPVuuT0VOjG3
Qa0i8BWlqAD0zKOui+5mXpcQIvwJU9gB/tT7SpVWWRJiUviWElVhiNo4nWswKG9CdSLqxl4i6gVH
rrousHxzk4FVZkWfjMBAgUujILDNR38UJciHZKAIsK+81OjM8tpq96DecxqD5s3+vF35e7UQ6Irf
VwDiPyH4n0xzINvoRuGuP2LoUqBYJojSCKgaoBDrEatbn5eNfjGJCqXJ++ttrpOAitnzEfEYw032
auAVK6BaUjyfMdECFnLx/6+p8hbfVcAa0hQwGRDi3wo1PxXlVi2N/V2xWUpsIAfjQPVs6ZR8wxOE
vpTnn2V+OhHhuMJiYMDcJ2G5AxWb+jEGcza7lGDHQgVZNzXKXI2OZaa+apZCjn6WEztDxawirdtW
1ifY3eTSfM7+LjnM0wBDPEHnqaT1DRlgGFBYK2hGAk9QAjZ4z9+nIaKyrPjlMYypZy+EIdQuqJmd
OFyP84EfjFYLy2gHI5JJRWWEonoVC/cbA99kvnwHCN5Z6eMtk4riVR2IYMRQ+YxULqi8y0xzUzPe
uuOTZF5iaW57avlsxdeRyKDVkDLSNKs/DMxuu6Pas+o0zsRPHg2FJty5erPAjbErZocx+E/1ZDHV
Rf/icXIsVJxzBm4dhhGy2a3iJo9kuNKUn+tolp1eyw7oxgPA4wEH8ZYP1KSnnV9yG8q/2FOmY818
yvLcVEgiV+fGjjzDyTvGfSyzjJjRjhQ9TL0EB70Fd++bPQXALtTYBipAvUZE1Ba7juMruMUXh1Fg
pHoL3S6IYeaQRsA1Fyky+K8oslHD3kTCznw7dFi6dJrGze9di4b6u0c+r/3OCBmiuFuVI+3gCvok
USRLBp3F0bi/u/6+5nXO9K0GXlotkONvas/+ICEBUHaRzOaGEEtOCLcZ3nAIzaCidAzk/NyrWsfs
guMj05jPWjFipIC5wF0VCRUA83jUq6Z7jIbUXnpmcQOLctLa/tUBXCeR6Q1pV+KPuA4y/xyLgNqO
wemMLcfnalUY4b87/L9NdjlM6JZdUASvqZAEg/P/SLPRWDvk6du2a1XR9TPBos25YQr+l0CTR80g
CP4Iej9oD71mbYWzWCPhRWY4p6Xc90AE5jTq3RQI/xQWFKoANswGF8SZywbc1A9936dzv+kpJ3as
JhBAAMTl6lnc8UEllCOJO0BgnZo1hdhI/LgYdSxG1JR0/FSLIoy5mu+Sew2nn/hiVNAF/oeo0/fm
w/4El0l+3vG6uBLbiAP2cpEEtvJuWs0iXdF75SdKzs4O1vgQknC6yVE/whabyKtGoH/3XY1nqGsJ
5gY7ZVVJNcmpdh2Bsb9k7/l+Ug6kF4FvUELPmqbPU/RCpIvxu54OPZw0JUY3pNQwDujzlxVslOKp
P/GWipNFErAIjl2njidvhyzuUklRkbPef/ca0+4yK6q7vG1k+ErP3bnHgy8uRCXZYNCYgebx7r+m
i3lVEkVAM64P7cPm7/kRU57Wla3BKHf9xBeWK0veFW5rCwnZKBRQMhR30MsP2neFpJmaXLnBvNrV
nvHOyxDDtgpev5zkZTES/5OxirdZMjnMuYebNoDN9CXvyyOQEJSbf2jIcQBokPXW04euhZdlRQno
64Pq9iBv8WttQ0KbpiuhXSjnV7obVBo4JzTAwbNCPOI9ooVPWsrwMZ2YGcs7/DaCUFUJ4dIaES2s
wvgDBjzDPNo94TRGh8uUuufLJ+1CuawmnteDVnyRtIU1owEh/7l5Ig6jnUTRMR+IzwBzrFmgigBo
QtMGVIW5ZkO+bgIZUlACalMgwu7AfM4l7LDVSlwuyVmp2RWPJxF5nkN2NjACArplxxDavptOE1sC
CD+WwShXujc9skqeOtlX6O5l5e00dS748uQwu0Z8NQnTt67C+pYVqbfYrvi+kuYendWTGiT4kEjE
ahLRS0sjOIZ/b2FcxM2HE2VOtiijOiN1rbA51Mv4S2EjR0iqFli3wTetI+so59X4OmbzGIINGkvi
DXZKqQZeB9RuUJjLiMOACu1pVhQQUVSUoOp4Bhwi0AAJQz1i81DaOnG8ATxjf+rX1DSFMNlDlcOe
xPdOeC92AMmCCZKMApr7dWvQz3OuGwzxBiBEQJO720WBc1pJp60i3EjSuMOSKNCx17W6gptF7w8Z
/omylRVoPAFNRt36b/1KaC4VU7gwhhRNQZPYMYGL89yhr+iDUqsDpT5bvu7d8OWfwVgCS5iWNCce
wO4POBIORz7dUW/PlKE1fO17sG0UQlLFVU7srhrgOWw4Tnxnf0C5wLJZqeR6UCS2VyC4x8MdLBnn
fGEOx1bTlfBvYM2C//3GQk8Bo3xDJXf8DKHL1D6Qpl0EhY7/DXkgRcCS4OeM1dMmJR3wLuSESpiP
qu0RK38CRSxyLIY0b6O40VW7nYFzZEgj2asTQUWrBgoCd0q4z4kLeTaUp/mFVp4YkbLby73FWoh6
sYOgTTs+pxKFB+xc8XpOnABS7xjy0UPHdQSTnh4yEwJaPqjd/JrIrTN23wfoXGRknCAltEk6MU/k
pzPceFSsLuPp7WruizlayPqhvTP6KOPMHGyf1uuWTQuT81RTAJI4icDnRTJEt01wbiRELL2syfcl
8HxXRXnNXJT60zGAHkqFOLpO6k+7egdhwdTCTB84IGw5bJQo+ihwzu1wmnbGF0lKwoMSw/ECTX64
KXpbphd3SYen/0VervZYpe76ZpwoK3b4MW9Q7ixo3YtFGZO5PNgpD8VNenDzjP9JnWuH8PrSkA9T
jV3+w7BbwpFZ+ov6O+5Ey/fOw+2C+qbe/4a2LRLD9N6Zcy5RvwVwwworzmUqtp3h7iyqGkDHnc2p
b5IPJTtNup3tdQpiFhfcu9HJ39LmCmvWTuGEURXXd1tQVJHVE24+rKEtkXeqQEz33+I8OSLnlYcM
boRH/CBVpvGQRRajRg7AdbYdwHQlgw0Mas9hCAz5YGvEgXufoYNJHrCLPjMRRPYTykw+ghGMfUPV
+CzF7v1Tx04g0rM7eFvK8TWmQg63Ub2yNva6g/MNiXtU2JbviRxuRaRy1Wwfa3lRW8GB7jaYIQeO
lF3XcGYPPxFP0loY5ItUazOrpwwOutlhhr4HXzjSIEBkvNlx2PZ0ULAaZKyAcXMXXgbilmx6dRFW
qmUi7W/REDNzWoUsUaLuHpydhCPqvda7Ijs4XpCCxMh/jF3drRk5dCoPEJfw4oxdM2a2Wp3EUkj2
fM7/oEHaSuD82Zk/kuB9jLeJfLBH1qwWmAuctUnJrCuyABlqZPNiR9nsU0TNAkAJHSReIJ+L1s4q
iJS7tYxUDUHtrzzKOSRhwDrGAtZZxjVOPJ2fTvPijMpVtgvrc9M4fPPtGXO7bfQsloch5BMR4lwl
yFGmr1IvX2CJ4OP9tA2wfcYltvAVm2J3sdd+L8MbDuZwinypR2YDoXX6acXg6t7Rkc7L56AI82mS
TKINYjgRYdK2IC/mwCE3XtYeu1pq0WVI5d+KEN0QinSGMcN5gxqihGpSepHZKu3jsVfRNTZi50+e
U2Jqmgl9sl+IP9bHhDxcUbA9uPpdP+hZj6EJEzFRAOmT/mkNGUlVVGQYo9KG6yDjgxsipfwY/Hn/
PXwWOQzCDAfLrQPKmAeEAv6dY3k2z99Epw4V7gdwyh33/wQH9pXMA5GxojarVPSbvFlSHzY2ghXa
CuE10AfU1Zx6lv2Z5eBNHXhBRF/gUWHyUG9Vw4+E2EchduR77GW9QCazFNmU/ILzA4w7rYh+sIro
EjN95sZZMeUBggRKtY8Ud6tTYbFWxyRcFnhAJSd+pkHzOzqSQdDkPk3cpNd78leJtcezReQWRQe4
gWf5DE1pFWXnl/AmKh/iVSw1XDh91A2MrJ2EyUH/anuRDvdWE4tNU5a9Y7aFvdE838dfp6jxoTSX
CZwuTpWk7TziMO/MC7o2GhkNmpdFwvDNBhLtz7UR6x8RXpKL29KysJHL53mbpNXfIEwbRgaw/Hci
ZAZmhaXvlaPllVBpX9iVSqan9QXi2Bs8zTMjxInVhcolBbxQIA0Gh1pIxkT1cOTweMmmqLtczUDf
hOfmGP07PXynQapbZxFUaKGSMltURuEkKUlRHyzf4CDZbMo/YLLKXC2nAUiC8bqlVHlH1Qz3nyLE
h+mGiDiQ4f4rYAzUvoH+WV8vbZ50zKOw+sAwecj+D1194FMBZowEWcpbpSnti8jvVp5EBXhQlIaF
em2JvQ3j9d6QCXrX4UIIV/2fPt0tRi74+k77vbGxACmZ4WgOFQl6GAEtw8HrYJLo53earp9qd6nA
42FOCdK3K0edFxWoiZJNJJPKS1f2TaDc5eUvTNsoIXL0jVf7emZH8REpSQgSJoQXK3DrEynaG/iA
5G03RZPWI7eAz0FPDhn/PbFbeCw5f+RaArMi0p73ewA3N3VZFlQNfl649M7zABaDGLqmFu0xVzzV
+UOTG3v3EfS//CzkQC8MfDk/dcsv5Tk5pifB4FzGlR7dJOnO94iIHF1ABCEODv17COPnE7lois9W
VKlgXM+Jjfss7wSp81vUxCmEhp3tHlzZ2X5oqWIoC7hWIyLg6SNyX1pGswl5QuXQtMZwupyVnMh0
P8JzfqwiZbPVMKwyit5RruLiIo8mQinqoKwv0W9qNZCJ04BF3G3dbDbrV+LAB8ow9qqQG4FwaVkC
5Xb5eXwGJziO1qvnScqDYIKodMy86XD47dYqUwwOpnbY8sgXKfk8vci1t5wRqi4ixv63Xojgx2uC
uFG82NGOB7u1WV7UuQVUBEWx560G7fYuXvZMLq6iR+VAIW5uLJJmI8EU7G6B+lJpuNQTk1gHYujR
1IHHOqOiY0zK24tVOx+icZcPHe2jmps0Xyn5/OUan5qxtsfSOtNzdue6suVp/md1GxjjOuT32vEa
FnFBMySF+eASs+fyrFwyJf7fe5QmOUHCahbaAe8FopwuajW0x7AYr4TLLxYtnGFqU/uGYhA3WujO
xO/xzVnrDD0uURfvVHKstWlxO5caI2i9vPjQLwgUfH6LpuaNSXF1mhvasK1mbE+QMlkTz8cwyysH
zi6+Z4KwrHJVE/1KhdV+vxoHkWrhtIpYrRRbeo59yPan7VbohrgnjNQrACIybRBWKIJpg7pd/L4n
3tRvWKAfeFoNEJAfGbinAzD74o8y1gjZu3r2GMatJ66n2PB395Oeh+BGwHFdGNDiGftvw9gcS5F7
14nQ6PSyyDx0n8vO2MPu0UoNTINLUvGcRi0Qse0a+ibZernPyNEwhkWtWx9ZiUrYT4XXq/wANnIk
4EuGyQmn/93X3B7FE0usy2Vsw15Qc4ZK02CDc+lQYxRailDBZdN5EfCrvMho4xsVfUsVczqcnEjd
ZrL64jHnfz2cVCSFvzWbXCSkYCYO97Upn1mRkOBBklWM27ZORPvCaRKDjNq99zDwsMG4cm8VeMs+
SZ993V451pRyEiIGWhWxIUbsMv2AL9x9yE9rnX1S70gA7qoVtWsi9HfT0qsTMMm1g/G2zcrIBkdZ
5TrM8cf02KZ7QjXMdZOwui1rJJM6qbbbhq+HFK3e+tqytobs03REfmAIC9YDeZ1cW7yNSseOZdVB
yS3UlXG8mZyrHBbM9EUPECreJ2lvQogEIl3nmtC5eI2rTCn4ed1ibVE2rJrAjbBLQAiWgXck3gSv
rUKKfB0tYH427DYQOHDMXlbcOYmpy4tXWTOWZnVbmaekJivAzWgKOcyTj8yaWyOKh42Ow5Krsnh9
49OMgK1lvcx8Ft7v2V5BVJtavHG91wI3zpQDPqRhavlB5u6+p0f3rvaq06LIL4kLxPaubP8x5CXf
3G8blREoCwE5T9YdAM6TWAywPB9om8jY07n9yslDCW4S1P4w84zv5LsZKnmSiEmcOa26kHgF3Nhh
6nqFBSnk/llusVhOFNTbyJJRfhlotKQL+PcyuUCpBOzukQQ4xQ6+etFAMO8xwxcwmdyNS33GzsLz
pjsfGnX7V6AYKkvCnEQhx8c9K78bziUdB93dIR3zWfiTQ/fMMlUHR4MibCqS7FZ1wb3ghLpRe7zG
1B/Y9mJzV6G8IMZjC2yd5umrtIHNFctyInF9lNdpt0JiPozwhmTo8YiWGmdEh6UP/EZaQhCK2OvY
ocpGMQ6uOhvr+XrYc5ylM7GPhR2Hm7TRKaeLioijmwKD3GuQM9JpaoCsrwwzpYjehTvE30QYxJw5
wfDbe5BWASk0KInSfNgZFj8HYb9o8jln7Y9AgTzW+Zge22n1rZzw4ybb2d5Qo88sMRRk+AhDfmt7
ageypvBsJo7lNdOPm8Njnl2rAIvgSt5t56rUPIpNsUjPgfH+evJzMtlPfVVyXkho0ifi2Ga7qttC
Q/dylTaP9TkKA2VfiBOpd9e4BM1h7h0HCZ3e9FdzXbuD5+aTI/tSKWXgiLQ6/5x0GqHHlpBfNszR
KPhqXVtuUaONcr4cfi6VdiheoVCj0xRRglnmSxBu/EFlwgY8H9a7H8Gd1uUkHlLE3A4NKZxuXWI1
V/rgzUh8REjXX0oZYYg0XHlkZ4+mBU1MCHinlRWP+0U8SYqckxMHtgbHmOqmU/HY2VREFSGtW3ID
gmYdIJwT5i2SpubtoFRTJID9z5iOKY432nhRkP2hrkGLDK9m2U9Tu2pFWawrFd8F/2H8XDrr3b18
3YpGbIn6oQ82D5shDxPCkHzxhEINAX8zwERFz4honaLWMiGl8NXP5iBsNC+/4+EX8EcsXT7dLelf
pd1c9Wu3QuHMlydh1/r5cHVdwtGBB4z+mbLDEUAzic12x83spF/n1eRo0AN1F/Oq/hlSjxwfkK2p
R8NwItiNWAIMe+xVGI99pNXap7oLkulylNxKzIx9EfnTxyvXaCDm1zQAIkMGnZ0dxq2FPcxK4ELc
p5rF6FluJ3Fqo432UJ1mxNmPiR350XOvxswbgDgI13YMCNkSIYBCcTvigJy+0hgX2qkZxecROGXq
tAGWaX5AHdgM+6LGeBHmQiMJZtr0pbuQKkD27mO6XhjIi/RD21dML7u5exJ23A+EZzbirJ3oOkv7
Z0oI9hoUMDhPGqDeyF1RYkqNbOZGuh6Du3ZCOXjakVIyr7mObcCoP0JxULaKm5rvtTkZEJzyTb3v
ZlH3/g7ta1LWAs+1pMJBNIXygm4RbNExOIQpmyNNxbdxzpzUAt8iajqLeetRquhXNO5ajFfv8y5c
yu6h80ccwWi9/z04mzFtOZeyF4kiZ2m0BuAHR9uSCGjwy6G4TCHdgdJt1P+069A8/4FygH40qkWU
yiaNmB5u3+t1DkqzqtV5dQ59hZjbBWHVRcLrdgQQA+giAuxC9QPJ2xteaj3Fq7wyoSdKxum1szSf
n4awsZI+AvdwWT2vTwB9zfG57DZTmB11lTV9R428KBhxmbOPfOxLbDzh2zZWZckk/Fg/JzSOmhKo
BF9xzPNdDuyPb2tuAk1gepgpiEYmTsLeVheVqVB1KhIPJhCVRy7pZfEXh5JrWc9Zxo3RmiBhs+Sw
z8Y9BapTdHIFFiT78gb2uIdr27lt+nUKq3qZzsxKrILN7TdTjuhtbtt6aeo8H5oeq4/5/JoELx4t
WN8180mDdZBUz5S0nPwzi6upnhxwqhP6Uc7fVBOyP1r6Fe1Nyg7F/Jq/HtSmlfjvely4+NPiXEW2
+r4OJ/+vuC09e1qpfTJPe+95yaX36TcJ5eg+T4oXWak8Hh5ewYFucP825x/PHApp5hASiroRPb1y
T9HOqOKEg3eJREgPMydGrU2KopvmqlsXX3cm3jTKhvKY2OVQRD8vJIW1Xzw8l8eeZGKBIFDyHFZW
Mz74ILEVvOtNOjd9BVfGYFOwHTgl8vOmNqobbdlu9lDJF6ds8Lyc+CJtLbTP2VQhU2iPLKJiUUrR
M5QBvL/AAGHTCxlfsXfxPQQlUirzSdeS74jyQWpqnMvsRS6jrEoQ0nKxgod8cHeE+F0oNWc+DfVr
vpY9s8LbvRm56t0qeUC9NQ5oIQDKJjYS8n0A2EUvWqgINlN4nODtXWQgkqRKopNsh0bcbknpPkN9
zpBTSYADqXYa4PdLWEbD8jnprZmbnUy6M+GsBCL1WYMHZ3V73wClQuq3HxuruofwTbwlXu3UsuS7
y6z8GR5awNCP4kcv0KxVH5SHi34ICJJtwub9MQ+ZgDJ4Lu3HJ2HLVgBiWN5/2qsEMUx8eXVGpqFR
bfw7QUvPB4ze5rt5ScCVz7LYqt5Jy+0O/JLh1411BXggXuU/Im28Dvr+TWtEsUKCvWSIXOtJz888
gz19ZN38B37WEshZCrdRYUO7k3zsgEYd91szLGT1XORfKTGe34Gmcl0I26NHlm+xC3/wSDl4qpR4
GFU8O2VNrKXKyNmqsjHo/ffRwhDTZNOrYaBDKy1vlYxLmSJHL1ZAtOAX7cylG1QTrd9DF7S/7VUW
aSXrKZ5j1znTZcppUSk9L9ezB20Q1Z9mWx5w/WFR0gDXX7qWZtDujQB5j6GUB48UaGXPxdhx6Nug
/KfIS4ePlE7DilxgjUt5n8XEhETsw4ZizG+9cA58qUYHGMBc7XWdf/4EdvjqSejEEu+xOFA407b0
VkB5c3ugbzEExSq7uayHchF3VHav4ZTpIgpUxxCmViXiPAKxXT9PthlorDmNh10mHGAifl33tsRL
EaWA6+ahxrNjq/hceNXaWuTQ1VE12COhldz1fGuGfVqj4GTBAYPL2RM9dd+Zm43Z8JRB9Dg67e9x
dL+BMWZdtZwFHHaQ0/uhM1i/UYFXlV0OK8AgJyi1pC9Jypttbx62wcc+q/J5RTmF/gGvQGYG2dHg
pG/Zhx6yweOmgM/vw/1h6K3Rvqzv0I9OJHQ0ARC0ivVEc0S8WgJyFfO80SNhLDAzL5GlIngqeSFL
4La3fs7sQnssOkvTbI+UoPX4CODeZnFsilSgDUWiPJ5wmgypC+apXCGHxOFH2P9iapRhWlql0HKf
uL8XZ7TMBt0ankykqWUzzOZsEqyIt4GYzKEMgbw+1+DYVz+LbAZSn+xYj/irv0gSnrue5ftjQRiW
KisuMwo/QVMxpOf7Rm3V0d5P/RgXlZR0WwxUN/a1fEHLOHlPZUtUBfBNBEBMuK9tJtl43zK1+szc
AnnEkWMViZhF0JXr2xXRXhZ6icr7wmUCchGr/IiUm/TBQu7F0sRdSimTp5DDCEBeNDnoFoE2Bz7g
3e3MCPsEFGXxH0TFVdDPseCchgfT2VWtaRbzLzDi+ttQC153S+fQOWLaGaWqUAr8ABpQ4IsAY8HY
sc2qk/NJyOY2Eq+tY4rESWq8amn4sDoDX08WINS5HfXFVCqZCMJHTg1+EZlnLLUQgFtZAursMxTr
QHfFx/Bc8c4Wx71hxFZ1NJHd5xrxsrVcqim8iAQCoHEwR8wfcdGgksZgGYQJPSSuJ8cP81yhmuDC
VAk8Rr68xh2nfr+A8JF9Wop9WgvQ4oIT6mOEmQjL/f8Lk3gOsELQ7WH1AGnGCV7alyttfnASOhsC
XY7RrEF0kImCpgTGhD3JIVxPnKNMjbFKhE0suu6EVF41aymGz1dLB8M/AGGOJz7QolwHPIR4Zusf
2fRecnj+qzK4Cr++2yjBUpamLVsL/8G/b5GW0sdJBATHmUVz91dbXggCVwADCRMpsghsmhf8CTq2
F4n+OafO+Jd4mi/VM3zL4AyzyLB7VMyimGv0Oq0p18+19PManEbFZtFQWldDmljJoc79wkm7brHy
bYR5m75amiQneX4qJYkmyONsIE9I0PaljaQ06knhXtB8IOR0ipNrEjvArxr4Ab84ftUJC1lfuizA
JMYnLkFycFGSrxPLHzo055P4ztHGS8BJ2P+ySWZ/zrvi2gP88TTBVci4GPUzeyk3fdK+x69PuWH2
5pd1E9jHGvxwUFpwfO8fYrHH+Ich91hc/eWnxrEpGLT+yug7vhOoQohNT6wq5IgrKOCU0Vn0aBCv
xaXZvGumUyJylei4/0HST++hrz29BT/vcGTIVlO5772ecs1NxbFN1D+n3Dk1/FT0fnQF8bmVHa2l
7AFuppTshpj0vK3c0etfDQ9/ENZKXKDCDw5+pYtiuVZOxlYTWtEr6C8PqL1vaMDJswN0VhrIcfY6
pbOU9zeDVCA6nAx/e6fZgLVIqOmVVUVux8T4Xdo8ZN2zGwvNCBPoWYWLuzLPVHM5+bjSeSDczqit
CyeAVpEsj7VrY36/YFe6j7OlM3CvTkccKXrr7KTeCv78tYIGXKB4ByIrLtzPYMKfxMO2NHYmNzbD
YCuzWFbwy+PeKZWKmRiPTO4+bImxsqyKxgW0bl7vqXzJSG4it7dWSOjqLbYrKzX6ODjAN2Dmvaqf
+e9NVLNrSTfI6RUd3RXarc/F0S9KhzwfZEHyyth1C0/cGTpdnnhjst2zHGjakvUjMIgcfwOhbOur
vNxGTRacD1J4waSgRsqxXY54X7Aqv/wI4Y3G/K1gK4IrDkWUT0GNFr289o2W/pt0JxNvYI2lHaQ5
JNON/DNnMVyptJNuAmIyPtYfGtFihDY0OaMSLyKOj0ifznl2Y7rA//WiIdhRgPiwXmFPfAzHtk4o
StaOE/8JVsbe6rnNu10hOzD6AMaWd9TztiDtz5q1zMtKAFtK84h85mH0FXgFlmDeVYvsIq0NiOgK
xgLkkq0X2dQ7nWrkjQnU7fxT8cD6QpOhhFSIB8MJpwxA5jA5YQ4u/MtJChAOB0zTiW9D9KdcGW66
ifKc2PY1fyID3uoh03BIL9jcoBJzHQpT6HvKfmgNNK6Hq3dizn9A+PujwzM1hvHsZaorHZm6geD+
BRRgYH1CYJ+ZnBBumkat/HAnrQGzFt9b4MkUlY4M3Thfur3lxnQms+IWIOzS1W97rl2jWan9Q/vn
p3FHAC66S7J+3ELlqTCydJKjzmrU6YDzVw3uo0EBvGY0AFyERWzTOrBXRDzM0vPq7wDnoEyowqe1
j8NdRJ5Gh/e/RCPQzPFDmHkLcCYzf3w0bymg5WXmYzIxpJNr1JK7UA198uCrw89g6gLm3Fbu9Qxd
MhakCKPtdp/6hA4bRZyB/7yEHNT2SOsxpnH/0PTIaMC0omg7kSrW8vOva9AWpDFdbWocftGk/DIG
RP+bdR5ZM3yNAEGKXFz8+gvxooSD8x09yid2wczfFTTsMGRxZ2MUKrZqCrEVvAIgQP6sZbhK6+Sr
mb3lJaaODAUjE6UTAx9pg4AO5Zz41DxpmJthvlQSBpJqrG/hDP+tgmIqFa9Dzc1da6BA9M1XHbUM
yjJGVk8xY9SHHVmJRtojSx3PsejtuU4ivr0HogaGPwcmA4ulsrNySNcMqYJX+YpJ4Xj8Mmn3B4h7
dZhyrayd46edkfO1kVGoN0MYnfUIbsvhqIb235fBh83GaJoDmViOj7uPVFmpeDva6imgr29pcuxw
Ff/Xtie63ocbVDMgb0bTg0ubUXtcwVH9ZZhOvWT/9VVwtAld6n/njpXp5d4eX/kRz9DWyBpDA4dR
pszUZkSQ8nj7qM/zsWlquxrX2Pkb9uXgooy0e3oL1W6qwPb7z5+Zlx84PuhY72U28ypxOBxmTKrn
bWQl1+rNklfTOYvahtNX8x5jYhO6mivM2DDURmJSNaOiwUkR/ObkmyUFIUN73wzoorTBD3CH4tE3
EpB/k8LFkR4j5+xruLSXHFGMACyTPj+4DSmsn/SqsUWTunb6GUQ7X1rQhApb6zy25exxJ/B2jmdL
KnPwxMZwxRYStD8lRSiQf6L3e/4Hgn7O4c7vLJOLv8fRF8zqdu6KCR6ySsCQwz6DkgXVbAzdmSN8
aUnLCLSoOGX9uWpLgkrmbZN8Ouamj3EYE4nUMql74qFIhdvM+bMEydX0J75I/u1o6JWrTL9p38ZB
xGKqeZuCG/mJIG0UZXQPEy8a98O6QZmwEn0oMldM4VoOY5fAP2ye7Citi5qJGMUt0hItCE18hUKE
Y+lMSgpmnfGkdGcC7G8ZegPWmH3o9lUGugEwUC8JKMLNkCNMS31Q5p4QAhxGoEY9/7wv2g7U0pVe
lU7cytkkOa/2hBoI8V8Yjcuvu+jXw0XAFzrtCpFgaz4Kney2GLMO2lM++tB3pC0S+s+dAQLHiX6G
eY6nokaZgzpwVXbAfPgXmxRo88QCiTXF0cbfm8oql1H6P63LMN8pe2kIZDSuAM8CC83erMptRMaX
W9kpFi2NEaxZg5ccAEUxQNKET9E9BVTDJ5UZlmTUeAF8UnPwma36R2OxhuGP7mUNth+HRrdRXrxN
W/grafaF57B3SIzLTJSWj2H5QAdihawnE9NZw6K6LYw4SF34A0Ogw4XD87RCZIUigtBMEMgWPqiR
pJt2HGtiwJ0w9/ZrDnmLXIZtePCPbVteXC3ZdHrSlWGHLHTEod5PGjVRcTwaGjOsertVlZ2Nlle/
gQTAPMMRqBIJjblMBrwZ//euHnkLSIui9TsAo3Gv/Z+Fwk5EmQE1ndfphwFiO4L0m+yqUQfoHXZF
J2jrQ1iNiksEu78ikpfuYke2yKsepp8vRipdpN8fD6FyQG13SbwezMzrEtjk6RJEWCf+tykcvgtP
HPhLymEGQJoDdm3HabGOhZXJdyYwOC40S0gWfVpK8k+Y/ZItEIsiAS18TerBF8GDP9htRIVnxnXf
ViSi/25n62GF679vGhrL0uTO0DFqbpT8+CGhMgE9JZUKDfz34nrha6VGUREmDCe2zyipkOM+YCcN
szQv6vx4duatvGhyEIIDhIyOZoo4PySVp/fKe9vN7w99QyPo90DKgIk+qXsoIKn1wnxDSpMxxOLF
/Gi7Yv4BM/Xaz50pX2EiEENMIrSKcKRpdxKTlmhn5KdrloQPlwrgVCaqXgkABDVvYuTOfLtK/xT3
JTHS8aPMIOSpC/8CSY/06D7yeQ7Pd6kaDGu8XVbyqWX5D08f+QY4hjftMP3+w7fDgD7Jl7zPw3ER
a4ZG0a80RycFvOdAjPda04GwhLagwZAGytiou7lglnNruUkDpG8hnAa0pAorRmkBW7PR6/3yFDmc
auiOTebQWoOyVorHCxX1OCORaygbOSKQQhIq1k8ks95S0ObF8QSAfnAHmWCYC9KxXrhrYIFL6XRS
hMv6WaSJLVy83b+tZ3XFZ246euS5DUE/iPIEX7d1AvdkNtYYlQpXSjSWhKMEt1vqgqO4rvpAJNXB
mbLxBrkl/ZFmDvCw0AlrghGVU0scKkFM+047bN8/TV3fF4u0KUujhwJHZlF1Ir6DW0vIqlKGM2Fh
yX30O9HwWypfbmpT7nF7alWVz/OxkmkW67m1a0TW2q2HtHgufltqHOPcGcH496r+0+zunYwj0vmI
XnyyabQkqSyYHtvhjougsypPzPzQiLdVwYa50NYalBmYWBrUtPtqWXUa+SrN8ZK+4vqiNItJMzOX
vCiHZ7z7snC/xBGhKQvZwuECQ2AwEGQJgC786a5BUKxl9PP9UWJkFILOEXjdLz3unRfzA7i2fz0w
mKckRkDV2YYz/cUZ8QsISuDD+3hsxUqFoHj+oke5qGbfGtzlknhYdn0jwFeLIyiUxdopEUiSHuQi
mOMi3Mhqk/c6IkY0bDHOrXJq4vt4i+6Qff62VuYK4sZVo9M4t/kojpc2mbSe3kReWqU6FVDA70KJ
sdOR1eDeM73/hZs9l0doEwDcFIDZnh+bq1/iKRm8FEBWuHTvCgdw4EmHgGLMr7mgNyRI1YkRoCV9
M22LeFq7e2q0YtYLAT4LRd/dVOogUnrCvXxNoU4/6po8gPbCDUAHjJHyuK0LCwXMt+vtkE96Aw3W
uu/hwj6Hp0sAFi7U8E4p+u4FSwfhrMgml+Kz6esE42mqfkF30SgtgeHaJB3v13nrFF/DMgf10WoW
UBwJdzQF3NEUusJGRVx8S72lWZpv0h0trg+GwxsKsW1uw/JpKYWjOoNS3iFv5uwvYEyrAi1f3xHa
CTMupk53zTa3Npcjw6oMAhNID/P+HSqnpM4ZAvohgnt5awi6iuwdSK8b6A8Z0FhSF2SzSiKM4stM
HDc2of0KxxvAzqcqa+EKgN9gllQAiUsYM10UqetSTN1I080c9facJkjXJ91yXwtKfonTq4UjWfZ0
GwbdG0gj93d+wihFS0IyWAyDquflGvrELZbSuWjHtVvaQpdIUP8CCqD7jNZNr/VkmTEZXH1KEtPW
kUPacVmGe0rZKQbW+glMQL+v1QVJuZRQUexPoITUM8RlV6QiyRevLY+6ET6boyuoJH0IaS6rhAK3
7zC2HyOZccuMy53YgIi5VCjWVUdHN40W1Ylkn6vP00eli1Md1V5Epcpzyat7dNeAwz2w87vi/mUS
0WL0ga/T6++ov1/tCHNzEw9nw54a3aCYFAHrje3+seeb/lHQ0NUaDmaMvOfBuNbccESlxiL8T9ob
D9SFNjkD3wPB/MmUzPH8P4NyQfYTfrrplbL7LL9325+kB0bjtRUZIKH8AEtgBbbT+6VGQKq5UUR1
nVpPxI5U6/WH5kR3RbtXMaYBNpkx9L5ReH0MNqeFvJeXAmu4ccFoygUgo97rH37brftPCeuGdVos
Q3xLAgA1fi/MKpySXU58rd1+uWv/WeRUB90bP6yhrms6j8+pGwZ/wKjRr0UYOpTpEfESKhYML8QA
pwHsj4qub/uBzJ7PpRHPLH/k5R7VNxa+qjjYaNY2MKGf903hoOrvtf0b/sb2GQkDTpeRj93VGmBR
mXsc/FDR2pFrwxOpu20tJeCXupMIu/IWtjx25Tu/uGjCY761yN399rHGdFzooycrpdGTvKJFJ5Aa
8C2uOktLB7pE+JmczMhzzJWTDIEc+Ewmuofqsf+DiQOJo7OOkpOV3yvMO5IMjmeCmayShpN1ajxk
gHik5DJvuu0RLCfgHm+j/YsMXM7majthN6MeC6qhjbpL6kfo2nKFbRJZ2vNr6Z2JkMzxBIaoUZ0h
6hd9AAB60dIrox3ehZShoH0zVkL8i59BS4s3IccfWWA/2t6WDJaltDZ6ytBjxu30YN5C5f9cbV/6
Ws6fznCnB2eqAOfYi+5jD4sJK9AIAMzJaKBqg20KjFkL33OS+spmGza2NluJwptnA7YOqAigiPZd
/EuI8H6f7i829CvBAhOCvmI/FoaclyfyDM/KwDFblWR8onCJrJ32hVG1GOC4wmkHpx/Yuzb78iU3
g5rbDsm69OEApUvzmSIjOh67p9REjyuTwb1e9IlpebT0E0VkhPQSHRiqk/LUV0PRuzEtVlBRE8BU
esBs0TQ4yRolo3sHtRhCW4Z0XEn+hAyHF4Xkcdc8hSgoz9CxKmOA/bzLLNOAhyEc6JdSTjgBqp0M
hbWTdlhNgmNMGkLoJYe3B4QLTW57iTQv4svDTNQ/GwCzaadb5LFQhIxzQ7zMt4kRu6vIruRyB0Ho
o/FaJFPaJdfbJ+hn/ohymBSWlO/CthAsl42PtFskMpO8E58NHZdLvzNl7+SKv+zVUwKyztmzmstZ
n/LA4Jz7x8n3hKcrHSHxgPeA3Vo3eVnCEVHrjZzom2xLU5Oj/HfjB3oKcoEFlgw6LyDQI2W69Vqe
xx0VKR+ZSARK4wAx/BMUYtgGStGr8bFUQmzVHhhoWOjjLDMkrPB+eeb+nmTgKHTWWakRZRo9fs9V
9qkJRmPmO2gj9UOV3MxNyaR6lDfWi1bUToq4l91E6Bl0x665/wtIhaMR7NJ0LoOPMEnJs4REE6vx
lC4TRdtD0Vf9aN/0EYmWEXauhlVu2v0R8xFNquxk7jWPB+YeRaH/ZYGKWwYafeQrzbAmJq8DwR4O
sorLqzezvlznLa1j8ASvCAMjGZ9EYA/Cp+uXRqxdSWdONuQVg//fAQyy2f47FlOIlE+5iHoV8frC
ZA4g+f94xL6rg0fD9Ya3eMKqFhW1r4Y6VImXrIB9QVc1TjGhjQ1+v56x6TseNSd5KHOYl1LGDRGo
QAcYJrCYp3gJ1EwqdhOglFKdJ+OLwK9wh0hrsq8ckWo0LHwOoni/PurS+0RIltrKKrsxlgvnJVkn
0xWQWdlnQ1GhNpPw3Ns42JQd//U+iGwQFjwArOT8ZEscR3ACIsqtAtF4RGl3hZVIo3Ya3TzAhWqZ
Z38b+FlAkQY6cDKGX1HsNaz/9TN+/L2kmrqNkX7EqxQN1YBT34PBny4MqAND55Px64tliL6SwvOr
WnnhnaVMRgSDXkLzNPkxRFfz+QneoCxtEL3Q+kTRyk1ZmXEDctmh5d6mFnuebFk5Ahw1gu9hlcxa
nKoM6FcWg+bsH/vah3FP3lbn4d40OoyUWg+ha43fYLH+9S12aRl9zn3+b0/iE6+MfABrtXGdUMG3
wfVy48R9aaRL2nQBHzFMv4lymhLL1N1PYbwzrU/wROyWq4tvJbQZ8Vo/etS9Zs1hJb3BDBc24GT3
gzrL+zn85WZAW/XJL3WiZE6YXqEBeqmuFbCOxwfTNXu4u8C05O1kCZCZ1AepoezOyiObECXpl2+9
DueaRBuo7fJJJ0ZMv7G7anH68GvAzvdN0z7LrUO9mR8mhP6hc+wCLzyERLButTPuFKxVAzeRaYFX
fwUKn4fcvp8F6hbQwKyE1st+HNOu2ygYuHp90WqGHzaejmhpR+YA4RUADN73Gj531yFHw1z+bv/G
Rq8Qhcbtxr/zriFOxXAN1hnrx/t49k91FRsDXfMnGthFXFxnlaoUSwTD6CNk5Rfy66kxi02x8ldi
XTgyzkPoAZ1FR3IGXcSBIRF2mliMH2CmovYftfI5LSh4mzjQX4Y1l56/1fn1ZUScgyCUUpqMmnK5
mriAzYTCCyUYwQL28BvUmFcnwYM7MXmAf2mw9uWMGrOLx2DrPX/Vq5BzFIi3uCyalZ6ucQtvtWHr
viDOW77PvuGwAEOXDx3SRu8/uuKNgrd+6v99M17ewsbPYQEZiXMdVjXSYVjrdlSnWoSwka0bc2CA
M2yqK4QmwG8wYD/ozTSWxkq5hOTjyyGC3Li2zTfZCcehWC7aL+YEceV+xst7QNqzMhGUZV8DkQ4e
R/TVfh5eMMRwxvS+iBMCNE5o1yLwzBqBMvlb5qv/utDHpY6KxYLHfMQ9I9+kUd4ZQyEyO5hQ+G7s
bTCZ+ACJcFW7M8o0kSfIRZPEEb5C5kdDHNsnWmFE3W6+eno7C4JRvXgBQXz0jCV1i+6TzmoqPlnG
ouDqF5IXV5I7MB5sAlK/XvUosUYgqI8a6eyubYWvDTKfQNoI6kwXc1/NJXjNeEYPFreIiiOwf1RA
pt+gFZWHzi3MJu8XVPxwDjTHjSst+6xChaBc/zBcwCIVsc7aEMPiqjzMYDZseNODkUA1j4MoWKSk
Qg/v4X6JFjTd/80pGCi6FpZKo/5+kzoOadprxUBsZrF0JxoDA7zhJPcOe522Wr+wOJN15dMx7x6D
wBe969tfrmhkTy9dBKl3Gq/CnjOCJKda1Y71xmEZml+nJGMi9xVRP8pV8XkKR8KnRx1s9s5WO4wz
fyg5iHLSiYd065qjuNIe0A6qy6Mf2v1uhsbkwKheD5KAz+HOsdofyB8Qp7OL9qsVhDuEJ5DTqh98
DkoBSR4RegM9yfbM/8kf/LnelYWMF6ka1crgkJ75d5+8288JVtxmDWuF7ZVOWXfjgkfUjznGY+VU
dMgToFNoXVhtfWQTTiqKawbIOSh3zA81MfbNNQjx88sxfRVXLJ14ea1cAONnu8wNGZmgKRIYJbDt
6Oz/5FqRgjaZAmp8Y7hj43AifUmb1I7pn7ApYIqnn/RZ/zL6SPCQTp4m1DvVf9vhFpCvu4GkyYHf
ytYSH1ni17pYly6WfXb71KgWX2ylCMT2ShzCZceD6ivFqVRfUUQxtAqDFBtqZZVh542t6Cefw/dr
AkX72HFP9xVKkVbB2/ZSf2LThtYRssPX9qStb95jiWoSN4hg5QOXVnp43DzxOF7hbuhGWJQdGLRq
a/S/rptAc63X7TU6HKD2Txj4Jkg7Uv/M+1UYC6ErPfTZQcupYxGU7Hb15jJk7gpFJUbB+OmIWQFb
O1byrhQnOcdqpYM4bs0t1dPEo+1yFUQSdrwL7U/xGVR1B2QanHqivGXRGbR8vSNDTAimOzhDMaEi
jFMxziQ+c1f84MH60AhOGxgbT/+cMRfKuQybn580sGi1tOnPgYRN+WHzcv8xMetywB0UXqEF2heW
gqS5d55XEE/E6X+w2z7ykCzLU9pLCs6QiumZywMJesoY9NckzQobzm+NzgGaw9PYoVk61Q1EMcLz
QUgVE26f3Yd0lNBn9aroRRhNPn6UeYCQETFDWCpWs3LY/+OTCiVvkqxsJO7E7/U4VMem5+Wy7YVc
nEnyO7+9AyJG6gFQoQq9UZG2rkVDot22aA/H1szPfpkRapZ3BQ7iQUifbM31gRCO2Nb8P5JntOb1
qsV+3eHKnbc0ueGXolRRFS9qccpTX0q5JQMPfKtnDtpvwUouaw8U0UZcS0+eYfGHmKJsrIQcAsCx
UJpz4/Gcv9h7GEuaU75kEO4mx2c8oCaXiTAqrIR4IOsh0Exe0GgUgByiF9YgR/1F8xdy1QQO4iyb
yKWSZ0dQjj6vN6imMpR6OczQxWH78Fz0ke9rRMXXiL64Kf/I1NAjVQLtfe91ma4N8uvrWpHzi7n5
HCrc9aPKhsA2F0Vh54tKiU3A4/GLXHq7olcF5c1lt6aCrpCp9vbVcwwgMMQLSjrJ1m7UgczeGI8o
aOG47KPL/Ch8wpEVUsaF6tojo1ZCo6smzW8QNsfMTn5YDodlz2IEiLo9k6AMEE4OW4m4Yuqv5lKH
Egp69ElvRnP/GWxCZDtdTceqXiw4oRt9ZkUMucK70SAH7o10t2W2GR8ztzPDEPkd8rNUHG7DuAcl
odP2IJDdvJ54g5dWKGbmarP/nEOOtBzqS4iLwwtc4V27UjIrzg1e0es6PYJNUuMMBNPzWhr2652Z
ymVPgBlxAvehRpi/g/fuhOWAl9RxQO3F/qwlBvavUg7wOzJKNaceKfX/DxBYGzqSiiFW1ZmSFljA
mlj+1APTyZnw/HuUqhmEDFcw47vSwtaXiEe89OlOjC/ifR4/IpDXo9ZcQ0cZ152HlXXnZUuLP7Zy
kse+X403knvRYpllWUv1OBPkTJAKNTO+qDLLAP6gx951CR+PTT3M+0xQKZzdt5/OZZ6e1n6INgJt
TUGKMWN+SY5H4L10B+OkGd0f0UKOTgCqKyuS/BYtQNuoDtqgT7QClGoGkvb/x1pSH0RQubuqRaB2
B0gJXlErFgVYxGGvbDKp9U7x+MyK2gQ/eWu9EmjvtmUn3dQkHfN+ZykhUX0CqqUDhoWFVQ4v6S/o
RYHDWc8XZV2df7JhUm6EEZs6TRts0riknjzPJeZgDcBON7OLJtfogDvxjDw3a5I6VM17BERmX3cJ
DaFqAb4AFbfP80T1TE2N3K9X0ALyMKTsEx5noEtY5tSAXloAAKU6y6QNBzbls1ITjyn4xeyx2shK
r+gotMX2xxr6JM1gK0rQNK7b4lLFwWb9So6RYUURNHXO/Aqn7I3NiAk0HgSrx046+CKOgbN5sO+f
0HqvbTuWdDMPNTLY9UNpQXaWasQnTwwvsKUkgE/2tOizWMSNuGDTlFfPgmKdIxK6WX8IuuDkAHYi
4y3NF2lFlCQ0cJXM/fJxY3sYDkzhYgu0s629wto5Pn4UCe5Bg9tyEr8KPBIl1Md6LZ1GEoLuUwih
kw/jXpxgbnij4OlAvJWeizDqa9FMcbseYWAjlB8L4WNDqbbi9rFSV2KlaigAJ3A7CTGA33Ib5ASz
HhAt4Fh3kk0IAzl/sAJph8C0IQWxM2gtjdTy7+SvJojtI/Gkm1CO+tMc7inQjCa3lnEVhoDQFIX/
ycEsclkaS2sW0rnPtKWiFNFX94xu2ZHPXmx50Mb2Wi1d6R30h9X3bibwJwKXmxKiwZnwfaqqlbZh
fa5mLwQl/8Wt/AB9mj+5U6CU49xdlTLmomXK/8loDxIg8gVId6R+2moigU3BzFqWj+4MU6TAmria
c9fmqhcE/0medzlkFhBKXEg4KkBCnuD6BdFyBgVUoiZpasfZGW9ji40ICHtmVduT+lxYz+V3WwEr
+f0XiRblhnUtq8JlihE8VHZng549Bn/e2NIjuFfm5hu4az/MQtJKqeM78UdJchSw40+XDARS2zbh
yZ9HKWiLbLU2tD8gp7F3Uton56BtaNeXdT7xMlJOhgve9zr5W/Pg1W/7gzq4d6okWozkg6241Gb5
cMxFr2PUWgTdRhTWdnDjJeOoMk6+/IMpPS2Gczq4xDcO7mCk3dgR6bHFKpe80Vo1zWy2K8SlXDFH
p6zI5S4mFYugnwrScqQkIEJD156sDboetZaj77J6TZxr6sqmG4GiACgJUxeJLxqUd38qt3dukKt7
73phfSnigqYtgVX1l1ulQtRUKy/7DJPiJqvBZzJl70C2Qja8DTXXNceBSpJSCb1ivP0uY4dN+ufu
7Aqd39ZQnLT6ifsbGpt7MXRB2EbUrUY+auBbZiWDBwosyZNqpvcKpTQTnltq8biG2NenkGD89stP
GKMieptF8YdIVhyV0bRntZ+X96ciHVMaQ/NLyx69p7UNVKvmg7mje2bZB6tXiTEk7CvyJm+Wkpmi
O0HZevV3jMmJIBnzeWzzlbR7UncHmMF0rzP7cb6bhJFKOX0nOTFdIHg5L3DG9ZirvhpsYOiW2Sbh
L9I5zkz1AkOwwZusNADnv+C+VA8P46oyMBuvBvJLVZL8bcy5SkPPLhFeCBYTFagqjGLiYF7U1kT2
xKK5N3zg1tMjeZsC50Lkluu4gzP7JD/BE3BLVot3CH4btD36TaoFvqNu3mqhYg8Vc7WJmBMoxkDz
+JVUaORNDRQqLUuQr8a/UzB50B4iPdlWzYLg4+kklG6M6TbykKCmpYevuqrNWJlVnpdU/mtNPH+i
sEC1OmqetaHgSClYtfd7/hm42Ev5N4wkYIPiLXvHRZefgVIrYPr2yrkm8YonjfapiGl0PHatwFWb
i39+5ksUgR5UfcIy6DPYqRwKyCeGH6YYMNV7JsKxWs/oj07cSVCbpLHZ1kTdfswucKDipFSFEEL/
rufx/M4Wr5724x00MZ4podcKt06TvzFcHJPfdJNmADFHDgk3Sq1EYugQQOC6QX9gkqLDoEV1CfTs
gKycuYORAplMQRUUSoBL77zwRa9bX0IK56sWD7ZdnXsVLSZKHR8DEI98Ex63l9lbOp+kKfiFRrSF
ZVbS+pPw8NwyzgF7eiBLWc/LREi7+AGKKFIAKyLhg7nwXS31dXaNIJ//tIO0nVFXQisuklRUhMbP
DVbFNObe2qrtZ/1NRexS/ml7K+M6uH2rh/uTNdFgiZFCcjQhtwEeFan1zFKaSHqjdrT0XOp76XQD
rdg5/ivEsZ6stL+DqZbG0uV0myRR8g9WI1nmTv2Y4hoeBwJIETmVO5eZhXWbl8s34Lg3RErqGgcX
diA/NclkOdweMpBThIQCv4eeNSNiLVy/guPPXMC2pV8HQzjC3mMz6ZKMsEA/jCeuTI+U2x1r4u8t
EVfkahPTDpuCfmWy47iyXFxw30i3JBhmtbPEA/54ty/RllJcymlQpRoyR90q7EN89mP+DZm82z5f
iQOIHWdvvcb/Fjea9P7UQxMEcnx/8nZDt//Wc2nAcUjFFfR/3L7KKJI5Sy1Imkupb2V3Pm8vM2SU
osZyijarRnVbOac/psW/k9VOvPh1WLMJQq1DQUAJUFHyJQttnlK3Tllk52fnupnBulA/ZoiZQr1c
0u8bgeDnrnLar+Vz2P9y5KjcD8NM9iVoLVVircCh24T4+VDlBfet6bK++j+XbjJSzf2sY3Cz2hFY
cyxNmEsfUiKvI4V4XMKViUk1YenR827T/pNRqI5CCiMpc09KaywWArHpU8i318sszyLMzLpJj6Lm
dm2dIpbemGpKstjSKKfILu1IvljdMM1n6Gj2N0pCR0+xOaD982UfstsaKlVZIcojmWkWkywWYOb0
iZxQKJV/lHwl0MSIaHKFE+YnL5bZf1bh2NxSvnPn2cKbvGqrQWnEDeOcp3NgT8rQ/MT3oqqpTRZJ
/drpYF5gsvfN1I+EEhE4L/MpvKsN/uQNCa0VrMn/nd41koSdMl05zXEovlfJ2HeJSpQ/vsNoJzbW
kC+1RLBYLODGLGjkqt5B2ZCIDcf1AmNvuj0jHQSzArnSrelzCsoAwmIQpE+BG6pr98Kd6+XbukVA
BvkHjyVDV579xFd2KfwEWwtEf4ImjSnOcAt+FgNoOL7UBdFD5m+alhjCV9xkdIMiH1LZBhIMcDIO
zAjSbZ8CcHrHROz8V/RR/oVijtxc9IgBPMcv1TzmREAh1spC+SicqoolzvFrA43Go26862sDke3B
+uqBL3U6Nxv26ZwKfJpAEzIFz22d0I9EHm2Xz42023ZjbKp6UUSQMCwVSqSFbIutahe+8lS2GEOO
3ZRui/8VhYaeQkNOjOpAZcD8dwVMz9HWrxjbauYxbWBWm6LDpADn2L9C0gMajqlmphlif+ULdWV3
9dyR63/lvwBxbI0tDHjfSuBTiXJU8k5MYnEkhcq/E1BdJjCdAXsidwWvyM/46YaXz9TYg/d0uiRb
VzUvVV9J9Jkw4xiUXjt5rLhGhG2A3RENePZksgHvuHgPmCILswUhPmVGdOcd5LZcVTL7Ss0mQZ7+
NAWYkjb+yd3e/QiDRgU8Gnr8dO8exspt7fnCupbuQgT7AIZTW+OimA4T4A+QU9WPMS9VRrNI8j4+
dZFlUYwqHxJG3+xZ9+Iq5Exdg9rwFH6lD1EPME44ETuDEI2N4lDFOUe0Nm3tEQKg+mMKhjrdY/M8
1HzN4bYIsggIkeRNg7299DBTN42DXV3ZR+z5BSodNWQ9w+KNZ95YiMxXvzZfmQyKHqPinLPPcQ+W
hcsJy4NTky2WldP95w48LtjHGTzdskMI6alAVRkIVMpPZl9uBrwxUZPG3Hcew9nmX+Ca1vqMHXwe
xr+ZptRIrnZ9ERA4vrcofNY8hvyAaOCwl8XJAAOgENqh6nCMAYLDoE+JyeW0HrdcYpjkCdOUX8Ef
rCKaNfAxOtPFcE5CH0LYtIt/oIwIp6c6tjhGUdkfkoO9y2no1aowVXbIjQVUPIOqas0+fnnC2r9H
DFHq2BmfuecBgXFz8b/0Jsp7ZEibySWf3u/QC9x3czbPruPvVFuM6vFwM8OFfZtpRloSD3/K4WcY
pILrxe2ylEu3Z/L47/Nlz0cjoFmpmjTuFmY1PZx+I4olhJIXfhYJb9Wg5A61naF2r00V3fQEM2fY
qETwb4w3CdV1QATKM/cTrxxmPT3pjrEHmVlJMvL4/Wh1E6uLoDUOgAYUbv4w86JCAlUsnoteqD3i
n/W11izqTheLHHYJhuKq/OKhcko1MlVQ2wtS2x9QZsOij8wCfYH2HNTqWFmWSROzjZ5QvIQ7vdsb
UuYLhHEbsbi4okcNZ54MTlxpRGDWLo9eA32tajJt2OxM6468Tqz/WXQOjCdK82MaCcxWgx+vbWAK
irqDtBSIw6dPbKfFuVi6BN9AVMGX+4tqnIfnUS9mLfIBQFfL7jxxBqPW2d2kcaX1PG97j2ZDNcWr
/5IQVK4ybFtYcNZnZ0e0Tlm3g0ll24ZoQ8sVgEb5aYkHWkqrsCPdx1yCQSrVwy/wQwp7/P/2Ebek
4OknpomgWarW5BjOB39v5xe4Mb5fRl7UY2x8Hu9Nn+YP/pCj4Z7JzBKrNMi4zNPl+vI6z3nru+1E
DUCc3hrUanCXekFa6VAcD6GCo8mOTt/4Me2jxqRxBPrGzc9vl4C8LBW9RSY+Z2mNhq1Mu0DL2vxx
1z/n9vqyGVeF4NenJ4bGyUydLFJyi4GWcxM8lQIXNugHDjEmwY3pVElXKqprp5kIktXQSplxnm1M
90KL2XLxCkZDX4XOen69CIF/q5Z/eVNFP2+ojg+8xnPe/BI5iaqN8VE8Lyz/bBfvjGctG1Aj1VIq
57AoXMnzVNSr1ZZRVOMLzWEStYdRzF3v5wb6VNftIRIhwWUomuf2uz6RSjbJYfAuigEJ/1ngbcmJ
iqUk6+XBBa0SBYSXp2z/yezRdXFldhnwGpyuDSNzlhF8f3Ovutniezkv+8gs0uRf+7Ei9EgimL3z
dvh6nedogF7Od1OZOgrc7M3PGE6Pbd4XjAxNacOVUw5ejCIoZs519SCPkaHPSdlRk3r+hwamvArf
HhjuNU/AEDPRQybzXctOuL4GawWPX7gXLc6UsiVGx5iT0dfSmm+UZtIWbydvnrnwQCacwDia+d4O
JaBZ15yRmdHDh35wTKNAPJnYWSASgC6kerepIRlxX4MWhoUD94Y8zgovVWcqSxot1OZ4ZspIK4Im
r8p3Suvmsi+CnUlFQFs39YLooEmWrvOOeZpuExbyRI/qCTcLAKWf7LJ92J/k/CIdLH4QLLUppTJo
I9FeTxrY9RE573jXRbQBF09yW+qwRRP1YEAKXQzmOeSjMwti+hWWLENmdK2hxp+BldQ2FqG7fvVD
ZP9ZitFkIfudQnzuxYZ39mV5ba//+sktuACuNJAg7vStofYj5oHMwBpQLTyEmVtFHKyzk5nHzuQN
e8L9F75SXZxVgtPlJJQ+eIOAjkzkH5XlBBn7DA8fEnNAYQl+cY+XXtTWVP6gVlEL0spuR2MQbKUf
NmE7N29MM7FDDOsM3BLuulFsrl9zPjkaHcHboKBFvDEj4u6seeAmhmvne1H6xCebD45/HOXVIrEp
lFrP1JXRHTIpDAbQozU2BnQv5hSVteO0XOF/msqhK/UvDXwbc+obMNgRUToSzP9OqwUMTOrMNemD
57pV6G/1EDpeZ0nIt+wb4SFHjqDMqVY/2X45sIfR9ihPvH9nSeDY9z2Kuw5GRTRPqtr0Tf3BMwDO
F+8eEf4XFPz19gK1mnGgaiEFnkxgaqZjHVE8CjuQHse0u5LPTPyKhnuIgIFPFlEdHCzXnDKeLPn4
9met4Z3nbSlnpTwalxIbX/5VahKgDMH8mHsJ67HE19x6Jg/FcSt8NgWgucxeGJ+W7xrbIsv/gA1p
jT02b7qkvBC85FhLSyFh6liHN7e+odiM6ULFSjuRr7rIjVOmxOagwAahgZMBNXJut4EBNJ1Gy9gM
XhyXEHWDErqKjIqQvlH8EEs8oKVABDPUOqVbx3kXD5VPoGcKJj1QOrlgh1GyV4YNxeGYjdOG4N5u
bR2f7PM/+wWZvpsAycheLSHUe7iUHlk01yr63VUmdH9g87V/VaJHRKKkniJY2i8fu4zV+s820KNZ
NjifApu8426jNS4L746FmaSuyTP2It7AK317rK1aXzHI2B7SyDmuxdxyF61lEMvx9rw1knYjfWYL
z81hV9XoMtE7VaaW58d7z+uBLMrN2aw5X/W8VM6ezN3UORZlAmtJkfLL9kCktOGyzCjMBdFFYHQR
YB0fEHjpqqisfHtLi+55PRo4jh1psd2OZoAqQ+qq14ekAWreXucuN8z+IX6His7MqBQACF7k0BK2
KcN9LduJeFf2pI6tdFI2jCOK+EokwVw29eygMh1l/5uVAZQykEwiprwpG7VVNZycQipgDz2yi1Nm
GiGGsdtegnbzoAw4PlTXVcV9gmpDCBogKoJGf0EIjyyHM9n+bdzV5tdBJF1i3Aue5bnwM30fFs47
gudHkY7AD9eQut8I6jYmoCjShaVWW03DtcOtSGnhViAvSv31alh+heiNtCsQt3csCIYa3dWNZlfh
zhs8+g8N+3LdatuUqzZueg1aeqN74hKsYW4fZQZF4qz21fCAFWWtFTnEqFk2jJ88TMUPw4v9k54P
/SfvYBE7LMAr8nxqmYdcwiu4Q3KgpMiTZeEY65Ne01nfxHnN44/rpuW4aSXfMzrgkTi7zpBqiCIc
AJXSUMoVf/huenvDSysX0qqfY3ZfXrq7g9gY89hfWPC6Jv+haZiHfLk70b3sO2NxOhqIusSWDbCM
6Ctlp0VgY8e2I/aq+gFo0hlLqP+yaI7dFJWlxKiN7LgdkBwMFkjB4UzX1LQJ8e07p7nsTv+BcLOw
Ljf5gG62wfTocfF/jNs61ggeOuv9XwesrRfVsgDB5RE8kdgdGX1DrCEq6dAQ3omSqooieVIwknzV
cveYFoJgMSHaNn0/pnyyMCqxUkHFvht8gc5QjQHm1L8FeJe+vn//bKswvdYbmnuoKaeGYMiwN4RG
dmKSp49IKwvo7EMbOuGxQE1pCkpLF9AfwOA2mzjXGyzj5InogG8MjtbFeS8PyQvUH1B9iXbQfFBi
KuAgjL8aASb54923AmpBKJAHKALtJuFN8s02V9k2uVrTKmX+USVvnm6lOXsNLe0gdyRoOJRyUDn/
xa+UEhdRPV55WXuD8jI4VVDGfTx7uUGTyF94c+YKyc8TJvuO30RPOE6gVW0q1TiYZYTO9z739/mu
L7EvAuzd0VNouzR7MeVrCdcdp/YA0QEYBy5vcmBbp3w0RIKKpXTf1+WrS9ju+od0Y/VsP35OTGNw
pDqTgxww4TF7lM7C2SiMvNZOFThcnyiVtR3m8rqW388AJXys7322QOJxACWJ/mfaau9JeCwX0t2z
B1duDtNXykqeZhbyeocgfhu7yXuIcrHHgiPltCIUmLy2lgxw0TtgSuVF2tQnifUjH5z8EGxm04rz
0fUAv2xISQvmNLpQ1cOLiIuzPWQ4xb2osf4Av5XfWDA1qKqw/thXYgWiQ5xy4lBJe1zJrzDOFiQt
WTBcq8f3TUIkrlH1V83o57P3O/3UT7tn+pEerJP3B4f+6fxJwVBhu83Eu6RZZSkZajhXDvCw3IH4
TlbzP1XZTD5cB2T+do+vmPtRMIBTqHhelvq9PveS+tEE4xivP3iRNcnRKEKfFBZnv3qsJYAHZeHZ
Chq6iBjCWLj/EipwOwroKj61D9ps8u0nAQI2FVSYaceO/jgTBLJp8Mto6KVS1dWMLGWY88dk4uO8
XGRBwK3umuXT5MZt8HHnFY7c9Prd/K/9WY5mM4ZBi0iDapL/DuCiFj9RasAND2cDgLfw5Hq74BkR
AYEUlwulAxa5FypE5ndFYnCDfgUUDYrMbcqGW7KlkckA76mSVxxZRlzkQgvRw99PTCy4fHWOzMSg
0hIiv9D3X6hUorT4U2ZNn/hciQOVtTkuv3LZEnWXxceKwb84uzsac8PR2E/71wlglTRsalFT+AGf
/RsalCx4G/PUJK68BSZZr6RklPobw7mEXWBRV9cSw6ZwWIs0OaAwP9CorKTweGdUDh7QYx1Je0zy
onUumA9DTuAe49nUZRyudzoErFj+RwKj2HMbZmx7880SaaHenKkR1G1IMobHfHTL2HAP+U9oHhN2
MiGqyWige5UIFbQoxS9vL8d+8Lzo4XBFoWgiVHbAH/Ie05WSPDRe/sdHLU26mo9X6KzSSLGUMW19
0QenVB6TPhyus8lwbzxfBatxNrdeq6/nx2NxaEFVXgzTSG1X7/zE5p4RPglHrmXQY79Yvl9qnWNY
jDbV+WIeXwnv1qMWWcWO7Gp0H7wRISnGbO/YTBrQ7lHPrjo5HzAAztF1BCQDYVVPbesuYIxK/GVk
Rkt4zZ+fxexMH9IQx2wmMQ/Lu7qUeP+QB3AvHX8ZisU2plJBXNg49SObZHK2htLFqvh6TdOk3tve
2Vro0XBnNECG/9inaYYA8PHUcojBehHlVFM5GvAxT0ZNkBzq0SdinjT/dQNTfjO3Z/0J/3O7T6/A
uSl/ovJDp0NMoQ4s0N8WBFo4uL/gdJhiBZcr/3ZuDEAkbjEjS7TGC6izCtmT9SDEsVGunrIpmCRP
LqWum9Ly24k3T0bGEWPUjyxBNCSOcZNvggNKrhr9AaBD6/rhBNikqz+nEEQmgUyw+cPNEKaKvXpf
YagqwwnYheBfzJ9pCvXtdZhRNS0m0xj0I8hpTo0la81WcaucLNP6caH8PT3B3GYHJJ3FcGiwtzyE
YPtmfuzj8R7GluZNhFhfp1iM/Hv29YksUybwsMhycl7wQX2l3hnY/MccUuWr1jPe8fWoS9FS+Pfz
ll2f56dj31u4EOlubONg0xBmQ2WgyHa/pLEOIQ3hCkUhesKV0IAafJKPL5T/cZlKsdyqj0JVjzPF
ysEu1iiMBgHUSpR100mHCsZuV2p9K076LZzTLGyas6Gmk5c6nJgbmUZE3cNfCHyTwmfG6JZvD5AX
s78v5YMfEHs84zg0/wEEPTUYv9irLpjt+uk9OhRIfLL07v22Xu2xnBkcpA4MhPlgUSx+JU2Ilwd5
q/B0Hr0XfkPE5OvQBSReUxIM2af22D9kRFyE8OOL8KkdHlKK1lAVjQUk29gz0bQFMrjMIHPjl/cF
99SEr7tALDpdS3Gmw5EDOQeEo/WbjilZVHlUTpDkOwt35eABS2SPb0CMoZBpj9fAfnVF1g/N0Nwu
Y4kfSk7JqtTDfnkIGBChMWcz2TqzBGGYvK2RhZX0+JcZT9JLx7gXFlK0JrtLJ9R4aXxkd6JyGr3g
d8AiG0J1VidS6H4MSrASVechmRfn91vA3BLcmuzBT3lqj+h2GTUDa55DR/AQv/mQ/aH3Mu+pfntF
+eFrfM+khgMX9T+dt56TB1uYN71dz/jUFcgHytUCnvUs/BcRQDeTlWtq16DSWdAhrKUN7Vm7j0/t
eKdqvjvMilrdqMsUfx2ttUs5V8bTa/vXaLAToLNY+6h4EqPFrN4PuQ/NUHU4ZQLfwsMeUORd2b3S
GTvuM5NmozV7sJRkIsZe0CgaBlLgGfMArwJGiogoHXhjaE6wmyLwu2JSF61oFOWzYcwLWBhXQq8Z
/8wx5h8rhyLzTxnPW64QG22Yn04yff8B6tQ/dZqGENz+n6ZKZ6qKma42EL5I8jh1ILi2kTRc4iBf
BlOCylK4D0RU7PjVTPBAJXRvj9eamY1f+XQ90xveRUuHI53SBZvamec6V+akhmNU9Ljb+MKzQ7xk
28pgaGwmefz92CCFFR8jkQGt7emCR5SwT8akiUfEpTWz0jNyNJSWDZR+iWG2MBVHaKYnT+JrGe7o
7+F2flGjIBCTGtGLyRr4ERIoSo4EPx1ztrpTzYBTnnoZ5msAg0062hndwXr2Q9uDfmFTDIxbLtlh
IRLsF3nKLz779E1pwEWrF4j0+bSW7jB7dlH2+PeRRm656m/QiyZTB2xKQUviPoVfHblxAG0RdGhV
7YIbOlRociNPn3BJ1aLVV4Y+qLjIdc2FWuffouFgxjolhVV1X1B82yKaqxkH7XNjhMEbnhMJOf/O
cVqgSLifGrehoqBfMX4aRfI2ZbpeodOerQhzZNZAddG3dORIo7olgX918Z73BN7DBqapSmqJF9eJ
OSrZQBw/XMWBfAUk+YDR+5fi4NQVIKmddPBczK+/FCCag3U3+xRwajCY7kpV51AY2gOUkcNsnG41
/qQqx1E4kHXpKRNTQ0Cr4Cjkw4t9OlsyQ8TIPREV6l5q0sD0GoSGMYzBiYC+knCLosZJ0aQz5Iey
4C22QWC0ntAorXhwKy6KwUCxDaKiY5kqI7d7N4SNue6vsCzRdbrHNuxgyopIHCyo5XaSeMRMIlvf
ipdtautpHdDOrpXMWACAAFSjXi1rGKuQZ5LfKJdFMCT97/uwJBFpPQvYy2ymD8GE7o/HiJus/AvT
iCdjbbKrqZTPPs8tgLCWdOqMLIPZqV45lmklEIPIrv/f5BlvW/gtoRlclU2DGJiXKD+EKtPSQSRP
q/lgn6/W/kD/4IpxU59GyXDdFBqpVmodu4anqYmt/+xvvVqG7g5eco1m9l+l3G+49+r+hTfide1J
9G6fbOmdDhI7H5I5a7L8ivdtGGZmEU3XlLGeUlrQede1a3RVK3tHWDfaByCmogo9Qbn5Gti8hYMc
AU3QZak6s8FUh+B8VCNg3L4opoo2EINokT10WYLNWcSc8NBABtvX2PPdOcwKBShzXSKcvBr2v8Sv
HwUwPYoDfY/acvtD+sZa2GMHJhd9+WRG+OUW+sEj7NjDELYNqfSUlxLva00meCTVCalhLyofRWi/
BtWjc6tNUolICbkZy/aHIP/XyHR0Aug3/5NPFfPy+2T+ShvAiJJibmjhTnJTS/RUIr4AydXS45+I
aRRug0QQst/TVyr51uUthr9ZV3C77jMMUWdZEun0mgY8IHV17t3B+I3J4ys0AgyV6Pv9yJ3vlJxH
AJwGNyVxtMXmysmJCuLL80ugr8LrrDnJkqI27WoWIYrQuMGAULfKLJoAY1z+og54N6uk2livm2Im
SpUreB6CWe2vPtmYhD8+HRVaaQGuTG/zfw/xeT7KuoX6cCP+IxPKEq8Tb5cQvtgmqUO0uk/yYatF
BB2lSoiOkoDzhMYJs6IcCFG3Tf25Bvrn9PrqZc9tuumNw5tZAOAifC25Wd4L9Rhkr0CeXFBOBSBr
Y3vBxogFoiNqpMBnDHOdLPCPDCqPeiLtN0phQ7VstlS0emjPMa/k/P3Ua+GFj6j+z0zauOSyoH3H
ZTuHEN9u6DGdPcmpTxGtKv43cDJG+bzTPP3cC+yfD4gVReS2MB1IzWx+eltOz8EJUTsGDliINks9
90Rc/PWjX7MrPp1cQ/+bXiGH14cSf2wpMS3g8JFae3vnb6AfbDjYNuTDVjvDUv3JwUrigFfgtWsF
mcgClwW5KuY2VpgHgCm4Cmlg07v80ilb519XIrBipP9iP6B2F/9Y0gBiVY7U0P+ud5i8PFjTklyI
ccG0or+vqiYrXDuoGsNsfE+a6wBNHtRCaPqf6h9/k/8tKb03nF3xOSlmRoF8Yxel+kAHR9wj1rCx
yEAHAf0nS6ZR17AwlvZ/D0NR+wbTFN8mpKdjM2s5PWl8t7YL9U1R2Xohc6ArHqd+QNWy+d1hYzak
+wwVkv8ZTOhkkIxhz6LXtwh0Lwf+Ez64+rNqEH6B0G5GLxp/2BiWONp/Yq4Ip8JeDJpyhOqM3Wg7
LGW82uC6Hvjpi3IxqzEajbLh4rqbolUYznf76RkMoF+gNM+oLYOGEdQE18BjROw9tFwzDT5Luot1
icCLSvF+EsRFxB2dx9aqV9CT6Ffx4j7lEcMNsjt6UK7J4oY95Uyrewu19gpHyXOAGa303Ze0zYnX
mCBrOQn0FqkGKt4Vwye+X3bnwrdXdZLOwYuQzmbG41j4Qf699Kz55rFlni1bdqGoTyG054ZacMsx
gGTrRFgqEyhIqvWTb9m8/qs5LNc9LmrWAyagH/qgl9C/OgyyEMXW7L4vcrJ1RCPllYobRSF8JgjN
tHAVR3SK4/IjYITpDbQaNhZZ16Wc/pFeZobnH1lJUJDZUD5lXlW+EJZGc2b7+HTgaxSMguuSa6um
u8Rj+TKaV5xUydmueDDm7ItJ3VCVF3RqVCN0LTjpmgPX+PT4P7zodFOrgAKl8tNLqiwUAlK/DJyg
B6w/kLg6QgXRwdQxNDv9GuI5BySKE/7aoUsH7zqvVcOxtXbvQjArUykmFn2qyZHq8ovkwXz112cY
OyuaHvSe0ODSrPHD1ouIqgcElaeazRNWOT9YqJA5lQFudJ25DUlxNHYs42aPD4Gum7azPNH1nj7G
15UF36L2JXsRHqgRhwd5pGKtwgR4DSK+zukZBpH5Vddn1ONqVdIAsmXhwCmtdTVUm+NoJS8n5mcH
FYO9WDHKMV7uM//duHHub3vNLAM5E1qMKJb6Mnd4KDxcVQPHPNW11evy5pDm3FJRSQuB60PYxraL
R5AehEKuZt2un8RoO15102PY3t43yqrqRzGwrgysUYHFUuLtTJDqS3Woyrj1G5nroCnq6JpfbU5e
JeFrBbPbx6yGMO1HmKdi/mML6qJ3VnNyW6yidaoY5xj3O50HEYWCQhy1yCVxm4J13GuwCvjH2AJY
3RUC/OtT5yog+U/br4vpZGF6sDQp/eZwvTWo2pMO2owGDqG0AAtNPvfnG3rOzvjuJsYWC6L/yjJX
HV/fJu5CLJN/RHRBsh3NWIa0zCZwytH2dz/oD5N23/ZOLBl20J0a0/qycmVYQmCP3Dxlget/g7Hj
nDB26Ff+cgojz7kts+yHZjO7+18GNz3hEU+kImW+VknwvgwcUIedcPQfe4Uh9CQ1MQin/bYBYhNT
86RklxvpUh/gGdmiwLAY3jHT4PA7aViY/nHxydwZ/yo5VkLRgAkGvRv6yOQQPGdtcvBCdmU3p60A
rFBG8HETg5AVCfJg236rABiabR8CGkeR+Thtt3i8ASxKmYMxKDIeaN1hDw/L/2Ras3L8+tCrwBeC
aed7rJpwKV9JTdP0Xq4TSGXJJ6ILbQJV1w8RzqLPe4iXtWYqAQS4Gga0T6GEnSC1SwTjSee5WpMx
ECmeme9o40A3qh2u/m4lTfFXtnxzmvd4AZN450hJoAuOuEh/W+R1E3ZflrcabWHMvxGB5VNOGk8q
VBUOiblW7fa2jIUwI91yPLeGkuuYBSvrLZl8UM4gjJnGuPwsqsyNo1nw/P4AM1A2h59fyUuWVZmi
jpHPp7/Lvv+F+w1jXeosMnzd/Y4rsyf/PDr2VZVio0dhHOFaNXmksQlVgMp3SQSSdunobrS+Ta/Z
Rq17ZEeFOM2oPBPYlw1s+mQ5LXBfsQV82CWp+Le/nXMD8KFKt4LELlrZV8fkq2K2IwmrJUybCDkX
PMHS7Dk1Sz/4w0wNMtqSl4x4hEPotyzqVExd3I990ewIPHOIif/Qc4qX4HfU/6GAMCF/evvpUUV5
xBhsA5mKnCM62sK9ahoCBJOSDZcxZRMlg+S+z9IlVLbwaPjzt48jRDpX4FMzjsk5mRRIlr2wsgYx
23jh96hiFufOqBDryoXpsdNGDM2C0JEEJPC1GfZ9pFXo+acho1cX5Yj+44xUO1utVkITAVlCiGaL
g5+MOL39/xOeRPZUdhy+KAtnTf1Yn6q/rAtAzkCeBDQd9hRnNV1xlfsZReqfkdhsLXkF9DDfJ+t4
cd8OJSt5MKrGwiO0ugE6FMZZeSxGtAaRtulhmLYycy9YM9ums6jurIYmBEwAgrk94A1Qy2fM3Qqr
3NcXUm77qFKkxJcsVCkklO34Cwc0g+NaiEwA1gkhvDDClHVqyDOB/8pP8t6Dx9+uktbO7BuXmRPV
0/u3O07URfyZtwbgb/LzkdekJUSRu8IIgtJoT5tjudLKdsGgmU3AtOPk9phnYAfmiEEVsekhGugt
LZChpOJPLjhTS0przlrKREHTK+b87n0pgv9Poxzab8HyjazLFi7WnDWQPZeeQqMXw3JxlBE3GFqo
zFE9h3l2JxtDL330K1bHLZO6vRYJO/eaQF8gtT0tfgzmnlyWWcQz6lS7zCB/2PDUc4mHLAuJFvY6
nZlpHme2+wCw10fvLyS8yYrPF8RdA0XRVAB5Q8v46VHZDZO7hfob1GtylyVRWXL0mcWoaA0bqNcv
flRUdS8saCmIesfwpZJxWUmqXGBgnRHd6yLQ4N64iqK9MPsFG5U7nctNE6Myf6e8qrSUMoROzV+/
yzl3mYUE1F7vDitBNPokBYoNqNKpdML5zZSANX4s688BnGvMuMP8J+Q9ILDHWtYmh7nrczfekwgS
fO++eOY3GhYSA9littF2MpDhbVtnxytJ81RkWCdU6Q76OZPnFXtHQ3pu0Fr+Ym00FNYkYcGoKjBe
CzcfDZw3/jPVWq3sZvGPQJCB4yjVLRzGYn/IqIv3n+LAh8QoRPp29YG6ojXVLZ1mxH7XYH/6CN6Y
0q7Fa5l/4GP9xr3iAzUXqMCnOQs1BYG4nlrMnuEXpG+tJcqz6QAVCX2mIJW50d/38dRt2yCcZ2Hi
cqlycvHF1T68jY1ej/wRL0XL5i7o0v+zDQsTjB4GgdhRattl0coDQfhkT65qVPhvp3A3FTgImCeP
AinCdkLPW6NMfrr8eJeqKNsNwwCGfKzRMJ9mkQJ61GRnKudv1k50vm+IudQId55ErxVL37vGV253
33Eyp+7IpwuWNeOxS45V20K1TulBQimgiweko0qb3MpMt3JH8FBsIgPt/qQxck6smLRJqmjkWXIY
obQA1Sm9zVg+OF1SVO2nW0CIOcuKrwvkAfMmny7nToKXU7DtpACkk9IoXSsstsiGnVP7gmfdAz0l
wWX3OQl8gKdsPy7UAim4Nyhw9Wy8HIedTeL3UJrkmKmrebmuLkKIThpcNkZHqzBeozKNE8oWyZSf
vO2vmlhfyFfSsSYU41ZfUXLvBSXWL1xaKVbSY2jRpS9MLjep4IFNLdTdf1gKo/EnKgkEaxCpYysy
s6YqWjd2mOicgsSaQXyo6cP9JL0FPd2hNXZCSFyQ7xLoMlCIHEraB2ON9VL9k0hqOzsJAL1fMyx5
W3ZbEMj49bLRJEaHbjuL0AHIjg9ehUS3BBDMnFdyiYQtrVNcipRWqYl7vzWTy5yRT6WdUUs01Dum
FLX3xc8BERskLzUNjE2TpOSiUG0VQI83iKv1s0aYETdurVWoc/2JWb/bxv5+ZyEtlkYOG1pQYb+L
Qw8gIxvq0Op5SZC/PsfiMsoI7vSirtVceO26yLNR5HR2cRfVBtpcPs87F1JUwUcAuCSkV7+9WDyE
WujOfOPfPxtOztyMs1phfBVPqRY8PR+kU2HxF9tHEGhQ1D+hAUhFEPddByE7v+Wz7ZWgYZcX+Kgr
mHFvtuE7QluWTe5/Vo0p8HWWgpT26moA6RkmYaxItl2AifXo+b2S4wtOElGKasP/q22p9+AKYR8q
ygiozIKpci929T0LpQ7oUqRY0JrgARcJZJCkiUT5KKqz/2xqgABgI/a+RjI+C+kR8nA4JZ5kyntv
CgeMEEbpEyvVzd4z3qPYE4VXHLp+fQo9mqesGGh++X3y6zXPDRVMbattj4MVl4MW0BQJZLHo7ODY
As62gGRew9K0WUQr95keVuAe0yUUbfM5HuDMUwFduJ5yNVQbplIzTzafygE2I+Z+2J3F31ouch4A
iKSq+FTgVrdqQuRp+2UXmeBkp9SbEBK/YZmkYIQXOFL7C/YiDUah8wxGux5ii6C2B9askECrgWAz
M5L+GoLanMH/L+zDudDKlU8fi9pkHsXSxZEpjHbSoW39ZiSTMkvQAETR5XI9AteDMwuLu5NOpMl+
q9VRk0q/NBAgnSFuXBbI7N4FAEdAJ5g+OlZGP3T1Ge5kO0DYz+cmDjJPMtdPqweNyk0HrPKZ5o6x
EBHuSDRJShJhDP2KRonXKNa+99MfrN+FoUMtHiTeTn8GzcrzSXJf+ZymsudZUK6NQahJzzcjjkjN
f0xr3Y3TUnEdCQqXA6GcXA/O2I/AgT1DsMhrPJ86CD0CwAhOyMa9dkwiDue+8vFgpDfPhRUZZjTu
u0LpROwYrly2kr1SwPqjKgeBzPA1E+f1NA1tZjbJ4dfnUmgtNoBWO+4bCG6FbSroeBOV5nxI6z7G
x7Mt+C2xywY4WSnoObJxDeEF80aHu8KfBJp3Z86yIzcNTMB5Zc/lHCG20aTA64iKYDjWbfILOQ2p
+46vQSEz9qYwA/SN39EQB51oS2seHtVPS1S/8xcE07987ETiArDpjs9xgBq27JBePmjZLCV8Anqm
sjyj2JCZA/WmfJpNtBHef0nEyhi483ci5zTKyRUq5dJ3uT6y0ZZJOhW9JwdYuu029YbN/p5Vypxv
oCJS7UaKRNuB0zqNX7WYywJ5L9vqx52FXi1Vx0bMFO+EIVjIYsZrxTem+sh4NBY0Xbsc9Ruc468z
ZRTr+jE8HmWG4HnTIEs6OqLIlw5DEIjq/aIC0hZgCAQCDadIoH9jqT2yw1QPZdCIfnj2eKbfV4sh
WsKXsHGRSA1e3xChAjt/iV6BGgBpoJqx86f5UwFku4wct1/Di1GcM85cLwSMPD37GJ2PMOoTzlMV
qiR7SSnZa+5YFmYlIVRKYrOGelBUQc96giLGkId4Y47iCAqPQtXO+KDVUcxubOxlOIsZzdzu+6Db
yjslkvUHD8QVGS9XanBwAaiyFXQm4E/okKeKFGIdZtnD+JsZufIzDkLMz+c+KwNpcgr9bxjnfJep
cFnNn3wW+TgC2QZC9+UaMV80xFQI4kjgbyX61olD1yvjCOgRN/V8rqdVOzgObQzwTYF9VA4YWnu/
GQYb2QGNNr7JkoDf5Ce0hjyBDFGZKPhCmFHQ4LtNdMY0dXZZvVjgpR46Re2w5F2rd+mVdF3U2h7p
N58VXdEKdu0Cfa5XkXWLbwiiqgEiM4nU0TdeVKDm2fbh13zLPTtrHg/hNrL/Ehvjq6TeEWdyXZb8
H3rUZhYKh1Eu2/jxeu2SNzu93+qTm/FcOOrWXhgtrb7OrPZO72L8mQxFQb38bUSpOV38Hdq4DIv9
wB12b3HTmVH9u+YwM8ZYlF0QG6K8LPcjFU1wRqdBkTi/ENtYpXWexTknFn4c9wdZc97n1NbOa+R7
oWMMEgcsETCTjtBRXzKEw187Bt2NeLfilCkp1cCwxJQD1sOePILkt3XE0y8xIQU4dbxgAdhAYasL
WYIt3/wm811+hfSCdPZ+6Lv3Sqc1C7lyOh/zu6tLADtmiTp+xkV3wGKCPBDI8IAu0PwaByKUEtMl
DOAaS6OT67VHuFR/0msJnroYgYSH7YlNRqMhGzDLqZUDKfK1FmUsLYNxtR10OHqc9nOrNhmqemwT
Dw8eq8EsuYCJVVRo6/re0zIOHHWnZy22MqcqgAC9hUr06WfgdgsaTsJcPSm4UyprFRC5doeFX2Jd
vL60s6wRIF8eet2PylkPTajrChfQBaqIQovqdB5/P0rqG3NDMbAyafMt30Y2UAs9hGfcBwLTi9E2
7Q8bfyvUdP6NDyIbf0pL9SpvghBOYSsTFsf+ME+4bMOBX+27WK6omu5/b76tbAMaV6CmfIVRcYge
3Fq7MGI/9bZCvNZgkVd32EMkZWQMwdrPDY9GDwp6DBWBIZO5mq3dLeBKj6WTAbNtLbBWEd8aGA6b
xwxLHGkcyeyCeQH8/Zuli85piSxTP/eDSyUqQ6qBfyYtjK3xFg+sgs8TkU8R4pI/MU6TMVetrIk0
ikBU5WVBJMeZYQoWFpkzjuDy2+AfA5ffTbTW3Urhp7CLiM3mPWIOC1XctdV6ge894YXupZ9l3U9d
9+SgaZK5jQ5cDJ9bocvrXheoS9UbSN2hRG43pnCAsSnijpCesMobFoCdxjMuM3H2mW16Yw3oA8OU
sQmqyqY7x9NEr3o1eS4BmwUG2bzozx91owtexNbYTBoKHedojW1+TPFohtWvMDc70+8/80JgYQxH
mtUpoTRFZ4ZXQFe47O360sZlUkJ3u5NANoL4EdrQOZYs/KQkkdRxDwnCtya1NPagiFhnIKLaou57
EZeA9yts83U/cw/QnClJq+HHyV+z0rZLt7CN8lplvC3okvibhKvuzW4n1XVvYY1duV5+KCqNFWmz
TMUqfsYa6OE2Pqh54K8Gbb1gEeugnJ2PfxzD7HDYDK6RptziaOIlo1+zcKccEV4l64jdxvE0ix2P
o4/Bh0itwm2hR9LwcHy+RuU4d1Bfxl8lCa69G4r8df3vLD16B8XxcJwB7VKitErhYlbRmiuuXX3b
ifdn6e/kkq01r2vyWuErx/vIYgGG4Knnh0WA118Wb0rLxPji/Xieeq1GeMDtCT4MTal/kB6bfqXa
o7Zk/FZklB/pEBSgu8IrxDJ4vU8msPo9T+KFeJqpJwGgbupYh0bhk6WIVrrDhncv+R61reMk6v/w
XG/0D1+8thJrlHiIqX1fsukQnOOTTF4oOq1P0b46FwKQFaUABjmde0MuD5M1XKqSeKnhqWinjJys
493WXRycuE0TTEm0YFExTEYBc7t78q0gZipUeT+ISRuZQWIgHl2IL52Uzy6ohWUzynYeljzSboIu
Mrbg0AhfNJkflIGVlseKOcLsQmQhCh9xb+4DovD2YPut52iVHlTNOV0tMp9vc5Ov83SHMQdWoEXm
WU/nY0sDmsNGayehURXwBAJxmHgeL8cRkxCJ9+UUT6X5AEiV1BE1KnoJkHAOwg/lNUIaLuR9RRcu
MvpxuvADmIwSc8MI2KP1xUDDmohgX6gwe7rqf708AOtsg+2tcN7sB7j6e4KJHYv/5RXozXJnDFHp
azYaWCLvO7qi+Qo0njY/URcUC5Ze6TrT0iMX8lQ4iw69IfDJN1xtzH88Wpa+BK/JDNvqt+BERZIc
+jaGFnI4zmT0mNTh3urxtgY39lqvOffdXcKSqZ8evfy1JUGhubYUzh5xiUe0Sbg2GzUDbBc7fB2f
HgFq3pj5L4q1Lkm6O0M1TWp1qgBO4SlojtQsNF2ziky6i/7d0X/lWAQBq3tHqJSRSDZbFEUE/AHl
HcDkIJQBwg6zQXAeXvh0xyASxMnc87j/qBNuM6VKM+PfoGk3PpBaRjAkoyMt9vGg9njLTgVB2qBI
CfIL8GW6xpbGKwtbTSR0HaecQ5W7pjRZIDzxov2i6i2Vysi5tIrjKxidTNdX+C6szgldvzvZ5Yst
u6tcX065a1stjORXImH/nXamx9JvXG58kCbPl53xa+e+E84HxTNY1S9IR7SAG408XAIjk5ntvfNN
5DeZZ3AqsHYjgWLEo0+lamnI5g8hGQ5yWuBV+CewIutS67zpUbUcwq0K90d0qFypk56ZXgz8ybWV
2yQHYYEhKQy0tIwOe2Mx7RWZN3JNffNSvsd8QzIaszofNxZZRybnn2N85MY9UMC//NUJhP0/tYNH
xoJf9ZWhtYMHdXn2xrfrEE/eRW4ncKYXVNhUvocai7A08vkelZnPGAXcde+VWIGI9fxJXgejHZpE
Z7e5p/79WfKib1M7UKMUAbDrGofDZCAZPxGV0udgpvL5cebVANJR3PzUpAkmZLUxfdGRtsN7XRm5
jruxnC4+g1X/qck1+irPzxr+LDIzWfRcber3ZLePVT5mQlnaPMO3VtJ4SpJEuSg+ynfW3Cay2cli
Ab81f6HZpNtK1WgDboJ2hIw4n3Y1qkhE5Qjfo+ijzEZ6R5w5U6D3DtptHmDfzkugnq5bfvrjDSim
mvehVY7ta+6/Dr92UvvZkEKNGgEKZ6QZ2LzsQLRia/1Xd1twrGPQAGYwub4OoYCIlNcVOzY9/Efz
w9W5rcMiigqrpd882xrBYZuvpyNKBnZAwG56Yp88cQ3/5vPIXXiPCjb1EgmZ5enwLo8MKBjO3A3v
VRtXR482XU4a7HbK69ifFctcJfDayOHgs9qYIY8cn2Kytvl8Y0kTVY34PxGwFtMcS367hZ74YO5n
Q0J8V/ya9EgbfZDCVJAfBiwXlK9R+LsCKeaalweFUYpusnUKcVXUg7pU7r/AE9b17tHUH8WRABui
+rt73SXCHeUj7KUR1OGivjaj0FApJqEMv1yA+gQzTo1wVzRzCFejkX+VHwQjFdk61DOuYZa8C+5+
30N9zyywy7x7FZe4jP0Z61epJ4DoXjc8MVsTTLZyvVPFGKXyTxnMlz9WKyHNG3bz6yLfqhfcy3AR
+SoXYMRxpGFQgj1ytiXDDBuEEon/X9TWqJxCVdPeabCul1FmN3zlFkmjeyWQCQLTeI7cU6DsB2Sa
a0V076KmFhk4FzteXDqVActmm1jhABKuf2dmSZSH669B0v1cLMnovmmTSdyrv+wHGRKWnJlVhCjV
J5M/WCb7cFEeN4OKL5I8I7L4Njtn447Yr1jguvwFHDFW8Hba80mfNpfvxq5At5v18iNkQbD7tQlG
r5FEgeCJwgIsdO9yxzb5heYG9qe5tjpdtV+nIGIaXhhEh8VAT7OHynkM7eusRbvXwLdRF3UkqA6P
dRUsY7222f6ZRk13b9XopSMyKRiSejPOUuofR/mjDh1APDNh1ZZF/yUZChyYCVApbJ8yFVLrO9VU
Qk8YL4nr8Ov+4u8p8tg62jhT8jA6aIucE95jmJgUZRWWAT38/SN9VFrGXGysXahPAHHJ7z+4qqSc
ee7mSfnZ1cBn5O35xHu/d/viGFlz8uvmCrcDyn4sj1PyNLCbtbMPHSvVlOdGOfn/4Iw0XY6D3E7+
vhTc8dqTHaIJ8/vxWl4IlwWwaXVcCwY8vnW6aaaqhtxdOWqf6vLf020WvXM4Po2rcp44VeVlegVc
Er8EWP63CQI5LZO8p8f7C3y6EUDCmlKS4INeTW9esm487AlisD10/LPTvS2B1xedGr80/rSt+Q6w
cFsdbPSDpfTKga3757eQ59X5e5HtHG3ypr9K0zyU28ZJN4S1vrK6KfRsnpdE6Ok6y3zaoJVpSFcC
X/OtVnXOMjmx0EtFOQMbUiQkD0kz1RfRm1zx6zTvfUEXCIIut5n7iV8e9EJlOLdWqsYnaTqKio+b
M1q5lLBhCrSwFVdGEOZ5k/D4PQs3K+EHhFSGOwTepc2Ohm5T6Q242tdtAq4Gx3xab1wkq5tAMzh8
hZ8V36Q0pw5RmqdWsDIXTQn1jbMdx0hrmDD0eklqkxrqfFoteug2+NqcK7RKKT7w3ycHI/R0ZLbz
wP0lh4d+iF4Kjnp016wDPKL2BxFGM2LgyqeqZ/mQEPxw9zkprn8NDP+vsCWtYirdc9ROPaOTkwRa
jBhRF6KBcAWQcsG1OHF4QVrEJ82UB1yBpLnnFHhOG4kSesxuwZWG09utoS16oQlEy8F9IFm4rVv+
9zJyzBBP4XkGypem60E08NAxrZdu0EAPyVTy8OqG9EBfKXJid1xOv60aMbmTDSz9Y5Yl5wJJ4+D+
qr1/g9suIPdA2A4FxeVVcUFVJD0VtaZXuSiknWb4MDfx6W/CBC8Hh+249kvPFvMefCxpYW2EcHhk
te9sEt20RWsxTZp3XJq//Urt96R4/1sDVkKbW9qogE/cq1ytfSZblGMQYUyH6gS8WENhKWgEtzjU
Upnya+8vcw5/jrl2amctedoiLnkqBO2bM1Bo3rRXv1Rd9pwut3zPtHd2S/VWLf75UvYuDT5UIvvs
NbkKERDEOzFUeTa4Elts8yUblx2udZhLZj1+sxRElGOCPj6ou2/5shx3rbZE6VfO97rh9k7HL6bn
7sgDV9f8+i6y9nTQ2hd2dUq5tP2ImqqxNaeJkAjLFtEfKkdTK/pKJFQ/JU1HOn1c6kkOg0AeAfUO
IhKPE1qsyz1NoGKer4qFXPzUFms5Aqn0bI1v1Brb8DCMxHyIF/qwnzXsFKSxyfN+EkOfOQ62eeMh
y5vpUh09X0mnFRAE3OC//BBAmtVdueGadzEZGrzUlh90I26y60RnuEtJXnYyq8Tiu+xInSSxYxgn
IE6tnz8rqLn1d0eQaGecYcBaBAZ9DIIG26cUVpvG39de5F5yLeszEg8tYt/+51KmRglZ1/FvALS6
PSoqvnEKi1amAud9FplQrPO++HZcTp8EMvoFRvEpkFY3DxJEgYgSwYP4IY9/iuhReMV9lugJHUio
/WwmsiHWzTEN4rufe5sbbMYDAPSuMoA38q9F5o4WCvgiY7fEbla72Gdoe5oPEMkFD0DibuXOyI+1
eS8xETTGJMn9vZihAzySbB1DlwpidShZ4jAgJqXMF73erL3TKA50/79zaQZJFCE1tfF+I7zDEUvO
+2jrk7Aek6MT3Q4kPHkb/8POHUuNNMf9rj8rOFByi15Y2UYDFrsF/FmCdAnmy6D2guTPOVl6eYnG
0Ye1IyPd8xPhEDntX57p/D/isVYBeKJ5k53LH4WA7rJGUcXGLgN75q4vn+slB0R5/BtXNjqMjuCj
QGwBeeVywJObw5boome+oEFjlYqk/f/amQa1mXWpACg/Gj2TGO1xQHJBf3Ng9bzeqndt+lG6LTOn
Fl7y486Dw6lFQrtSjGPcrRTXIYkNtDravzIvt0hAsZ0yEYJm5JSNbRXBQoJl/GmHLFsmHOIAjg85
wdHvcIpqHPUv4xy/hqgntXydpZNLS3P6Pv6BDmLG+/7UHrRGZ5h3lz5McNLn1PjCWPQp0ZFBjfvl
oIn3kISgOtvxcctnUB+HwGhSOZ+NlGBh6QjX76q2keYXTVmJcExgltO7u8J6zxyTC+8piFPCKtTy
eekZN+OgppIYDvdvhHk8Y25n02C3e8pwi7HXq9BH7YsfA+Ocq93RLzYpd0OiAPP9E8LvzKnYj5JT
F2fp+i0Dj5zFJ5FAqMjgrm8oQVhgH4BLf1SaS93NcGLF8yxWoiiINRBkwrNNnGQcUaHu/4j9B/SM
n5gwLogxLoXMxifEIo/JdMPrpNPg+XQFgs0fMYzV9PLHkXw9RRzMLfWa6pH4GFl90LeY+RYH+auv
eoNFoYZbpoNBkJPHLjYGNFQgv6D9pmPU/vNVUeI1/uOganTGWeuzNl1BBJ3r47xvYqYzudvckIMy
X+6fpyR+kFC8RCRlL0462aXKHfrRoNIXQwPGCJda6dNDBOeSaLjqm8lYR+cskm+82q2JZUDRahlD
H0i4un/djJPYeUlN3tYSI4GtXDVdGeqSZ0zW320YPCe1AM7URhMLStwvHbJ2XEAodbWORJDP5VRt
UDr6uFqmgCBXG1P51dD5dyjAWsUSBolxTzvWpTRvadq8+wXPyif5Y3bchFPnE3r2x+VVB/MRf2BA
MGBFRloO2YVMWC2VRlQucJ7mWjX/k3L5WTU90eceiVvrt0urTsaOHwvS3vAhj2mD8cRWQFrFuPx+
suTt9igeLCiUYRuAzCpK9oTo3ICd17xBVXh6oct4rqdvRobXQzm8UT0pHJJtuD1lXFvPkcQ7pItZ
6sy24ZtTVaGekh813MhCw83Gq+lUTUhe5SbanjvS6R6JiJKF68ZO50pBI9YMPOU61QmkaXpBFmCR
xwa+LaCSW7NfgkX6d7bN1iSDlUDmGpXW4C3sts1RP8LT27wJ4CcKkEwdZzU5MDugJWucSI+qZvCb
RelFuYimBdEaYQKJdLSO3lqeHI1gStNoUwY9ecg9NKW7DjPuvMW5JO8kM0QgjmDAQnSjBZFIwFOk
Ty9GhD8ZpR+0Fbam8YBaFjlCaEQtctRc37MNLl9BhM7Rha5MVF2bQp4msXyIvz7mmikgDWzNMZ4w
Rgg7YV3UeaeSuzKGdc2WER4nCofbMkERc0hdMx2Vj+tG7FuOPStOJiEDI5MhG3rFQ1e1d0K1Z8FR
bzoKCDp2ADo6poDLHR3ohiP2BKw2YjkTHN1wBS/kJAIYcmY1/sF3eAvHIhL3zAKmxnMsOZ+5RrQ3
pxGInv3gohpczXxGA7KGZ2tJMvo88nEku5e7xZzH6ZDfb+LpgRNeQ9uVebXMbr9ci/cZYrQ3xlCu
gBj+xjW2th3f2VtAzuit+8S0lRRfpyMMJhOu2lasaCTSgA7kD1KuKqKh/Xz5Gc7itJvdxe1ufLpP
IChNci+VySTebUU0GG7uK0kskhxSwgvGDKF+zV1If+OoG4x9/QgWfmkLCkqFgE1id2DlIT7mHs+6
QOaqliw4bI+ME4eqPU/OwKL9gsjKYt93vfziteFGD5eZtKScF12iyEb3jjJus8eGfc7krlDKBhFd
HizGqK8aomHFE7I1cxXVZjLeEs8U7vMxiKV0acWr1pkjvwjAfuBqasxMvejmNO+zA5BRMMnVPUea
7jlk152X3gffCri9A6kUIvg0IH3iK0M3Klwfy9y7g7A77SfhHzp8QumvvGQFAO7ny412VYkyRfpi
7LOCqavDI3QZXLtCVYXXNmqIGdV6u7l/RvhUerN1J4SZnq+gl9rMzFcSMrGmT7nLWvpZm3bwEShx
oPgdbAdTGGHmLTmCrYlomiy3Ip4Z5YKQNlwCz7IOG+FD0xeJVFFtwBcBpgM8kCSXuJyq7hIuW7pm
EsILP/1CgaOyux4iIm7/hnJkcL9vQ4kPh642nT5a4Mnp748synIjoDw+/ytkjfGWZRbeEJe+FbXr
dVmGYECHzVcnLKfcbwRFLIFTAiJeh3qwM+ll2Z3LGhaBYtxgsLJfPnaxaefzK94HGQsMgvxCUcBr
liyHRBWwsHbK03vyRHgRpy3y6qjsZofAsLdOTpNV+5Nc+KRIl8OYH+CFJZ+WXeXYQDB9Emk/DZKa
BUGzrb6x+Pdb7WN83PgyXA0ICQm/5sZQ/IHJrcXh7hhXLYW2ZEIQXuDI4kBPmbbo7fRHnsL4ME1z
yC+QGrCleR+N0zdA9QfPe/+XGJAkjVVwarakfALCYxUFxeFdN4uzLKzuA5syrT3EufzsteRCDXy3
vcHxNytL84ac+ljiZoCZ0yzguxFeMHU6S6Q37Gfj41r/MTSO9nugna/Orkfz5Mo7+Hcqyxp4GWvl
D8pVsfPzpx1mm1R0CtXP/4uwy1mkNXtSJtZNhVVscBkxP4ML8JjwAfXY/KnQjYu50ONWRx2ywz1w
trnC+CPHPSm7PUO6d3VbNazgFseEFWSR/m6R6J4EDlZg6LTXO4s4Hzoq1Ba2CsGxTjviGySR1e19
zuRPoFkKe68gJ1gSm3yInLU4xI+mq+EiP/DVvpMzzXT//FQOc5LRh1HSqWYaSSIvhPJqoasa62ul
ISyjNrvwKDE71goa2ZnXZpPc4z+jNIL8quT9ifz6wiO34dnAUh1VyG+G9Z1ffnoUhh3Fxu6VPA/+
aw04A9+XjzoE0iyxO35BHqhbsfcpCr+AQjg/qleoIaOU9hO65sheNikCULN7K86SA2Gq4cxSPP7a
zZRdS+ssPnA5TlipdCBbeUiW3hsdcAuCKQkHA5usL3p/uBB3McxUoQq2Jhnyk3V4HiReSE2ZvZqM
/BRJ19YXBZ6nvfSFSsOP+x2a+mcum/gzlp3sCNN8F8BLVYNGnyyEQW0VZUXuErVvs2M7Be/AaN+/
XpYUbWCYY8a44aNOS/5Lwhl8IDu8SjFtLd0igxpoUxAbn2z0sFsBUk9sn64aIH9ZXTPhHYMmb3rm
6D9XU/j+jf/WP7bjM9vwJ/ROuErmxG/Cuhpy6yH1vZZ4h8Norh152pBpUgqGipw2osZHM2t82mUA
zUX0d9ELJ2ckrjQW7Cp9sD16WZ1ewVwf3xBzMVHmUvWDjllEc2d+8LBNeUMfGspR8O17j/mqZJT/
25MB2Bnu17/UpYRNj4hNBTfUZc7M/S8vt5q6gT05842IkMLEsw4PKErm3BrwOMkDHTjBTGYOjeTW
hMQ2xURF1nbbYlnnMNSHxLHny1txmkPrwcIVHDP3oP5brP8kJubNR1RmP0G1ZCojeRDMOjY48szU
EQWOUvjEK+napw0wGpFba8iuSelAus2gFSKBX1tLi8xA/PFXoYtOEcAxxsHlk4g62XFVIqcyCUiE
s2+hWC4sJujaC9fkImGSOMdGeqfozXx69GPFXZ5bMPwvFA4MVNYhfop10fyz6Gy8blFbgUZi3WeN
xRrYFSGx2XaboO3d3cqcP8InU0iP+ARjX+oaEnKdZypltFj1rZ2hTNBz+MlZNJSCcky4vmfDSYlz
AldUlG/T+1ohhhf8ibRmLLecrstHc6y/bRuMjCcfFq1QhVoIuKPsTqCXSmaZOO/bmI2lyZx1Kfik
hxDGSXMZH3P+PacUWtvWNsYzoXNjg9YxsEZv3Z6PowNDSOM4ESUdg578g3TMuaAe3U7i4QnYkE3+
+2DSGXgbLObcBD41QqKXGZc0fRtKF89pu8jf56MMAfNjZwiO8E7Ug77/9hZJbRzvgXJR792vzfm8
QVNmPXOV8yG0Qt7lVvLcLXWJC3l9vm2VbbQYalA63iv9UvkjcSbDUh18/+lGmFwxSQUmidpDbG4f
s3Hlc70CMKgGRsKGm2qGjZRYI0omvhs4UJjPsETMurpFGtaRYdrUwxTv/QHdh/VKwPEVb0P7Y3ex
UBV3OlcG/F68z6HZDlVdtdg7aG3CA0eQBBLtDRj4HIqbfLNYH73itvd5H0BBQIh15hCLVmEY9NCb
JhBqV8NkyOIYQBV9hCofzoSffTaJCb+kpl5L8DS50QKyji/0+QYw/mb7OMfDA2S+xkF3EakZsosQ
5rh4EnOlq3gb90D8Zrp5plNx8s6QVyjx9yiSBJWwK/rTQvm3TLbyeYvmH5+7e/oVay2yBk+whM3Q
a0QSweql8SBktuyngCIANUblJaVFKSJFDYBi31nXUxXBZmkLUr9EEiJPWFyz2Rfj+RSEYLKaC30F
y+5wsTk1/vtv4Z7KMJApWozpkInYvJF/aK9k/gglIJq4faxl0Xmav7+0n8J7CdMidNyGaq7yEXPR
Fc8p0v+w0KTCeULbzRUNa+wroSv0BS0kfqVjI9/LN1UVF5LM2nkAVGtvyWEqjHSDAsrV+uHO9Up0
M7r+L/Sa5r0tF0PmAqlAlleYrzmf71shL3MeWndgHjr/3ATVR2J4eihid35MjVDxQlsmQCcvozkT
aRJ4T/cwHFsl7FeR/4g/tRbVH1S9jl98AMgtp1gxrF91t/xJKBAQRljAy1Fk1b+A+I5kFr8Qf1Yn
EVyr5KhPvWu8taDOgr+YITcdTKub06tGuNoE2sngPRLeaB6LiimxbcERj2rUYWSqDPk8wEkwHXvn
tXsB0MSJB+c1m9HkzGle8OD2ahX+bcR+ehvKPe/zkJx6cLnnm45PSef8qZiLxrjZYSISq8LodBHz
d5QlGdFKAKl3I32go49jPzQv1hi0MJd+Y1IZMNVXxCihYhw7Pw/UlCCnZg1Qs2G9edPFzqTiOIiG
V58QfTJlmNiw0IGA2H5WmEWkC0pyHFJ6TYmtYUiD/21X2aT/ZVbN0YU8dCbYmDrSrCY+knhvdLXZ
zmDtIwbuQcZZ/k4i39C4rLyeToSf5qUHT8yycfnJOqNVBbH/V2LK9ykBtOjAm+gskayFumsoqidN
ScL/7ecJv5q/HfDNWdNqVKVB06Y0axOX6o3EMLmqDUVwu66EKmA17sxue3rPSAo+kV1kYza4Zaii
D4Nw4t9WIJvxXxKhZXeEgeJqS3sLrBw2rScxTZxcZsTgWF0ZP0sLn/3RJG/5fISjx58GI5PUIrjS
sQDhGej1djxwyCTjbpsIoXZQe+7IqDL6lMpdTY3yqU7ws0D0PM2yXGlpOGUlHJznwlBLUJQ73lRc
oIPq5vd3hheH/C7vRRzGTQeV+Yh62DTjV/OEzxy+JtEU1WAG2jdm51499NME1GcnCWxtD8ShRmlu
2vpZuQR/lWDwGl86PWsEef/xHYw4OkmU8ZiguhWmHz8ycehENd9fC4uOU9Q6uJLz4rYtTvrXUIU5
Ahrg5Ht2bQgQaaIlkUUPqpvZu3KJJspyC6jBeYvTllcbO21P2Ot9cRfQJsseexqDDYMJow2oTOng
W+k8d7oTZOL9ZThi8WCmXDDYn9xybC/xUkqEgqr9jXlnX98q32lJko7aGnc+Tgjr2ia36yiSbm3u
Kh0myBbmPq+TL9WtuW/iHpEQ/nD25blR5eVNfVk9H+rcKCZa1VegxXLS8/j18Eudn010925hJdb/
yES0Dtg7Dr2uvMuhae+BidW8UHr/Dq+5BKUF2usqdMI6XudqF4OCUqmk2vP8NPVho+NYFjJVTQSE
6kQFeddZ1cn/OQfAmDYLWp3b5BTmkKZX5sSevTLi3zg/fBfp2YgJ+4g1HWaGBoS4rm4fikr+tlkC
KYYxaHPj6P5AHbs3YOcTYOVDSdcE+r9UvqcS6MLBuDhmqq43tYEh7GdDq4XF1OTkm+9rG8HvTYgy
4xqq4pvstFlMKhJsZ/Rb4NBp439P1DhUtpJ5fLqzaSIyUy01Z1tsdEar2VYijkzJr1c1FokGk5PF
hfkp+gwKhwGKYE88psM9S2gtBJl0I9yaXv6qE5Z1tO2gocKfB/bVkkZpAYhiBIAa1lxeODllouVE
Hk1Dg60SbNLWGCNHw4VOlW3kiRw1mQHYb10MVpPm3I5UXxQstp7RcUe/8m+B8sO2xDQwfFtHPACj
JJcvMfVDPbdfX5NIKBdCTNWg/ywbRQ1Jkua7jPZtPKPS80v5GvFZEudqfV1GrUTV0RYb6AiCUhzp
VRTW+bW8zSPGkfaHPWDyJ9V+Go3g+i5hGet65IxOwtwFz8kQBRlHa62R3iiYCtv0EtuT31ptl9et
ruwX+E0pAEtfJRU5+Ynh1IEWo3JdW+KtZbZAwbLhE1n+lrzL10Wg+widzv3SeGa2i4f6w+6o2+o1
Y13juP9HKGCiJ5o7gHjh2M6xl0c0Pcak3L8/4uWzvVF5pvhgX7uJLDFM2gpc740ySP8sloEzniNS
5CZkl3OzXaUfr/M/ykum6/nl2jPBvjIcmTb6iJSXroBLtLpTWX+sLgfFwaj8kJvUPuxHbsReo9C2
7RSbIZwA5ddouVa6aabB+gVylT2NzcW3Ke21n2LtBnxSSwNMFVqsirMuPCYZKex839SPbGt/JsGC
3G/qL20Clzh+SE0LUIDAoOy5XDEUa2CPA9GzcON4xzcL/DSfSHIDimDDUfKZkxZD7DtnqZAH0LJo
UROhbMftu/VRx30MUk2DEGHPoSfVpPESU4vQfx/pJyTgXhLwidHMWqk8ZPS4uvycXRd3g6YjDgJK
KLTOSTAkVHZ3yMYa6xC+xvrMKmapM4095I+Mkd0ZDg0KXbIya3CJPc2mM8+5XlWh0KLBfU8cmbpM
5LEY7H63Y1wRuU8yT1dUqWxOHqKxizeQxOY7UTMVRbvksMqvJLpOA5GF/mGwoTEx2k3VnM+SHMGe
Wmvp1hn06zdJ9YFxPiM/4pTnxcOFdwNnD1Xg+0Vo2vMw5xnuBV40pK41/49J7lHPRf6PiZXAqXOU
zhKgp2Jf2DJtvNsGYzZWZrOXeG3BpDdZD7LMHg8M9Klg4PCIHZUuYv6SqhC7w6MF53wYji257nVS
MblTDOJ0cxt2pBhw1z8py55dPl4zsGpEeWP6E1n5AQxvO01BIXQk2nL6O7H4YNnrtvjduHiVjsaF
RZ+usVMm9QjUML95EcAFQbWkJNUhxdHH4ye06BVpWmww4sx4+IOdeKkz0lvhHJg6gT7X/Pty/SPT
eAD8t+JdWe64jsOdMpAudGIsIDNgpGz7JypxcFfXOUwX75/WeNMhisrGkdv3Bn20o7fdmGMFE3HE
zpf3TlLOd/bRRMlYprNTpDxwvbx/Syu6XkECOIRBYK1JuTpx5QSh0MKikFzNpKDT/8yZKYUuerFl
x8TqWXbWaXOGSO02o2rho1JeJsypfq7u7J7MFj2F0Itxb34mQor7KyrtT5Mi7q5Tnk7RzaUBftW3
omlOsxL8TSnPDz2S+yk+zrC8vaAe9GI4dadJujDzIQc6n53twUsTcXqPzWY8AKPfVxFl+rGC/Ult
2UeSjNJFuC/X685RUTChoY9nKfx2BtTgv/nF/qC69luedIdcnUcOQ5FzOEnylCQJCbuuZr/58yhL
4k+KN4+pGYFHLxF6DQqxmtXO4bV34qrIBTkzZ1MlzfKSwyEpcorTO4AvtvdpaOxuZftXVMF1saYL
o52FBSCJZhaYZ4msom3DsRTdB1pwC2BIaRtpy2kEtDzf3Tod74BteuqmlhtjmyPF1yrGL1QuoRJJ
9E72I7XVYm6JcegPR1kU7VgEKDr1Z2rdBlXREnT/NvKvXgGIcw0rfwUMui29F7D91aczyv8C2rfF
DeUlracB90HdoJiRYHZNzcqndLg/8j59qIvSPqwtck5os1t6P++QoO8UxqARSO2fFa3tc1l5sCgg
VLLhmtVRQWYXHsJiilIFx7Z8vnjV/94Zo+ytJxnQyEDq7jzlStgsjU4wODhdAOh95KyB4v7z2/zX
7if5mOrCzAA2NytAjDhmWN1is1l4f6MbPGFzhfoVrYA2Ipk5IeA8YB67E+pIxMEWCM8xDwvaOJsm
WEu14m23xtcAeIZgDdyz+1h61pfi9e4+pA6nngfclu++sjpUf3L/uURRtRqSKJmTwazO+F9UaU2S
WWfM5X6a+4jIZCVwPrWysXM86/p3LChst5VIqdQBxDZGg4jU6TL1hjmYm0JquzBJgLuAwCTqIPvj
LkKQIHEA54539br5J+fMXPeijCiUrAFn735ym/8C7yiLNk10QGUAsCACi7nVbTxVOI9mSWfrntBG
TR7R6EFaEYjxPk8nOgPeWHJ1i5ORjjcLGGFHXGZvKIA3VffwOo568bO/vIWkR5GamTsVcKu27lhz
COd6ffmXp/L1Jc0cUwpCLVfNc/7/fHmvbxkzPLH6yARdxvhSed7Ha3lNZYsxywU9V+X6DYbw0bO9
Z5jLyKeP/1yqsMvG+DWCRccN3iCJBY48C8nu70s5dCtprkClt2v6ik2w/qi8Gs1CppLv4/HaNN4Z
NDNmpCZdjaGos7o9UKpP/2eYn4BWnO22WoMagf/N5omvRB1cuHXDU7yHJCcxLa5jV87Ql28qk75t
PQDRjY6Mwgh/LzZLCMWLszkUy63s4dwxB2OMx4vi5sl2ziKaYgoEBUfF4hPZlUaFfOlFn+3VPhs8
z/8GSA4ZyBnEXDNGyubjwzgE/czysF0apsOxbCcGKxPRoNfhpLG0sFZMAIxC+VNFh+VE8F0shC2E
rGVaF2Y6L+/GacE56pSanwB74/QuXZQjsNbjZPnvar6W6Z1YWbV0lRpF/DXoLukpLlZu/OLqFIyn
PLQ0gFDkL9X7fL6dHK/FTIBC19PjCSXOB6sYRFHoUp+EUv6rYbjrZZT3N8meyNG9TYJjztayiDNX
8jP+QwLeDRvQMcqtXhu2HY2/bjxx+EcDBeB0xJAjgAUZz42KsJxiVnUTPMO7V86n7KQm9Yk132US
hRzIhrVh+dtefGbXZe3XgJR1uIcQBeuk+x7Y6bzXZEEJ+kofN6mqrutC8HGxT4UAOUARVJg8CpNd
XXF8PzpGkef4KGo0ATFeYoh0djtjeivG0zM/OKM0kVqP5ssbBCnIhCRIinrkdaMDgOlF+IlLUws+
bA97/DcRPekjS36FCKB6OkWKNBIJOnMIs72o+/8Wqd6CFVQFIqT3NICwUwiYUhvObPJNcJFN0eBw
T3N9azxXWCPbZyeDk+/3syUzbR7xIU7Fg1kY6qgIbNqHzcyyQJA1vlk51o68UTk+rI1EipxbBOk9
jVYXP0nKHnOdfhN1emeJedJorkWA0c3uD5FDYHiDVNHUCbPNABRaoCdhy0xCGaGFx66cPnoiluCH
B1+BrGUdqNm/DS0KkrqzFbyzJlg8C7SyhAPgVJ1foRM2azJOyCqZ7JfiTNBiHK1qQaxESqYL0Vui
qjGbOd6DOEfq8pHk5R+MhxsmMmD43LEQI2LfzXcFx0zDP/A1TFGJ0FOxL8Ln3tlrWXftNQiT+Xh1
Gr35JYGX/Oj/S1z9oBF3rIZcT1RqqpoyxLeJWq5c7zCpXmDSIZvXO/cC3/6bc2l3mV+m3dLEHv5J
MsTxW2uscx8NFlDlMBAjcbAclSNS+W74T3ANWzTwHsSsnDGet0A6KPhQDvveF6sOsSUJuyxG07gA
0+MODHJK+7c9uTuQIpmTeDbw5/VmSF0AYnpmiTdjvaCYMmJ4RDoJe5IUWSwd7DONqbX749EEygx7
i4bMcVsdUWnGOUIRC7GfvZS/1UipOnEUMlTRulsf9Q1epJXN+AyOHRkFbS2A+NnZIKeW5+EzxCtX
3n4fgDXZEXChCRPU4tkJs3Vt5+eccaRM3WA8TnjyTmmm/kZeHTp9Ubmkc49s4OmMX69czoVkbMCz
mz5qmRb+F08fnQxzFHUYJS+Rrrk5lh77kzKzMZ0JDavDfOoT8ZashkelgEHZnM87XfPFAcQPe9e7
YLw+NrNgbaiy2/jqXqACk6R7IRcoGCezPrf0qOvdy1bPnIdNqGB7UDGq5SdCkHzR7OqnIM44Gd4i
hd6ijgaktlbvHcpk0lzDU5Kt/R2VSc/D4IELdDe6EYQTu4U0UCYC/rTeZvFVD6ltWUpcWk5yfdVP
ZM/zC7BFXbmmS2/cy7P+ZGEBTWiWBUlZn43r1MPp9ASNbv++HGqa9HG8hID6tOFrk+9gE7ykyabQ
0i2IoPAFEPo1mKBqPOTu0Oz0n+l49BmkqkhUC+3xMoUqqis1PuN8fg1vzxx1nVPYc/xpbQmHtIv8
M/RNIAGvHNj625crNrMnAqm8YBe1DpcEifZiK7jkjgVEMktNpeW0CVBAfvG4GXEsx+vEyC8ar3Jh
fRAMfvS3MA99Hgzdot8gtY8e2cXT+5BxOwi8tOGFZMOs3udPM6OPUzb6d5JmQZ2t6bdWgqQCjxVC
MOkGhlzLjqlbOOxchWNhEMfh21ZX+2SADlwZyulFo6bJFkPTZ8xlCjJPIBnts0ZKL8Ql166ivF2n
HEli74wkVAdxV2hm+YgczBhIjUzQnJu1H1Pr4bVg4zgD8OhO6mryogbV6juilpDvftL6Sk8QVltF
s4ushTnCgC3868Qexb3DvRgGV2kFFRhl2zcB9OVE/PFlnxA+6Ql156s+w9wttlb0rvLWBRlnf2rv
YjkvsJI+Sl6cJIOiEoYbWOxwgG6BfqWMHzCzAvUbdMxbXWlWXqV6TL4i8dRW2/RoCVFyxaucxHkU
kH0eu9rnzQwhJWmZuHmkCq6Whd9Rk/GNWr2CdAoR/UWaez70X74kWnKlO9yeNUq+m8PNksqWpp6m
32F//7RYhxDpn3wj/0YhfuYL9tofyQvHC/0+1WMw8fET7Y/u4lOtSSVPh/96pFOzXJC14aIhRaUH
fSfnzcZhAaLizawLvVLKFBKeEpc3Bgxqfm+Jij6QQNhXQmQ9O6L42j/vTR5KG7seVgfnDIYoBi3O
lZlI6B+ltO8kyTMfr1pkoIiZayncuSobHb2ticl0RqImd7u8n0wbQst5PA4qxkz4xZmE4m8Krus/
l5naid85RZUhupJWBCX+XwJYSeZCsjekWVYDM1Rcu6enGca+g3klX+gz4AsxR7y99+cEtUtRcgwe
AyE5FkzgF3Rn0qzuZbXWLJId0//1CDgKk9EXkKLQQsz+xJtGv+5dzRSzedS34JMZX3eSlVKtA0OZ
Ef63bmx+1k0IgD5IvTM5eMRr7xB90X7WdsAPl0as7MYkGZP8w5Ut5PiJNv/teot/B1U/lJeyTaol
bduPaAvsN8kEwgd9JmwDXT7FtWOvos9PEUy17lrrQEV8BT8X9Sgoes68HJ5w8zsra3Rk2Xv2Z9iL
1RZ8E6P4sKliEDtb48WCgLi4W1yXlyEqlaXCk+anrh3/UnJdAB92KJqVfR0/gEvKYoYl5qr7N0/J
w/idz2Oj3m7OL4QBxIWinRtgJ7Qlu7zOzb2w2FMFN+1dLCQAkrJvk9PDKtgqTqWD/P5fQYmccnYy
lko/w7FG0idXU2niuFe1ykaGvvOZxHO6/vyVlVrgOKf+AYj0T6BnAM7OXtuOA1CweODZzO5KBoQy
Xjg4xFoTdUxyWGxBk1Kih2SPjlOSG9Ovm8nTOePCku8DICWzyIY3789rp4+HzPWpEdI7bE6Rn5Ff
0rVPYMkt3MGpUDNYlsWjV4krhrlZZ1i7YSK1W6wyv5NYZOlbFaKRFD/ORo6ClHyo4K0q+dR7XI2K
2m9whUnCRMIrqFmKFj/lAZYU5CIxZQIiDXCSOAIq4EDJuMWGyTTE/isL7fqC2suGV6as4TAbT63h
6tB1PnvETHT+WwlN20QIpyeptFTmn8C1V8qPEM/FiJh+uDElHSLFehkHTXRq5d10Pe6OJm+TX9uT
ET8PqQyRETZOt1y8EwgApVyx6HsF9P5Gpp7mGauBUsUNcnrqa4/Gjs7dAC+bKyYlYxTwEhZmePte
MwBuuBYQqhoK7WyqmjFWsEXH9DAB85G4dpLIDItUeOLkookmzrK1NVsv0LcVJXDz/BtJ/3CyyF6v
+YmFmzUVF06VpCD8xn93SH6lW10qDhvj4CZBNhb+BkXxqjAvr3M8ETeldOVOniykHy1FMZ4xys7Y
a/p78CTGZxzL8/wgiZEjb4LBZK89WW7r07f8Brbzp17QqMuBViA3Qy9sLMy2xjfNqqdvn0Yp0CtP
UiAX7873+eBy4jwCujUKTEPrzmfYTMgmOx8hzFQHCX/YW55nF0ZGnhTrSj/lNLGBuWmRBl/WDHmd
Y9JZvEdcZOFKiAabddp1vUPcIwyBrrgYjObu+t/mUmQA399IvQa842AwNsm3Ohm1m33lTXO1ksoG
cqvHqvStpMKLB+95MLhz5rdsntTDJ56X18xKWFjPCNcEaUN66MS21A3bpryzYcbyapcXDadWOEP1
N6BXZhEE5koepm0oYIlWbX2hGymr8jgl8ugmYIlnzvmEBW0NB96zK4hXv0aGcUOUgbfSrltaXWmZ
P8zL2xNjfajg3Qta9GAefYgTrqtMTAAR0SYB5JfA4JkLZ861YUHYsweqeoUeUYMcVQHKKgtC5e5S
QDPgrzW5nJASfC+3fyC6vuvTbX5rMhQDp148FhBmo9FT1Oh5JI/MIhAygpzF76MrOLKjACNXWWyN
1xM0lizHLA+DdUjf3J1nWHbbch5NSUylyWAtMfePSkmLB8cl1iKcrNRcm1S/YFKsi5pRBeIeXFls
VHaFIXz0iHbhnnsE0wttFCKEhrR3zzoLRvOsopLR6SKjsvPCFQywv09o2yp8wO9KtR82ogf4dYda
4cNx42+GhraPfpV3AbrHr8cC7qx8h7rpgFKQ9W43UIWG69kIoiO7lbWyOz7frbdDVcbcJzp1hhDI
b7J7c7Ix70bJlZuD20E+oTaqtEYSfFrBVju4hoa0GeZtx3u23jhXR5BOlH0ik0RhyMWCVMr4DGmZ
9ydqoh3DplkYKMWwpIQQtzSZrC7IJhx9B/Auu2YV/t6gVTmYu8t778KJb+EezechfAvgGsCFsHWf
ORbacbhBgxuPEDMiK4RAQ4Es1flsqx9F+HR1uY2xpyD94IOGURjVQ/qGIHaSfwrkaunexgooeI99
bZWX4Fo8LHcSQU+jZYGYhDN4oNkoOco57JRvs04fxd9yP/ZeeZcBlHBVmzvXzhFcYbS3KULS6p7Q
p4CQwtAgAHWAxgoecRsHNHxCaXCxh+h4/lCKyELKLptuJnGFWmPp2RR6CT4PA98BFwGiLqvLgvfS
FEuMTllvm0EYylurX8y/vka5Q52HPoEaVPwqHMCBbPFMfjTgWmxZ2ME5sTTm35zRWSLE6Qs55x/Z
7XjF4mpJwELapNTIufYOTYQw6cTTyfRDVrKW+R4gpl3ssUQG9OVrLC71XHGKERQ2cW0oIYKuwoBg
9XJI1cp6TnPq0xcMSYHMOtr/COx+mO2NmZX1x8KjGqVxYskTeoGDPrW/HPhpIim4Hc2K833UoOHF
g0OuFoPV6IjvTJtUoaC7VJpDXsgJ1TEcgqqzMtCtz+8+RFdrxJbVTVKq37VsRTUjd59eBlq0xT+h
Qqjj8kUImKUEMpM5kBEVqYq7BKJbX/Hqj7uE/ofw+xMwBPBBH0TYH+tOpxd5L5n+eNs8VuLwM6yg
nZrBiQ+WW9VYkh4Y2dcHu1cArSwjkqOerXOKRMgzoKrZc/XVNvzb6f70ANrmTlDiqOCjGHo585Kw
rSaPbXy526I+gRDNGJTIRcEdUc84Vyv0l2HCPCEQ37MRd0BQWpsUAuB8c5d3HrXUxwoY6j/sgHnN
J1Ac7u/WGDFrbiyYfUbA/fu0r6lijnC3AsS4xKW9/rYqR0hT3hTpwZ7VfnupuQRjkgrhCkfX7wUr
9j8mteVerSMiXALI3b8X+KgttWTNcBIanZlAeqX5FecMdEnGkF267MTsLvhk9NKMVU+FnYVSLuAI
kJ4nzkK6xBwX12hmWGK4ZNjDKxZqqkoD6KHvZoXms7N2008vprSonX7VyKwsoW2xerDzjLgOj9FK
nNidfQn5PSdeqaNarkspQRNDfXX9Sm3Xo+m5SMHqBukO72lKfbNzbd6H+INxXVxXaj5zJLDJyVv7
5C86Q2T2hjpOKbo/FkAEVx0pCYLmoIprIAl5T4Af+EuVPSlSZB3jUZI/+eqvY2h4qYcaHPL5uxhs
wuqBLjGgAJ7Fl8KEFG4JWL57IRBiWBDCpvhSuW5yFf9sx5NnimW5RbtDpfCAcMrWRAHyjJUQtX2e
hpbxOpoQc+bUTGK96jCDAcGR7tuWuNzOl6J2zd8BcTQHt+MmHM6kIB14F99HSoHxGrow7eoHMUO0
NMyVDWgQ9pZFhR3/NxtBQE2WKTsdjJTB4b+7rNODO9KSRwV33Ow84K4ceak+TO554sN0aTVh42gu
kHchARj3PORFyvKk20h/XBIiwCJkcdda6Cs6ECR+S++KxQVvz1nAXSBdWnw/rBoALqxCMaP1jFhT
5Zf6GIO4FcHB5cjsjKNRF+uaRdgBCUuEnQxZOqRFSQW74a+yItQeusTwkSKb3fbgxwOeTiz8MSG6
MTQgs4Oj2vPG7Y+I21l1r0bccw+3e/XVrCgQr+PyXOS8w+nLF0NYIoSX+fZE0wNF4rermb5ZsrI5
d680Y0giMzmlHjITiweWXOCPRSuECZ/dbq8gpCqGo6B0HX1zmsKWkhaa4ik0k7nYzOBYDMPhhDee
fnSQC4Dv3LJAcqdddfUtihr/frcTnBQbv/+5otH2V3w/Hjjx0TRPkBjiyOZ7/nmKR4dZQ8KiMAeF
Knh4fbU+WID54O7d8ecUeJBnEtRK3xLVlWWMYCWUoWu3B1za8Rqc+12jCuZHC/yIeokpjiP4zE6a
rlFyLCUSi1nSjbwl0UCqAibqPbi4wqfoDK8YU2ogLdMJe1JMQYJ/KPFe8b3Y4YVc2B33NCvt/zdv
XB8EYxKQ7Ptvvx/5xA2opIhRsoAC1Z8MLervkNlBg7f9rVRn/Urtd1dr4rjL3wC5VD/A6kVvqB69
xRj4FkelOjR+NvPCatZj+tFf6qKQQrYCz/2+zLzV14qMuQTuk0xYKO+GuSSn4tNOjt7idYxUCl/l
AWhvyA4rbJo9MeiJsLo2jykw9uNUucAftb0nIQYv/vEq5B1GjSABUwMdy7wKcBBiJSIgV4f8qFiQ
3XVsSTvU73K0i+qdlycPJpN8K+wV22rDWf0RrG3WWmLaCJk16GyKrdA2cOCHhl55tE3mQq1fHDE1
pTYl090/lCLjFrKHwAFEbyhV7AGe69vLc/96urVFM88fOqK4urRMWU0OqChdmZ750wogyNaBcSVM
5aVxSrQuPve44AbsMzh0KB45Uyzia0BTL0vKXesW21EFT8a0yKI4p7rzap/vdpyOsnPp0adyyDSc
e4CQ1gubpT5uFyONy9w4P3IROHwflk34nbUGYzwuRxyGBoUWaQvS2qQA0EwoGqMOPJrkQYl1RNsc
ZL2hPNTUugjdpfUNFR2wL9wQXxhYGgE4LmsmPaWD1eAYBPYSx5MUrfL9ge7JnttsxFMgy8Jp7QGb
7WrCB3zd7pglm+00cnoWG3rHWOZ6Qsal/TrLw7zRuCho4coSDG48mu8BSxeAnJH4kfYS8+xvYCw3
DesViazVss1CkhdzqYU2c3CbH9Yxv0M9uI/qi9LHCnkBsQHo7eMjGZD6Ev+4LvRosaHgQd6uF4JL
bfYHJU5uSclvKykjtJ/B2mUjBdymfxQSO5zyJnZnK++oJt7cDCbSKG04YO0PZu41roF6j6O0Uug4
x7RYDKtpgm69WGCCxoDJjnQVFhnMJnyoQKYfNuESf96r4MQHMK5xWe20O3lo52hanGOi+03Bpuws
aiimeIkx+eiM1I+CkquA0y+xO2gLLfjSmbSav7MFVmw93E6jrqLCWdf2BcjvqzGoHdo2tl6Y4aKA
XRP2tVg87f2prFofh+YhcAClTyl01RF44SCtWDp/jQgg8xCHIULsUWshMdw7vEnp/5N0C0YwnOOR
rx8iZfU0rlsXOCFCMVlYoetG9aYXEPy1i48YT9/6TUsEpguuB5SagLma/Wq10brWhM+bb4HkegNk
3BeSKW2UZRQgDDU+yY2ncJohb3Nzq/MhYfNjLRgF86/0Cd+gDBhBu6IXpkVHNjEopNfUb+7A7cqO
Z+kNM8shq8kHJ0f15J8Mof1O4Y/rNiPM+lZ+yvjChootSU/Skgz6T02gablyU+ZtvNOIO/34M1TY
71vQKVJ4wc+toQlKgsd4qvAMweSj9wj5SO8bqSMCzaQGMyMo963wgDSjAk/ZvMnhS5VVkZjfFy1l
CHO6BBW6MY7zR91cwVdUWp2tgfGaEAdt5i5Q4Fm2TpAUYSA79jBrY5GE3Y0YZvIASTFZM6YdEdSN
BCmk2P7dT9AaxOR4erxxQVBPFVlqw6jDwlnPm+H/4b+hR870vV+EF/AjjMYrEx4pouJF3b1mqBYT
8FVwA6TqL2ar7WfamUPbKNjGEagqgys1vG9IkavuTVDj8bR/j3n6Vj+nqm40OmIcoCa2pA/oqNZa
jdZobMPY/akcHJw0h2FkN1RN1h6YJo66LT/r3WSEiDIfHa7GjJJcKmCpSqSZo2P1mo8kHd0969Kk
eBdsAJrGEqaX1aWQweBNs1cG9sZ1CFCf6wYNcHAR7v9W4sZyRfXnSFC9GA7JwRnjiH9Vh491ImqE
iBsuk/zoHIkId/yXqx0v1FcS6xsCrLtcysEGpqOJZlIPwqXLtCgbALxa7WU7sFbgHjAIYhb4xU1p
pZUxfHfQCAFy1cJOurOZc2+dC5aM2a7YG4CtncBT0goyXWaMR4K7nQ1MXe+9A3cwmzg9bm5krleB
EQC0+3bFfOD19C85lavaWsFHAlzO7ktmKaAh37VlOkWPKhhjNdAowmeycBML22mUFZrFzUAOQs1E
X41erKQ58hZ70LZ7t6e5aHH6uI4StfQ1A8xKubCXlCh82NWEfHnxMBZs4lBKmd3AeOo1v51hrB8Z
80lfpKw8WjFZELJcmRHTmuObPDjr6/DnBMsUiAYhVDM3pf8cWM3qUv4dJeBgeoQWcFRS2tl214ZD
NGXrn9aBFVsPi153Qy+677q+dmhsu0YWlUpM+CE2AYfayM2y78y2yfea30Lk6d0YtbmtZhNPZumj
36GMcAND7klZbqrWTph/Zx6ZTvI2tVlUsk0wKp+BU/YpMbfD+NsTvZ864e+wiKPFjOt3sHpRuwLF
0+SUqrg/5/B33eKAYOJJB4SwRt1H8KUOi8Vbc5Nxlf+qVNoItngfn7k8pClnoDuQT9sqgefK2/OE
x1jWOVfJM5ARnYkPEsCXoC76i2OjdZjAXbkASZEvUrbq2IoTgKGUea9zz5+vNraddPU9qg2LvmGw
It1KH2ndk82dkycwowTQ+bmND9aTS1xVOrzLsNWWnACc0hvpHeVzeN9hiczqD3/buO6Ob6MujphM
gIzw8AqAy8WYMSC287X3aLhSWUBWQ6BU0axwtAwqy9znlOud1wvGfeANNlSeQCrRljO60NoEOCCE
Mr6L+0EBBB3mX4fxTcl7riOXNaAwgkXjJIaAbBDVMNzKIwAG1Bonp158syFLS40Ih7EsAUvdfQ1F
zq6afgw1IfUs6J1e492kC7EZyR+1nuZrYUN/p9nT2EVkIjjLgWm0vYYpr1APRXVmF5Ph82+xZbCl
GxVjMk4WQVhaEC1lFsuuRhzPqEH15IInsWnvBQTSlK/XMzru92nHLzX668bUYqg9MIXcJdllibWS
pbWrzDkaiXHvwKYrAcYkuTpB/E3uTuVcBMEGZesQPemg1Dim304OY+BqsbqiY9mxDVMLJC5tbDUW
6NrDMN2hFE4DgC9I472eXnOkkLXkOklSQ7IF6oRVyCFZX5zr1L1ZOpVo8GEBykxVMYbb69cnB9BR
v2znhdWqFxCkgzQyYlcax1ClO/6PxjCTeu9dP3oSinArEK22AoZ6HzmsOQFtFNLKqaFe1xIfxoqT
nvFpaf0Pabh8cAJhGZrr02YayCtQLlsYnhPHlkJMNASU348MFF3DWNHNdLVYbqFFpVnVDXPJr5Ji
fIgk3X5wzSPIjrmMWjZ8K3C2hZqkdZrSMLJKKOUE/+6rHkRj6ZYrEMcxYUtnNNqiK1vc1ED/500V
ZNuSR8J3uGvUPGXhFU0tvwNTnOHS8/C7ceDjyP3btY/nCV2fEPKVMbnpdtSjFwLLIBlkx0PHsK13
YcTYR/4wvWwOIl3YOztQ9+zbnz51deB0SAx63VhiJJ0KorTfVBqrZuw3tcEyMDPf19mBWuWhluzE
FX+HEzun2eiqreftFN9OE0yRWcLB3pP021Y1nP6LNu2aQSaT0wVUdEeaEnWwtGr4xjVupfnGIK4a
MdbOdkIcLUisAp0paAUePRlFf6VRimwsg0HBtPJfCtbsnzAciBPYpPrAvWPobCGwKC7c1l6nK4iJ
zQ/xTTrvQNKBMW00A+DbPYGhPryostWbH1Yrq0QAIOXdOo2kj2YEEj0uLz+CZjaJFtLvdCaceZ5T
x6q+IJROJy4yGMlLSWhnv/J7UmRZ/iy/tDuOuRoRwx8akByCRR+9tU2vUzJ8Hi9/XYcE6MBxCtks
kkj/okSEovKBepjFBYt9eapdfQK72r1Q0eHlxRi1A7DbLM3lmSacMMbfjmDq2LuJKz6SjqrtdhZf
sNam9qPD6h5F6gd9kXOzx5Pd//ddHs1o/RKZG2TGdqdjo23oGCjDfv+8/bh9xNlaRHPbhMhxhixR
b+QHxgwJVHD1o75dd38IsUKqsIF8h976+6qh7In2xnjyOw8y0hzwfFZtvUGvgPg/ZP6S9lEMAhsB
cH4dmb5nOmeeaoeOvWCJAm/qHhdoFPSXFnXp1Bquc/9hjP6kqsmj5JRw7ik53d1LkG+5LyjkrFn4
P3Kh+zr2kcP6e3+g7qYYRI6ehBQnfWVStR7TIMMv5DltcSWqzWyytgYHXz2cTnfl2HesSwVKuA0Z
ywSwQ2T/aUV+KqecDEF54gCjXJ13QF1Clxu6M7SCD6Tkuksp3xTINIXfx0Ja13iafPM+PRBNCY8r
Gb+Vu56g6Nj15dJHenDA2sfFLidSkWIy0AqOpHz2HPUWXCoa0VV7YZc/l1iqGFs+Hb30djabke6q
JWr/6lT7X+tMAGSu3rGUKwNwrrPCduqgcs0BM97aZqoiau7vXJNXYgsAr0tX4b+dzmhpML7tnojo
Op/Zzckd0zvCnm/nLKIMdc8Pe61zAGbY3dbdH2gAxMvf9DkqBAmJ9SOW9CjqZeoCJxKfDsVaW08b
pr8UD8HupQ8EXYer5KUmPXU9gnWv52qDfDDhzciQgdUEoLt1NEv4itppb8xESR19GsXTJH3y96LQ
XyAMnxxdzDCYn2jgJQeUV7y+eedqJX8jkKUU15+IqJtDgbOf564Irw1joXXRVhOANuSWvse4XDuV
pifgILwKSUCg55ApTGQM0Ma36K8g7Lx2PyUcQwntqS0bj8KEzlZVBrGaje6p1lE8x9/Hz35tpKKB
8Fffdxn/ldcF6gqI/YLNw2QH3e7wmTkon++uLcVDahz6fW4gSYUMUZ6fzYvWCtAxCslbtdmaO7S+
2jvmNOzWAxbh9bckOmpg6czXg8VnuDthGWIFuptaXas5GIEqmCJ2l2nih3poWwi4y7BDytYt4bv8
aO0tblgxUeq69DBwEhNQJuAtJre2pNBgV0T22SYQDsLpwX0YXvk4pqcPuxkw0HIVpe6q3sCVtK+Y
Gi4hX2fc5sHfW8A9H9pC6Hl7i0jCMrOaz5LmCPk7aGzWGyrUqqq1urXEqasyxacYRBmfUlCvioJm
41pip/SIq3Avvh1eBw6CK2UmhBTAtMY2/Jy8HGBDS1Lw8siX6efMrfl1yO8Dm3couMjR0+eRYTzY
DgnfNb+QrnQ7idAHcAl8ejPaaNL1R81MY9BM094RlJDKKGjoIUoRJq3f9aBZoSRDvJ/iGjPz+ErN
Txo8SIi4eipH3JNniqTDgRs54EtZmxjGZeb5b9zaEoCUIo+BSQf2WiI7NXAxU+4ui3IIonPCUAfF
gBfIpLg4QfMwu8SNmoJApU8tmXpgmbddfeHl0zysjMuzscKggDQGBC6kwsvizzGPzIZEsS7/wrPL
Mejtzd7L+dE2nD86ONaN5CqJTFdyTAARZzs/rT6zX99+bs982TBhl6jZ5T1h99Lyy4uGWYmTJkM4
pVl3d41ULJ27D/Lv7eESkYntt7f5+mfp4uh4Fe0qJrsZbjDExs1DS/QRDfmXR8GNK7hYhJo8ZnIB
Q+9uhhmjbKieayL3YkqTsnAeGNpE5BrQrLCOa52oVvTE/ZAQgRHnhvHYOw85L04BCB2aii0wbf53
KZoSkj/doprDoMKt9Ykz+/1Xes50P9Gkfd+KVzRGdcFd2EtblCCLLWNwhLn/4qYCqeahuRDF0HmE
VYGjiEifsSKMeOXIQBTDFnEBb4wCq7L1pfFpiuJTHZ3bvz8JQU44ddN6nmUWKWamgoBIeYi5/24d
WL8u/qBvP019hHBw0q0ttU4FFgMFj+Aq7M4e7Ct0HzVvkaZWzn0xMppbYLPDRUyvVP1shxuEwiYp
MOI6zMYKzGCqHUuWvCLXthwfY+RjTp/LPJKiOglLGH9l2mpZUKoz5g5d+TbzGmX1KI0L5FkG2ntT
C6Y21Us/TAeWRB279Q0ZfVOaVeRooLT23nT3oTx4F85AhJiXy0dXvSn+pjFJamJdEe6xT2XYhTWa
FckLFy5+3tq3RIIALEmKeYSfjikd+NqGOXKVFsMDDd9fjlXtHsD5UPAwtNqUSmViMaVvuaEETdN4
ZyJpKZvVmqm8YYbxktmUjJqu0PJePvinoeiJiGwxOAXcdRdZVcJ6FL8mRGppxPj1rku3Q1boyIJ2
x45Z4rg2g3GFNq0khcbnzKxZThrzUNfNUUZXpeTqdSEFLBYMkhEJlP1SwqbtV7PzV2vZ27XXfqum
pTSVl69wRUbiWus2QjX6izCRaCHL1UWFYXqBtvWwcoJ9QagStrFdnR0pb6262LiyrIK0j37zltde
UZYVwUgjEODeK5PByD2GqVdFNrvYAhe4gPr+ANWP5Ec8OUJB4y2CUD2JrFAuuu7JPXF1AY4pdqu2
o8a7i9n4dyu/ZQvE4KMp0b+9h+a30EAbaCqQIF9Jl1z4bgPTVQCptQmEWPzMz+hVepECcPk4tNd9
jA5RwTBc6IP8VmMF4M61hPFClw3oV1m6H5Qec3mwiYSVq7ocuqS0/3u1IpKN820AyvelMRGicH92
vB9xywqUl5HZDRVm8S9o1roFstHVEkRWeQ+MEZ4+gQGjOsWoGNldW4WawBbe/Vej+p9x6QyLDPkJ
bD0QxKNQ0crZSfDaccJvUlnkobN1uhDRr87fr0TkM+NoWhfrLWF0mJ/tDxVW9a5tmFqZiK8+6G1t
b3bQlvOP210Bc2yoHh1tnIHzjMjOxn+6/mmUubkQ3lgSEnEdYso4MFc5R+eCTXVwgehTYE+yadiF
yhxnagKb3Q3rcT1H6OEu7CQc7AEqG2IWYMUTKr/70AWLWKE/gZKDC/8f3o4oStMvsxYxukac2Fi0
70WTBy5GdcMsJnkFVaORdDevEYIfsO4o0UdRbyiMIwmOE6ncLn2PviOdzhAS0jryomjPdM4XiQrv
mdZ16Aii7Tx6DryFXGWEoKb+cSTvzRFSGfv9quHgQUyH25hdTYFmXQPY+ECDOVMFXrOYJ4Oh3CQD
amSSeaoKgCggIHOzzjY0qKfgxWVYtL78xi1SVC/5qBEizDTr1pP2hFKdf8bT8zbNlVknvW9U3e70
T1fXB1kdrWrE9dCyT7YTu3PfZWPKU/E23bydWU6uqaw7AFZftiJ2HjwbRf3pcWxgd4RG6eO91+bq
9T4LUZF/L4JcChm/LrAfojnmS6OrDRy2XQGBpJgXGgIHOYNr9j4/EAvAAcqANpiI+ABXUUmWTcfy
r8EsIH/Lx9KMwjYYZ9Pyyl9Q55EqouudUPrAryYUUs2KSCcdpUFqSzFXnob+EjUvEnu6z4F7ZPl1
grAL08by97yjP+KXEGv1zwMFCXDVUTtBb8AyDn7KoeyUbnkmmSah+mEj6IwEvRkQp4IRsFHtTVbw
oq+Ognia405KESSkT+pQo7FFTd8YIyefswP8iz34KP4Z4IozCKf3RnhEMQdJIcF0v2qXex6ImejO
97/R+8F8XEPm0M9HWE+D4kWS0lxwHf/KPxh0Qlaj7H/0NooIkXCuE6DYVTCJjZJRwXcXEbFXcw5V
VDAIB34qJU04dgnJh0lAUZZg1A54uPTUII7V2LmhoQkY0hATvozPav4K4rAzP4D8en+tMmG0bv+X
H5/P3FFbYhEbPtLNXnENOpvcb8eR/dmbEkanLzXKdJmcz9kcxV5UY/dP83k2RCuIEVMMNvUDLHT5
gcTMZ8c7Y2O5DoUofppgwLHZ7ZpBoojeSSG/GwoedByKDjKwisaZpk8AB1Qx5fke3Ymmo9/OmnoX
zY31EfTPeTA7/kCDNC7CI6VHf9HX1bVA08JAaBjYvDYXG0OJlX7gjN4igU4Djd7l5HBsSJCUDpWJ
vU2xFGLIcUpsdgdSEVvcmYQB2y2eyP9jYvLOyroaWKFSgyA+5b7N9+84Kq21IR5IGJ8ZU6DDTgO+
H6RGoRfU0y/wsmvOLSX2HeA6mUEZs1XCxDJCdjuFQHen56QdTXVpqWK5P70BrOh5OltvUNpSNRLk
FHCAm1Le9n8oILGrpB6MYIzBzZ8EzTcUybYEOEWPg1hfMquE9/1Y4pz/+BJYiJwlglte1In/AXDt
77p6dzOf/rwXT5wVJdKBQUXpWkga8qBJBNTC+KrvWHKD8iJvTzi7TRkoJLz0iOuHWorCZp8f8HJl
id5rjdEDtx0kc6Q6L/vFeiWtFYZX/WUxQYbGebSJRms9b/pPzU0Klb3BfNLz3nLXvt6wLCsIRm9r
VE/B9aSS5Wl0+0NPaA4Kv0M1cg7la3CIy498WGrEyGE8N2h3z9TKd6zJ8R9dqKDlh8U7Jufz4Y3l
tOp49qEQFr6vuEIK4orEDuEnt0jjgKP/6N1HicP64UMM4OfdS35eHMjL4+ZkwWzOeZH6Bku7RPv5
GLq/iCDH5OlUVeP20c0K3zYOaxQ0WqLXGGFosO7ZiSLYdr87JcAH9tK3oVmo4rTQ6Wwl9az/UJ+0
2TbOMUbWnbYzMODHA4GF8+/9RB2CC95GtvusajRFYHJx1BxqOreilATeoTD0I2GR85uSsxaQDkjL
faZ5tJx43NgNIlZqva+LrV/l+rJhVqF5UuxePRguBFzIDaV16cn+l525bbgDzIw0J7rvgiKc22ya
onbjFnFjQ0A4PrYvLnlmkwpN3NgUAnnO/u+FOTW1jb0ZrPqFX9fT+Jp1nCGFMh6J2YaCBEwVTGhj
VaxiQCrx3qUbsCUJ/QfoYH8pbNGAA6Pa59PIVMw0ndMJhNdfVnza5uTd/S5H7dMkmEh+kwLbNt5N
OLYnOvUO/T9O9UhQ89YntKLhl+fVi3uhQCDF/8zwDKce2rrdtgy6g/RZPSGg2cj7F3lPfmjJpi1v
MpQrTLvMJdWG3IPm0T+3vLMocRG6mfodXlWb9WtvqSAD9QxcnNiMna53VwA9hSfVR8iDvkHpN6u0
UNYT7nL3zvZDnULIJMrPrOr6WfC23xXIipUNRafpCaj44M9ykPKcI90VgRBse4r1vHFlzZVjFFOp
83vSoBf7hIB3VOX4/pbtZEiiUD6Ips2S3mbqgupjnkmAq5qGINANgbhqo+gPEnMkeEqqxWkTlX2S
aPXkunydlO2lGAZ0Tfeun0Zl+kF9nU30YIxwlqx+dOAJnAZQC+FtZK4nQXMJP5dvmy4Flo8GapoM
EosZODNTA/FpAkU5dR+DhjJmX7H7LNsuLEmRwsxyKnVGCQcB9z2qoLZZ0nmRKPxWaqN2/vULMHMw
ochGi4fQPNEg2BVi2sOn2PJlnwZtIyQKVsww79qYzB6a83wlZ9E5uCr3znfq8yYCtF46SkWXQImO
dfRsEk9LVDtIwRTCvahUSocgE2QzHHBFhthYDfu1Gs82mgy1NYcR6T/WFBcGAWJmU8iKB2V8T0Ds
5y6ggsEh8yms/JFtwiw1GCFJKewrEOWTU+iARMTcijtOrZ14Vi+v1uE0z7TcNxdMidV2/IIEqCRL
gtdCLfal4NThDc1eteSQfGLluxVaETAmIprzVP5rIAYNr2JST07Xh4Nu6WrtMuY6uC0G8vNWUzR8
GBTPemivAAubqbzE/gDcRvcLuDnuPXmYDgqNcEvASVdinBUq9IOV7Se4ic7GxwMZo73NM7ToWoZ1
WOtVHbE0TA3g81Kfs55ckqp7q44keSiRrYjQzLuATHf7YeN1viCgtopJq58HcWoaDZFKLH/iYJ9/
utOn4J3gRPgTf3bC6EnfZuOPShfLfVtk963vXw5lpreFs1b6gz26fcLOpcYMgp6aTZ+Zq0nZZDKu
Ny2ThUH7EdSh/Jgxe27+flaUUdQ2zHZYfiqvCgqBeUn4ZqP58sZkJ7dsaAmzqGOsN0N05EMYgHN6
DbuUuTPd2YkM95GentNp/P6TYtaZ6f3NSENJAvxGvObesPnKmj9fpaS39PQ1XAxn85cnT0nHwaln
ASE2xMYJK+4A3vffD2wAIgt3l7RLM97cfQKd2Vr0y20KFB1ovo9WYh4WgUxVHAgnMVUz6Cs/UUpY
NAGTBQE7DgV7LWWDQeoB0Ste73p22idHB5c7IHbArYMFXUqn/TxkmdrNhQmatTwC8XwWvgyXXCcK
qrPewdILZJf0Lv+9Ta+dRYPuxcYDMFQckY0KGbjoBZtiLRA31JhvQLuo5rgMCrP7y/qUt0qcB3o9
R2HxnlThj+WTVT3fbj1RmK28qEtyOv4h3bzgSbPN74gmGqz42QbZaRN0OkLYY7xVHVmnEbyO0cyp
e/RVP/RHuznCjwPNEg1/l9Cco8aU1pnE/kcLmn2gRYv/3on/dbwxvYghbzz2Vmtj3DQv7AW148ru
lvAwBlxNwcgJrzW8LzxFhidmtqwa84bVbLgVMpRN/KoZekIBfmV6KZxNQiUz6cfhdUde449rxaGb
6PSUrdEha4WXIq4mJQxPFmS4llSS+JncMUPDkZRBxq94qZJXbaLQbxVY68hDZ6qtut31wkLRgJzB
RoJ20Olle9lW9YOyEpBkOJqGP3kQn2CFOCgFYWqTKe++keS9xRwR3g50voTbGbRXbMMAQ1iNxrtC
EOVopMQ3GSbD7j8g7WnVRg1qp/LiXiBkWOdRHit8QJCBD9rd6IjX76HJdjrvH/KHEphUM7B39e4l
WV4viNm1+Zv+9JX0BuH3pYjHAUril4nQf68nhX4+nqO5/IDGixa0Eg62n+YQycotXkWNk7q8MlJc
+tp4yg8OgLCnuPAUJAOIrs/8S6ZLX9ddJhCn06kihi+eCxCf0vq/EBivC8amzAebdf2O5uvqUFwW
7nK4DPnRkdLXSXuvpTcmnBsSed10ZOFfI3k5KlgBUsHdBoFoN1htg1CHme8TpBG+Y39W3yQHK31z
g45FzzgS+yQnBPO74lj8nyfMedjrQx9eoO70B9RCVLhq8VppYzSUXBFwJ1VP3P7olgVdHY0cL5yu
UIUqSWtRfMzTL01BlLQhWH9sGF3JEmBzvMPWtisMsgEAXL60FR8rO/47COuuiWXVA3/LIK59FTGM
F96CKjRpDSO9E32ze7SRs8VJjiS03OEWIhtfDQJC/WZrzdgXIAZUlJm5NYWBwJTXhFjlH65X1PHB
9DczkBdVqAvKB34BFecOEpGuVeNjurPbXzg6wHV9GLiqyjQjwQde44L7G1YbVEsxs2RChgDoebl+
URVn1VQqAdOOp+cEZGFYVJJOZp95fyLTP7KiMdxqhA1QP8/hcmOYtZ7zFIJ0mmbsh4D09p/tojzg
J0SdcJFMxJDa7p5TS7nH+Io0UrsqRckDRyWh1eoi+n2orfruG9inJlywMWj5qSqxObtAinQy6y40
uptoIHt5ZqrkEM5J+ZguI8026VmEVHgTdwII3MW65HNT52VuY6fCX3TrKUBz6qYFEz7oIIfgB/Rv
pAJSa+bysXaRJaiRlg57Lo26kFl5NzDpabIXVBmZllZBHe18wRCJf/mFFxPCuE5pjV3JC8Bdza9L
ekUNdhcV/DN9XHbC7sl8Q2Z4buUQjajuJJ5b78oxFfNid6fESKxFZCtZp3ntFZSD9rlHu2HpgOI5
kmb7z6uvZoXnciAfAAIrOYMTr6CJRqD26Hx1hY0VxF3IydSZVXwAMVywUYjqBkwl0cREXws0ydJI
B52kxJ5C+XhsBg/Leq9rlje9iIDXF7wbbcAeOIq3fVG/00JBI2bt4Rhatsqwq3sjW7H55rpJDXac
FF5b5uf7WjYlUbAcVqBnWwfkDeK8IK38zvLrONMvGmBz7daxLJm9KwNSSyQTW4/irfZ0aU/bPE8h
wwfo0jYg+8ZEGoW9e2HwAMhomFXCKcQ069a5xmQAtMijdsGYgtvra8y04ebB5hgq/xEHinw1iV3c
KJFmpwpO4XwAoPn3hf1ZkV1ovTsT2TawvebyiykiIkVQzXOyc5PzERybfxg7bK1P+yP5HoANjTvt
U6th9Wpv8D6DLMDt3T7R99sEQ8sberfemqAJ3WMtCteFH05OAByrDmj6f/sQEl5DbLkOF6WC9NOv
3cCw31p7YmZ5kRJtxT/TO9+WmIn/WbvGVwiPgxL9rrDZSsqfDp50ZIQMjO5DOcXAtr91QWqyVM8N
g1wVZAjrf9uVgX4ub6JGv2XE1zaxPQM2RebtZkJcPlTFYHBOgVL+gBlaBLNexHXiTgzbUr34RQjv
7Yo8rhH8dF9sJcuQRw604otun4akups1QF8IXS/F7S6xuZVont7/pW4VOC1HyDOFKy2Bc9oxS43G
CtJJzY3w3HrCpMDIZXUbHoH4DSLT/US1kq00WYG/TZEzVZ/xQNp/Y9/ab50izkyJ1t1BWQlGdpEy
ThCuiETo4mKIWHl66kQnEk5/GvpfdYLXxvPboB799XnqbMP6V+Sdrx0QuxwKR3KYqQYk/eqoirh7
DbbqZqHilz/dSZED+VrJ8T17T2niqrKUttzA23ujsXX0UntRTC1WbPH1ED9V9KC3Ogqc9KzPH+b6
FAEPI1TOr2t/n4zso6JSmrLDLV25NtzIogvjrenPfJ3TdvPP7uG6tP8bNOjdRe1RVA6ouJnJWkbb
2PZxosv8kJJnWcKkypxghHzgfvumRtvIQuAf/s7F3mNy+0oB+GM54/8rqPragJ8tgPH/1XlY4d3+
9WIA7aMn9Z+R3b7Gt/FdxSlHivdO+SyIXWhn6RsOSxKVtgmWGoOd9sT59VdrsRP448L3uOoEkO7W
0veWq7GzQT1c9eFBRia5tcLGk7/YXrGAPmb24uz9WWeXCRvGLDepp+6H/Ns8aL51bDnsnkcy56gz
ADCyizqA6maxdOxGa40Y4a5iU3q2MEfqoXuTUlccCP/k1xBzNCddlBzCavSRpGJXLU3mTdOqKb5e
+UIOwsrpJtdpdFCcPMQY/DEbTlk6iJKCYVmTolgWn4reMiAjgsC3gw7ya7hluDNyY4TY49cZ/av3
e9mpJb28q0RmaVhlr4Gw48+xDyJyS1f0GTMxqRwf79tebPlvEFIh04Ibfd76zlBB8vYdm6NPi86d
oFyhrZczaFzo+QwiyHyYo1tuqc2gwT1YJnq00pTa/5RIMw2IEIB6MA52ZgLq2WC6TDDkPAp8uZpJ
uY4A5Hp2fe8Tew72m4oXQqWay7AZUqGy/GEYDdCvE4sc/i6B5/D/Slv4kmDw9FVPPGk4mfBNitF5
+zlLJZmBqz6eC3vlwSwXsAJyV15pKOnc/hY7l8T48kpD6PZI6EqBl/vqKz49TF1HFVBIdAtXPUO+
wy+Z/VUnUywYBr92mvlxykGVWJ9CurpwTsBvfBhH+ntu3VXc9ayt17EpFMOZPG+pU5/DhqA6pQON
2CUUxcuX/LpOgrRUcLmxHrjg5ePQI6dqXoienKpNJpX+0tMKAX4V19jLTNDYGvgVcvUAFNyEcgjK
rxTYbdLK3ThfIF4h0Jq6OnUEapQPwJUvlVMH3zSqfk83d08hRRww6ZPguDrfOEmdHu0cEEXOAX0I
b9ve7PtO3D9EC5WvOTiCLqoMW0sOvBVGZIJCOJRd8zC3M0B27fnuJAHin1/RKfQiTEW89wnSV9h/
zuowEW9XijfkMX0WJkxq4eD+k3gjtE5JWEdiQWa8Lnyqg9yerwRy+7ll7QiPfhviAKwgynacPaov
F3yW0fLUH+ribzkPL2rE3g/gDjcNdjKJmxnsSo9dM4b5upT7HjUcx5iIsr/CMriBCr/F2JQdvwQi
KBn7kRL144hmehSShWU/+8N2dieCE9xkZxzcn6Fu7k4UDpZoL/V+Xkc+UJIXIzyDJfFGxc3e800W
9b88fbO2CC+ehbgiaXglNlMEIGaM1/PJUR7qVTkW8BUXWJDh2AzxRntbTBvl5LPPJqF15fRIc/Br
esWhvMKKAcM15XZKp3AocBl3BIOrEcvQ3prQbHnrW/nmzoyOxzr+5oNWMxmLMIpf3rsdhuhLwlCu
kdzmQUACBayKSVm+F8BcpEg6x0mpjzy5jBiTVVnf2BSkU+cfqZobW7qI0TeubDEe+pqNJ3L10WnB
K+ahpsLUMNhcXMjrXLGd5Bdsh4mwY5zVkOyvfG9EZrYjs21UVEckfkqMAZB1eKASIijthTWkFe9r
Fir74A8fVl/U7tTaCkYz/m9ZYlkQ6zpmqmwXTEZvSjtBDTmFyI4Anvu4hugVy7I6qzxcHNmEdF7W
beAUNZgI4e9QnRMSaokhRUHdVE3pU1XP2Fx4xGqqxt36dD+KMsIsDWoiRJLTE2LgsJxZwpftsTgW
Z/aNR9UfQcHGdHhKqQyafegFAzZG0WP8335LfrcV7TK7S2dxWKqxeoSpkAq5OxiWqe7OSmJft7aP
2GZBEzw5EJtsZqTyzEHHvsjKnzuaAj2TmrnmGYXyEPt31JhrQDo2to2cvM0LgD58vPcjMJGkCN2L
XQB8VBZtT/H1OwmDCykK6ETDA4aAQ4LmQFg404yZsiYpofLFu8NCy1HYQXIE1LUe/FqXlIgcnu07
m5xeMfW+kg2IUxtBi3rkR8+TQCnHaZiDUBseRL24Ci3z6lyrW5SQKS6w0H02Yonw0cQhLwbAZz1L
Ah/1xzql4b9phJRT2zX4zpzQPMRS10c0dqNlsQ9mioFr+leTejthFb91m0U1wEvmb0r4xn7q9UeP
HFJhrEyHQ6f0v11vh3EbiO8bsdPPDx6OgLrdigJ02mUQgGPPLttij8uJOh0LMDoWNKQwdL9njEid
3VIiWZipYqF2wR+i/6klH6io8KVa0luCQw2nQHp+8FCZp4vZakYFKnGKU2osrSNxWC3T7zIsKpYm
1MmJCOqkJmXKsA80eMOM1IgtGWYRqkd8xTnmIcjDkcsHjABfZXqd3Dxd20u+fBuqmUdcuZCsuXRR
/AgDPIamEH7t/YMxNUB1gO8uQYa31xsAlX8OUhVZeO0r+fx5XaG5U0jpbjY9JrQ6Ngyq6GfHWaUF
eMvwTsw5zXJmrZ3+jRKij8oR/hWpYMioYAPPSQwoyAtvlZI+902/ZxSJZe8pU+0I+nd0kCTXBaK4
6S9qH8mGnSlCbpnOmK74Wam7LlLcmuONz7ySY6otu1yXeSVCt0XmeOte5eGYT9fUUIibmqJPR0Nn
p7ags+Src2nwO6a5gR+x6bHB4rYltKi94bUm4/KfvYtAKl094l29LZI28CEeIuTY/6ApJ4RWW69Z
i3jmyu32e/246mQSLFcwwRP8YYgiGF8jzDhuPDg6VNBVEzeBeEGfmB3jGIK4JwJ5/D0SWspLmTVq
UxT6L/yJrEzRxwdIe78YeOK5DONoIVb5ODl+FElBOu/J5b1nulN70qtpfw/y7U/gJcKZPmRINQwB
kuwP8Iqatd4yb/WiG69rPzncwBDonniAd8SM+POzZf8EDBt9G8pSxP/MuSen3N69ZpvuKuNg6RjW
x+tkw97y/Juj9z4GotTlE2ZvsDF5GVrpFs61sXcM6jjG9vD3FqbtfHu93PNj+Yrcm50qN1G7LHEQ
YOs/d6kUcQb+E0vjX0RDaZA1zCpD1U6zCascz4VQ28BQwzde+w9r4BqDIBmenSaYO2mMkWZptVwI
OEbXxBpJjPtIEG/UWmdXBt2BiJJo3pYI0WQ6IVnEF/VNrPmJGsVXzfa/rIXBKfN/IDXeH6nCNaOL
i9sT4Swf02hA8leQRQQ52nNhbxkugXpu62rLmA/MG0UKLIOiMEhXKmpaVJ+B55ZD0FL50Ag3VRo8
svwYepZqNQqaF0SOVWejmEbDek5nKZwzkVmkCnOCz8F+3XOlzoD+2PsD7kVL22uwBaFooOajX0/O
IPGd5QbjxjNu3MdcoZe5b12sfi1yUUgBRX1XTGBA3V4P33H+Ba4TvK5iN50Ob4r7I5SRbJpkpuP9
xfOZg9SJukWbso7KqAysvNkCacOuIPzHiFAMgN0phhN65vdAnfzGNxx1oXl+xylJ45BnbxMhGAH+
dlawlcLnBF9rxa1s/JixwD0eFeBhyzuE9HjaXF11KBKgyMNg14Chbc0AxE4AHUcDYjn9UcQ6Jzy3
oLpiUCsLv0i/xvZzk2y0RyiYFRn3JgtuZPMZErTzokGgIVN0LWgGbCEzdzuWoxEFbp0lHYVENbxg
08TvtOomhf9fwWvUTmWDDqH0p8Wf556xxFp0UJR0hCShhdAqqgvQnEqNhfRJP6FJft3vAxzs9au8
jcEAARaV3CWqls6MBuyoZJcnMeopbO9cEKMHT3bTmmxNzpx3IdJYUzbxdhP4V/kLpo4B3LFyinr0
fqHnHZlUSalsvCGDvgAMO69rnDDpQKDsrjnbvLFvfO6NlzmX8nDS2kiRX8MQq21aXbGu2lmWm3m1
geewUbwblHbd5cIHjwx9Xu1KMUIXhETEfgvufN3bevY/D3EBlshq5I/VmxOzw04Kkyt6X+iZH5Rf
/BbXA6aVt1TwijBtWMSmLKrGlXT5O6booyiEN+y+QBcarNsWnjBnJh37+ydPG7tKiGAnX4OTEJvq
HgOYGEewfYBv9MOhdR0Hf9TuKJ7nvZuoiiCQUH/A/yLLNyuSSCzCqTZ3kaDUxBhG6xQKQucwnjes
qcgXu+Rm9PRo7xCnCLaCB+H6/NJihlAfukEBWUjzTt+AhCKXz+tCJEjYgMcUPc3zu4575uUwRQaU
SYo1uUHqt1ldU00XVXBnk0qX1Fm++lenc/CcmovUutWK40ZyPoBhfBLvIUH/nxBxQCFMh9wQqnzE
ehkNvYVx+dw+0bX/M36SWWsqFIjWNbps20MKJg0KSzbGxIOcVHFn+i1BokSW7lx00fuMXOSb+Sfs
LDfJe3+rBQmTTLJmqHuEvCEvC+UclLf1PPYIYLsVdghpQ6FSsz2ZZUt8FzSIyb/ePw5/k6C1wVo/
Xqia+ZgNGL1TAJ7HESZ88EKzOQGuWU3hGmO4IpyuABEPVHXzh9ZiEVOM/uz5HMp237cIU6A1hq6U
DQV4XSNbyf8yzWaxZLA08eNE9zkdcXuu1Ift4//vDQcwF90i81cVzpT2BxKV/PjIaMDQP4wi5kNW
KyTQIfqtJWp4wdj2Ekcn/10VieJHUqnKrtI6fSUhEnAFtGk7oMScnSFwg797kMRwD+6B1fh6+DUJ
YgDMJH+KmoEj5pvk/CtKFhooQX0etj4Rx5SIReFQJU68bqtAcxO2Vqa/B5oiPu/Uj7hnoYpI5YTk
xGioEJ6r15axcgauDylNy8E2IdWHQAyXMBVSgtvTGoRixIV0iB/MSZcRz+CbO+eIKfr4aRjKxv39
Ewp6w5mHocB58GuDH4OolVLnl3L3zhuBqU/iluzZ1n2cWWN/Ul4hN3Ao4ZnwGJyugG5MTV0Bypq6
yVw2xIyJTonbrVB49YmPR9/gPdLB9O75cIJCqewDhVp0YPvFATpEjkPNxzjI3g95JQzyFP3CDDrf
H2LDFyBQCPgmQa4uI+P14DMRhwltf/C1AY6bpPsRBL0x81FpYVE1cBHc40aaJ22HlNm0FEmm0gyC
26W51lCWn3zOj1u05Jl2JpVY40h8P0iDP3QdhXWoQocyMKH9rKiey88qhDQfHHXLcYlfna8hnJ5H
KIlqAPl/CzhRkC+DmZuq6QTuDRYMUc0Uy+EbqxIbtPDnOWJkOvxkdgRVu86OA9yq1ifb2Zbwyng2
CgpFRQCFXfrWfbK/qYzg5acSsM/9CThElRRSLjAlsYvOzzZpN1/6d9OhxrSUUvQ30FxM26Z+T6h9
bavtV3qtCQNck9soR26oB7q/gv1Y88xjJ3j26YE28cH5CEBwsBUau+e90VjxvzNXoslsZkL55zbx
OPGCW1JdUr64Tj5LG/vjCllWqTvM1ffp8N/TuOlBeQp5I1ZAJ0WwYPmD1k26LYs9OEwovgVaLR91
FeMGv8Z2N0wBTcrPrP/uYP6Sfmrp5RI0Zph7VriEe43fHrtR0sU7H71fo+TC9DFM8XWYXUmc2e0z
Iv+o7eOqUogivdVKziVrtsnWb9CmQOcPCQdszYXx3DpuL6oAQo5VK94RLz7hczLDB5nGi0l2qoBN
QK5bZydFjDQfl1zqWw1QhdpKPFITISw//Kiofci61tkE+1dNL7a3JDGCX1JxtatnPNFsnfQy7wUI
l0PSUnGDqfj6aNBR0ObYbLth50wZPrUJA4zl9gfEqQwz+0RsGedWsbTW7++IVbgNWEFyr6De7/Up
oRL5rgu087h6H1tpnM60zbnOvwz8QSP++xGuaLNOzfWFbxyQkLVfNckVYmjmSWnrHAivjZpgMEuO
K1y8JAN1PaschOugapNqu+5J3dia58FqNZ6+l7SpdsXj4nXbWgUh+MPcwZXB15uj+HUm9puTBT+J
ErHzUZXZ9SOKnZieEz8mMvpTy+R23FcqncPh82SUIreEfDq2Vqnzra1EDha3oIpwdkcRYYHk7QIx
+8dCvar2Ev63Q/H8+iWa5aukrWwzNCeEH4tmZV74FYEqZ0LHT6D3i6C/ZPj0hdZLQoxdCu36CkXL
CTAzV6GF3aODtb9NbFzlAiDCxwYnrqlKYXuWspaLtyujduojAAyJzj9pVre927tvTT3Hj4h/PafR
1bY8X4jLc+KIPNw+kgFeyl+GDl1RuK2T8aP8cJchXzQr7+t/Xp5myz6Iabz043dYVQyxB+U+DED3
xdi6/Tw2UMMji84m6ZInSvQXsyePqcL6uShtM4QUdRJB6T9KlXdR0r2ffZNLOIpBgJ6I1qYIDCC+
fCO4qyQMIr2LL317H5WW4vvSJ40zyHqL5LEW4E7V8iuuG+e4Kk1XBpMV8JejaCg6cRI9AL1FglHM
I6yDgKQmYxLvvpC+y+ulQhUHHTGR7yml6QYKHWGA9I58XcEdmiwuxLCqXfB6F5pTuD+8WlRtspWp
0OUCZeMSIRgDZMfNuqYGQpFMAXqPNGloZaHOx+bSdnzk8PJGokZOwnufMyMcrs59RPJNIB3zGI0Z
IbZskZAQ4HimM04y0F8G/h/76LyZaYA/OLRoJajrYpBVNU4pMpsX/g7Wq0A656XmHCZVhU0zvKCJ
dfr/vSFgkuJwT16YMue0epb8u/He76A2AO/13fq0ecJjWS6DYaPJgWQyKc81ja8/Fj6V1cxk0EJ4
cC4zx7LCkBNK/EEsgvHkYNqnOSDnqvvLphRQ7X/N0139skMv7vPVSRnV2C6cqkuaRpWswpADnag9
ydlPZtVmK0JICjE+hQib7d9pwaO7VnJUJYuw5cA2J/kTecy1peJbW31e3BQbv5sXUf3iZxhZB30x
TQnsfWHyBHVFTGNNAdb8hq33RsYWpXxM1mC9T4VLaVasakjAtM5LghKOo1H2AYFJd6pj4acIVmBr
Y0Qn245Lm51vDVGShgu3J5ANCnqR0gDmXXAvrp09pI1Pr9heyCqt+/EU7qPlSEcadZjsIbQcthut
NFMxJC21JgEbgejaglE2u+/C3UjsASsl4H/9nadzQsyvveW1re+mBIKsg6hJ9PfPRS7UPBzNjQhM
rKOl96usjSwToAGvfnVACprzXPwM25tvFiL6l+ycw2S3jEJwxgKA/5ZdHLrd9/kcCKTscTEFV2gw
OEZb3IHuiJmBGwWqttBbIuwOB3G2k8Nx3GRjVjv/9uWPa/3BLYKK3iozF2R/FfGRYqwQMETuyOj+
+P7v5Fu8XuoTaIY0icCgTf1omxqmPfC9rqkUx7kxY5ofwD26Z6PZ05xlm7QCCb9pGD5qme70pGnG
Qp9JVxDG+DF+wDDSJvWQoH+b9kAduWFBOEca5/XdbMP7q6MUCZ90Of8psiy5yGE+Hc7bhPEAS1gy
eTwBFr2g/dEZB5NAnPlDrTu25dWi29lqZDUz5Ald1TaYuf25zjIdQAo1K6rciVVlHaENAA9qz+4Z
w7rVI/Can4fc1m/YD/PV150BZ2baMsuY/fmnk52oIinwnBnQXfMW+82f91rpTiguvdvDoiWJtdLH
sDWn3/ueQjdNsf7EkMkyH8jmeVxdZ+Lz8A/wUlFQNvXlgvKdqF4vklIqDcR+kEkUWvpiBV53mz8C
6zeXplHmmSnxjTeld68fFN8NEp+ATzB/OWUgHRhj4jqPd3xMg/UDRIQ9SpI3GzcS/h4r4dSw3+g7
qfwjT7RruGQbScp0EIrJ5eSbFZmAuoHrT1Ql+98/6iSLz+JXpiZD9Hr9q2AMTnLdzCAr4+0yXTMn
V3A0AXDYaAYF/3OHR2SONcvrEMmWaAcjwwNXdf1XFsrCMo10fZTiuSidaKCBMbmdcqW9VunFrJy0
2cnGuLkKwHZ8nxsDrZf+D5ZjrEPlFgXTShYEjhVmQNu8PLyvBPmpZuwRCqKBnqktvo9YiJyf9jQA
beoII13iWj+nSbsCxWz9tB/DZtLyN83zNINxQxxcnDv1YMyKbmSXYNXcDCdg0FbO/ZcebqiX0cXm
TlJNsdaDoo+Hg0uTym+pzadtEe8jF1hSm1rDTQOSp/pgHZN8G9KFOZLZhK1WX3yIGxcOMpueCMol
N9YmV2B+/vi+RwEX9mj+EqNmduizqXvwa8MuoUth+PA6oPIehOoSSQvNWenaYKV7LvSCjV8w8eIU
c9VktshfeLJCCnYhFOn1ScfT5fDeOez0YkyAcvOOh2v4HSZc3nhFJciKWN/xCOr6pNAlHFeAjy+I
b8WMVE+SWBwQB0UGxvb9jV9lKh8gUFFZaahQU2WlshnNFuSgXmHhhF9EQnwfaMjBrN59RdHCRIif
lBMoTzoEUj1NKSgYR9HO8hhPChwkBnnijTTs+BQ/LmqfhyvuWroHuu3gMKr3+I+PGf1WbdPNocj5
nHaGtKeNxk8u9JIQrm8MFFdsMX7LVIsDfB+oWj9zRF91Wf988LKPZUVlqO5+JWE2K5Czdg0lP7xP
Vt0WoQyWtQX9iwH/O13M6TQbpDsu9sHwVT6AGNlXsj+83gNlFueCdDZrSKcj4aTABE9mt1pnMFB9
QP0dZtfx6g4oSMaXXdqdUh7FK6xGksswkJ0ov12pQ7+H1mm1g3VQb5t5LIVlpUW2VTLMCwwyIKm9
0V8P0Eziu+R+z9B5N7DNiSTaXVdyOfAdvrjeOadAChkWEzSbCrr+vJ95t6c5wtqQTIPkLbqag3qy
a3OJyfx9kfFt44P0w+Q2BXLr9GrO4Z5bQ37YqW1Xu9VhUr/z2rkNdll14LMMILHCP8loySmYNBX0
+yVqmrn2wHJbwJdZcHyHnVC0embQP0Daer4NYgDTwLBy3XOAr1aRy0Eu4cT6P99p0BOlLApsaicl
j7jQtnrE+vptCnxltNXFxxbSltA+ULnSun+KTnf2Wffssg8lj7Jn4eUT/Uql1SdFO9QI90jnl2V3
71+NFuQpKY4ReWHxz/qNTRe/5g4dsjyiMND2Hyt4qS8Em2gjZQgsZGRxv23HYSfqY9Tsx6WXaVUK
DIz2SSrfd11s/WjC/ZRxN4CI9UjqiesPbDSQMuCq/sFGoqlrT/ZVEa/BZcvMAGXalMPbeC7xzSM3
DCCNmchfMnCPWFvz3M227zQVIW7hFayYmGOnle9OYqU51r50sm6IgullMErTvBKTgZ7DXx5rLAiZ
z0JJVOqUkLsOqOD8s8Gao0BPlWV7xg4kftA4uYRgoLC7/wNjb90PIkaQf/+zPInZR59GAwOCXgl1
qpxWz4OftFLzGqErhf0haAslM5Ffz2VzsqUYCO+N4RFf9ctenC/SEgcQgCIBNG7GaGMP6XsTJCn3
dBDvCF2EVtRjdscFgCISZfeC0TwcRW0oLWCtsPKQhxxHxnmI7iArJF+/eKyMurYERJGxZHvIcf5v
HPLxgwxzlhLfM+3DmXCIs7L844ZnaUuvbgqmQqcna9pCVOjXw3yLhRVJ70w+7CB47qyZTXHvWadr
ZiQPaRweinot3IqqAO721bOQdLQuLX8tEJvwRIB/7UUBdYFNrCVSUCgXuWkMUBtcQGeH1qq9cGwb
iO1XvNvdtsysFtmgOtAxzWhms0Ev1oombX4GzVTE80vMIyczkJjkvP5BQXLFJVud4Hsa87pbpsCH
tEZ0CPRahHWDxOf4YAEcgYxW00Ek2/IIvOADxRHbkeGNUGs/Zj2FybentftiaMBVvtEg4kvw+VZO
GN7U2/Q3SIknh/pJGnm93qJFUVzy4jbBafbpSRewf+yZeGRDDFrdthwJoOT0r1oU2q4QvOn21age
/Rpj69h2FqlGIZpiCStTP6/h9+bfKH0zyNiczfpe/lqZSWdOrU/RVAL3V9DEOVTPyY65PQPmCBFs
4w/wv/549S7KdhdXVYWrPMBEeTuCnrXX49Un7S2BpqsEWdOQIiHFca6wca2kGU9f4MvVv1yKfS/G
rwoz04or/okUlXxfCRWmD61wdLYDlDNCpFzk9d7Jx0PFF/QVlSh+onHZ/ZJaTsgvThYsg/k1qeiX
o4DFpxhHS0eI3FiffoUamL0u9fTHdxEutl+Fut4Hn0VgTrlIquWH7+exfFr6ky6gwx+XK/3lS/Yg
+GhoR9Mfnv3vmzcJ0gkDFEymU56i2/NwRtPrCkPfoLFzqenx4bNRB0IzDHbHng+znshKVOekBuJQ
7xQTGAWBqdnexPktdFZJh4yilv1hw1hoZVv9hBB5wIbf/BClsLPeDyyj8Lewr5q1D4AcTS5ZJ4Ev
rR3vRYd55cg2+qnEBbjt8jgW7OCACikaO5D2FyrLDa8ocp9AaTcLT02J3MehLxgjmv9fB1wqCwj+
jsNhUbbcAJT1n027F3wST9wyUJBZitCKTa8mdsNoiy3G/Mh2HMMuV/8zNnOIaf3DxBDQMBFvH2o6
OVYu7M2uD+r7UMGuhLOVHuzCBhV5wHqcyDsltkO43HTcqPY0ERiwfNt7AItJwkUPM45x6Cm/AyYq
B3/AoYO+4ReTE4VRbGRrxuBFYy2Dy5aCi36Nk1+RYCAEEKFpg/p3t11z65QWmur4X8TIfRKOTbNu
YkYmHtODoGc94gWcrEjG00HfO1yY6mUk9oZyBdNE/hb0Mv3Oy1/mLp0bLoE+NcmoFenYocCEiDT2
U7sKGu6yVgmGEDGvKIdNwZPBRZWVEcpRCiwPyc00QZQ6ZJXq14ZKAXOLyr4OugSHwqkjrXCaF+FQ
rwwWOWZO6QLnGoNGUuOtOIrzSQjNGM0qVvYSAJtGiJ91j5mw+Xsga51d0Ks6kxH2srM9mbay1R47
ps2UgXCYnnnEQP0AOwLgaAo0xsWzUPbUNpy2vY9CuFzlblONTmNkmmVJiGyroayHBsTIeA+Klyr9
02kGORjdgKpaFBCQ1CD44Ol92VIZs+VDbNgq4HS/1FCVBrLROEVtS7hTRCDcKrhZc3vbhl6ovSC+
DWfqrGFODrk5RaVttoKRV8l+hyDiIO3281yX+sqVqWc4/t7lJAmfkyUJ/LwotU4SHMyZTFuGtQHI
FOE4hA21xUkBnlETPDVI543rCDyelPycA6rrPXo9STqgORfJHxZkfmeO+iTyVgfUIeC5ECLoL/ru
NNTknlcowd/GJHAKMckMon4cSpak98i0nOBAvVGgEsA8MCu1adtItdmoFpkf5Y20GqPIefuqYB+K
rmFQVnwTdcw9TLzOODtZAEjfrYd5nQcDBscC+Kd3YDz5fPZUrjjofH3APcESf75JTsDHRIfie6Lk
7mshbbatpRBD3ByOReRTRyGpsb4Ke7yPYaV7BinZDWVckRzYf6XsWxiba1Ol4DIt0Re2JfKHBu8e
OiBgVNggYb3Ev8i1L9JYlcrzYnE6U0qvWNtPvTEwI2Hu9GSU7njN9CavJX20ePX3lQKWe5aon7qv
U/4q2/N3r2NTa/lm4BSGEOPhxkPJ+smLzqrqGpcY8c04jTYcd5+swszdDuD144f3DF3LGJLBqxav
WxOO+wdTTCHeW06+AS645SWJbBYGIRIWPN17KlUIbvcU8BDgCFKr8TsJs6pA7OTIMYwwBq01mLzC
eiJ2bzYwQxkSzQL7Xv1b7Lsn11kqhOz6ztXeczkXuWi0t9nkFAsBFQkKenDyCrsmej52nJUzgrq8
KYVqqcMl2/46iNISd6/0alosxdMGmlnqj7wPWyDsWwpEGWEtQZRtzl9Iq45QqwxK9kZ1HJRZ42Gh
o7X17HB1LYoE5PO0NWhop3hAvtO1gElM98cPFOa9GqMvQ2SAxoSNzOTlHti8jFyZZ/z2kkjSd5Rw
pyQD0kVYtFvrVVQ+71wCSnvpJzkobjFcmY4mGnVKpyzjEfEGOj1f1FRQHCfqBjtVA/OmSFFIyLa5
xmi2bdM29nE71EobxC7h/L0FOdSa9A/aT9OrLlXvj4Gewy1IMSuWEQjq/qZLPrzUiwPQF/NLVviu
iP5D0CDkZm/u3qyMzL2VmPxx50Ckum2WSLQZ2T6BAgOI9LTusBOJNUW6/0xRlJoMPkGKjmfk/QMe
FD0JLLIkai0CAj2kRAGMUatN3C6QuPnwSGGd1GeUEZHkWfK332JpDaLgK0YMxfdHelcCrdJvLc81
eOQl1EXlnFRsbMZvqxVrEFwDySnJBCYvw7n10o+Eb0ZsRDYyRtrACFaTHLGXbXWjKsrd+/2PoBhf
7KweeSYMxoIL14f2LBqeO0d1uk3c0K5bFLXw2scpVq6usyX2FHNujBwgTlLspUMtflwODY7JPISz
tc6zoail7fQrWWj4Sw+HuU6zf7NIdu1egZz6CJBeSRWdq+v9Kms2ZQk41G3PIUZUOZ68Dw1Ngsga
25rkjcsB7pi4qg6W8kRqZ5WpElOdLeVxGVJK+DGReG0X2Uym+HJlFYfajJ5P4Q+yLNV6rVqBzszA
T/r20IV4BFueBpHBFLmLjcibM9eEBPI9XXkSBgfnNeG6Tdd7esUzqY4+KeVY6o4izHw3WkgTtoRE
OEF0nDeofqCvzNZVpcBiBei5MUCvlxnw9yMbzliKi+mVJBB8wsITptoi1Ok71hLmrDK26MVND7Wy
uVWppa7caJMB4NuNr1NwVvwx7aObvikpRrvD9AIW9IO+KnXnTXb8dpe5lzxdYxej1oFuem9K/SX6
cqX2Mivii40avCvGjko8uXWlH2JFbvK8fQDiWeD9vIxlxzMYtR1rocAUsKntlCzerR0qSi3jNG6/
B/7sFdfgnOxaqt+39RGj+Nlon444KfDslXJr2Gq8NCak6rW3giwoCe4bomnpbhvcsnhGCU9X3Ske
85ug2cn/c0+XSfoHBbMkVQgGVED6QOf39pBx4nx7co6k2UldeNthEbwmpf/BQ40YnJXO45k5qH0p
biXdQDmzEorg2RZa6bX8cwoMW1byi+BoCC4AbHlcKTtSOLqiJ/bqorACQqzYsuC6SmM8vKkt20pS
faip20/Fcqx9EtG28BBdIi/yyKp8s7jHxnzyMkX8/e89/QWvw35ayJaoa6PS5ODxkNvOWgHpb3Yc
xmgxYELCg7Tj5bT2ZHzF3WzuUNEvbZjOSg+4G1sE8XGfhnTGnNIetgQ3GeMt1OubNNK8zGCdqMSI
S8C4TANCXzzK/z4gccAVKM+ez5hAXHAy0yoTx6QfCHNMx+xAErPC6HflgF3u7bjFnZBwOuxhe7jb
VZ2n/cfhXqArvT3h5gn4VaqP4QnscTbtOzLXZ/9PAfSfjjwhhuRqac0E0Y53WXKv97CHbD+8WT/G
4ykHNR9cz8PwPzTAqXax9alOa2bTx1n8T4peKmqzeGO2YgnqQPLZoqe2PWofW/hlcYftluLYcfPT
eqFJqR82pSdv2mN8sAQoZZrehmIts0BXsLLx3kXd+U1F/6RZC1tMroB2OiflxZcT6s7bDh9Y/haj
SBy6aVuifyEpAwMNGh/kugYCcxOBqxf7VWIVQACRVbhFnneb4oJG0HM4apaPu/dfWaWXN53EMkEd
hS43AdQw9liDvZdWYbXrXLCRWFHM0SbvidhBnVY5cz/eW9ZbQ84sX/o20E8fi5ZwIiinEBI3lpwc
vW0PczYbbqT+WWwst/hdYEw/iIjHcrMRJ8rv/UU1JTPsDyjAdxO0pLACwo669h5TKlROHZyZNhra
3SocvrD/p7ZgCUdE4aoYTCeW75HMl3aGOzzQQ9Meoh+hfZWmOyhtjpeQWY/FvwmX3tmGB0GmHF/U
9VM9BTY+vy6BVufW3sVE1BBzJs0LDUNLK6hraH7nfR32QUAcZ+1CK591qXWxYeSXHkPLIPtECZyk
4DM0jrAyYTftk7w5tFNRmWQgLxdvVGgNcT56inwFOshGT6ZpvWZYcWuQ1xV1J75k1xzQNwdot8TU
AhchkMzBugFcZf+GE4mwoWdfCyp+Pcx07P6J6AQePiHjzLztn1FkPnZY/pKVIr4z31/enffGCOC3
uYer4Du3I1O09/fV4qfIWXtekJbM+hGuraz1hZMLR+wKqECKVuJBQ39u7IbZvZNaMA8reJsAKgEa
YNj27P9U8/osHDdyAUAXM8aYD0nGcColfvyKP+iT9alpTXgf09BvzDwagEaLYHXh5pPhG15I/obo
kG0iEYzP6ohQws4r9LQmSOYyfvuesqZ6MNNztmteyndSnfjfJ7Qu2vZdNTgY5Dy1OQBDW9UgUJ0r
WI0w6OogAqazXdrBSe1XRlRWp41IPG7+hHM0GyaNbrBjkl4/LLxGO4qXe1DpfUKZjEJ+DLUtizpz
Hk0xAOpMSB9MgL7o2vglkzg0U2iLzXsZZ+VworYiCrA3Fx4ieXx3E/GBlK6Fh8Fag0PAeq1JLDjD
ATGyZpuKx/cyI0Nm96DhRXg6iu4fSQb+VSj3bujKnAJyPac70VWEYFPhCBG9idrgAnZREmcqgEOt
cCJyxRrIGps+URL7iciJfSP4Fh8uWf+Dv+2RzXw63y6J/E5Vkj2XNZnJ48STpoTXMbAyZIOKdytI
VkNO7scXr8D4uz9cMIcSvjF5IcO1ju5N2Es0NwjrGyO8s4wcinBqsGr+dNCSNRsKE1MVG8emlCYq
Sw1KMCS0VMjIIB9uC5dCwqE/6Hoh9vofu3mXQo6g44qmS6d9UwSttD3o+ciFaoh+Rra84BG+91e8
hOjSGxorIQbFeUT2iwLcvaeTxcKiRnVgIq7IGDwmciNxRNtY2cRfX+hJ1c8SxE+fFpG8f4Ykdw4U
x+BZF8NxROekH6+urJoBi1nuhHHGymM09wysonjJy+TMZNTmkLw940QDzM6mUUuK7RSkXB+xDnk/
Tx+iYA1kYkxrcrpSj1xZpVmproQWReT4eZNte+eNnCmIgnb4Tl9XfVk0xESKtUOkGvJciE7o7Jbt
0SnOkBjIRTMc0WTMH8a7ERbj0TJ0c5ob2TTFYUn+zgXhkrUeGfp9rd0tMAI0qBxUX4b47c5aW+IQ
9ZXbjDqKMgDqk0MM8vDg5zLzfEC32945zCdvMV7qJmWk/MkAWe0qpPCJjppnid5QFDnFK9VlBP8j
QG7q4rRZUwp54dkKzGtKMeUMEwoUhcvPUT4lKpaXxey3+llyrefrjoXTyT/Sdw7oIqZ5BruqykUu
2LNTnOFDBZxe8hCiHbeOUyXgH4BbqMeuUYnqwG+4LCL1ei+JZqvkRNVPmDvgz57il0OWYqjft7uG
1c3VzN5YQtg2pmgOgkTp7czq59uLCvphXtl5t+ZXFfgP4oCe+vwOWxBqOus08phneJzp5rz5POfg
opN1n5xz5G7+pOhWT7bRjvj3DW8OvbdOvSuyNmwviWRq8v4lpc7rKESn8dNTjUnsTDFeZDvwSoC4
+pMucgqm4Th/9gjPomenC6KTvLOWPT7qOzX5J705VCU06uLSb6MUcTAPEM5zxWyMbGLDuEGVXI/X
HrZY6J0yiq1+ylRuAtQ0yIx8o0sNioa0jCUJ0Ny2QHtlJI0ueuB8nRHsrkfnnZkdLtspGqQypRuu
6wlqueVk/iNYmat85f/YogEh37a2xgDgm/bu/cpDuK0bHkhbzXfJLVwniwiWGGiNwLVNYd4sbAkX
acDKcnX0k2CRDi8TOUwP8cjs5tBX33QfvXaA9LVLD4obz9OtxvEIVAHOBavBFcw5WIZE9rw1ZCmZ
8S95Kd0I/aKCc4uIHsSRDvHpyU227nmK/LFh+U+DNP28p7tURdQ8N1R3x4nSyeUunJWcxIc5/A8E
4nkZoiFGbHjCNBwXxZzfrzKs1Jd3GRk9N+Ooh1Rr4ClQxHRUx67WTaLJ2ygRIQUXBjoZGCGwDtjb
G0lUhsr+xRv7V6XtOb59ptpZTSlN0OcJ/wVyEVqKI9rNDkzX41jFo8gfkD7PWEVNDHiuNLkQ+AIc
ho4+CecDZ/HYnOjSCf0Wm6X+QCxpDDr0R8Fra++5N7CpHDFBlvfNRk3WxbbLNILKKzw498iaF94M
G3PHABKP9tTYzuWKiINte/UktcRvjljNQR4bd7H4Vq5C+gV5331xqJGnQ3vImEzDTqGBw8sJlOnT
LPt+mrsTHZsKt+Pu3wxCV8jb1+F2kNl2DXXedniAdMce/mXEe3PkgNstuH/Q0ajWzxO73CMQiZyT
m8lhZ6pdTAgPleKLygdsdaAWeoUurbJBQR2txNuIVtgFanjaqy3t8oPkVeYv/7fLnf/qJ41lKR7k
V3j4mRwh4uNpz/MHxQFkJbmdPvv5s3+kTLv68J4ZGHBpJlPT9qZQrY001KxM13m1F6SEIj9mBv+J
kl/z4JWI3KnEHqoE7jme3rG0jp5nUIZfcvQ8E16sxbpU1sW998QdcYzqDE2sX7fax3LRQdSYhz1T
ewFacYBGD1IpajYf8jHUmgrznZhxqnQuWue1WK2bUAK4Vg43i4HhImBAoQe1kSe1zAFlIlL39+LT
BchoVC4nEpMrGnWzodEPXSSyhB0AWwb76aKYbAre/WXC8jIKuh4jYscoRuRzeQvVSzaxtX+a0/5d
f+IDhdzzMSVb/6eIRVhW/6odgHsy+TbBEYtvyzawWVfdMgPAfM6YOLO1PiGU+6mhBMTI1KFSrpWf
fpa/KBtE6QkyCgY/8QI50rZf/7HOj6GyK+jqX9uhATig4H1UVvLQJDJf700czEpFJHrjyTCvcwNb
kgqBa57XlIbGRS8Ot6ILxh6ejcLkGSDyUaFJ6NiEJhBSLtygopxX+QI/glreSmJg51dRL7qdtOyq
u4h4eQtSb+esVrxj8TsxTEMtFtL6weSTsnEa0jUkqv/bUuKOmQujtBlx5LvL6OVXxqHaKSU4URvE
qWxEdbpypYbXKlWpvnmNrVA8EMmL034U+u9iGEiVuywEx9jmfNI/Xa5fzX7n1uAC6fMSSKYz1vUh
rPtGwgGpoLDskX+F/J0cMgIOwucidMm+UHm0W2B/2mcPFGPBbrjpbvwflJtKyldcI1Ny/O9mMWHa
240zTcbH2GSvgXgoq32qCFYOxa6ktMMhxKJfj+7qqA0a7KKhw6v9IC21UFh7Yh6c4EZ+1iaHQ3ae
rZs45D0keeoqhHlhkeK3dogaoYS98wRrpeSoOIJdBXTsJXYgEHpjzuy6Jo5vu1O3Il3UyF4WW8Zc
9yAzTqJAtREPTTJdntZPs8qF4ovin0mLmS1/4x+oVnKlAgsLaSvwynsWdsQTNaXO1Dj3EeQAHer1
9DC3KWOp0go0kGWiv9tJUDQLtCTv8H4THHzIF9wYQdErZlp/OdHJWlAcCjkfATnI0jxI8iAS6nWO
ERMPytO6llRIkWQWCiJYHlPxUmMOafUeUl4SYD8CmsTelxBwXEv38vSVzWYOlUoCX1JT3lJlSy9R
eggT2zn4CbfvVYG6IOak+68teGQ/tbzdev2KwupslR19YuSqSaBNhylUkegjHGgUeR8z1em04w88
vWaW90VMoCpZt/gwM+3Myhc9ZFL9jVgy602TquXImbkLR4a0b6jpipI6BoZ6BESSu18bpl0S080m
yjpX+eNwu2i5V9g40cttc2KxgjpChlHnDq7nxREwKeLGazGKTxsWL178ZMuvgD22qR8orvWQcZyE
bBBALCKffNRK366TU/MA+oSuokDGHuIVP7erer753f3zkSDwWcyg0n4CI/oFQ89npo4gqFoDX3xw
7NeuK+d62EsoOvXSmiFuTpLTomxvBpAZ5Br3/NWy4jAJoMzx2E+PdB80UO2S7h/MhJ9KPZhwrQD1
bl6c3bQ9TYvZVb2TW+/un4T3SyVu9CbzSNZumNoPMwbuCZz/vynAXO+fgWmsfK3mYxzow8oYr73t
FCOfrd0Y6SASJ5smVk4/qwsapL7c2jtcNLLbSHYH1lIQNHTdcEBeZPDsyJYnkQebPbvNXFXWFowP
vVyD/upEEKKwOdla4UZDboS2Fbgr1xTFrDWKXF1aWnDzvMx5kLx45HEaugwPau7CMaQG5MpWrhMz
jQf+fTFqlz9PXZYqPs+pWwC27DJsK0ecxqHucwtYqJ3D+ixYzVF16NbmvCOacNK479jG+SMV59m4
7p76pgeYAg762KmIdm+hIV1kmJlLvpdILuZkHS6MtOtVXqB+hPgn+mgFELLa920uKdLqdB4v4F3b
U3L4zM2Nsd7OE+Q667ZR9y/V0VInA6Jifd8TgquqaffdgQ7d2lDCcQAe8goQYbBTLDDK50j1zbz7
N6uv5Ef+xPDIEM5dkqhNI82jS+IyAPMW8hmS/jlSmGJ17Z5WoWd+Nb/HxFpiITcTKclFrQZXZT70
QIFcYceKrQw0ithxeNgyxSAVzmft/t1/IoVDve2llQPm+BP5+9ieilJZw0YfPL2r8bo2CqpkEqv2
9i1YkKMkT89NVppBXfveJXaChRY/hxOH5oQ5Wb+1PmfnD7Eh2JJKHg4q1MvPbetqOVD+Hryv7XMx
Suex+US8ONzmA6uM2seH8xEgM8fGjRBinmd7EkCtrOOVf9sDgk9prg8lK3tco05tciGmC21b+lF/
zzo8RALjEz/QEtp47KGb21iofBJa7ZR0tg22yB+mcEJ8cn09yHyoBcEHN4yC9Z2HTY1+G0r71fTI
gxiNLmlrqfxrTXq1WU+isOjeCNvcTPm8u/Doh6hUbXXjfkmMaY7XlQ61zVr3sPBg8xHdIQo1GRMv
AuP//3lrKYLiCuuR4JXhEn8uwk5qmMplSiWqvnN9Dxin+NBVqCD9Dlhdm0l3wqYvPlhUICbEvZKH
g4tZyfMn4iRbOmWhNiKn5pJ3KBEmrdJRqzubUcsDcQuTObGcwlsLAjKdv1JfrzUXbRJDEp/eaOWI
i650Ug3t7l+kHc8As+ke2WiyxUFQd7oun55XVD9+ZfXcQ5ekKIlZg5PskGZxYR/vLCvhCxqeYAKP
Vmthz8N/tDMM8ma3ZH5ZatN1AqXvgmOBbdXUQ6x0tw1pNJEcPIBOovmJ/2oMxsr6+vgyLW4AnLYc
TGlLreswiqsOdW2qObozDqZDlldV4yqPHNgDFXL3Q7gFDybeQY7ugZfiyz4RDN+IiwdpCxt/cqXm
XuST5yEVddy5+okpM3XZffcOonn4Uo+nDnjXO8XDw+D3bEMJQvORmtvscaHk9R4IZgcrEnkGBb7y
fxKvsS0GrvhFgO3FMfpIndAcftT14ViVFoReys93/eaSE67vb3BkGY9GE9gKYOSlQ1NdpnrRy1al
eaS7q2pITLjMALytANPsUKXjFzfC7BU2nyZUJVCtuYAnxDd0DRjz4osaudttwc1naLwil43h8ZGo
6Ve0DWMkKPlhPtXH4mv7wgVMyZlgWf2/3FadP68QjNYg/hfkmm+Ck+SswQQtA58darX9klSbwyzj
EKlpojtyuX0X6QbEk88wixESKO1TVVpx99XGcfKj5PMtaA8ugs91kgQJJOQSVExfgB6QRgbp14Ub
wTz8OPaYyjy4put3TG4PBQuJW89rFf5ODp9JC2Qto3OdivRwJRCNXDfV4BChLkzHbQBEQxCBTmza
vlz3XUnHCQtdAyMu/mdO8gaiIWjkjkW2AWHxr0Iw+UqmlPoyPh79Ic05ZslNRzXGoVlWtwyGW/8d
RJPsS4hpHxmXsYHQ9rnheBUOyTVZ/al7CY9Ryf+MNm16QMswJ+gs5hcxgJ5tkipnde3/XKMCvYhn
ruVWVGRGe7QBZ+AdAZE2gwubb/pgA2wbRmk6pC2Hi53Q8QIRncw5cXeeeASB14lUUIe5uSc6dLdR
G+sY92W0RaBU0q62PM6FtxEIP7GLJRW1dABFyeObTpmg9cbc3HoQCpx1/346MaD5T5hMWVYPf6DC
MoalHag3aUl40jfmvgD9EKjKgQy6WOvNEn0juPULTBA3hRjljbi7SIz0yLP/bCJvJfzrq2JQ3H0K
lrieCY8Sh7DhuZzOwifyH6Ape8TbBI/IkJoXBLSxUvpXVOCuPKHFDTR3NdeGDOlQZhylf8PeF0Qh
3DdU4Bm6XkX0VGyjFWGaM0E+60CQEzWGrM2O1VRCXXjOGBRkLj6km/WSDgdLK0Q4Q6kdEueU/th1
oj5zpp/xbyWUGNaYwGwswxZhgo9RXJPDDxBZeGKycNJB/+9bu0AxvWZy0wgzPsIHmBSq+UvIAOLC
n0pQ5nwwQOQQBoHubWpL2nQR1DtNPCvGcZzY2o1V0x+Bm5801zIRYsjC06r0qOrZjk6QuovwGP98
zZeFpm0lheosdNaY1c/S3yrGRvc3HU0+WzEWdHxBu8nkfcGjiQ/2CN1o3CNaIlUaWJazYzRu3v47
llbfrM0xgrNE2pliZzcLHvbtPZBQ2UMV6U9mTMfhbN2kp2kOwMoKUEnTirNU7bnAnjVz3YHP5zdN
aXYrm/Hwj3pucvV3vW507KdRf4lvbc1r0U6ZsfFe0HouRdzwL0JqKGTftFqRtaezQMoc2wN1u3sG
gfBedVM6Vjk4nkH/yV4fIP0K1naQjvi2qclQ90dZmA2PQFm1ZhzogAOisI0rG2hLiTJGQcnseS7Q
cuwzwL5ZDEdxX06b9IJKQGhpE75yoLDUqdGiifEeOxoTgpxFAkY0asoOKx0OTRHpsJ5zmA7PBK2G
EGyPURm1KlTl2shnKFk9qrjJmHdeSohEgHdva5+gRciJgyYmPkD02VZR/qDTuX5UKNr7P3KXQCmf
GsyTpCmr+8rpM8yc51Q1d6ZkeI5/1B9/0LCLIJO6hvRajCbGn76Pxrxw/99IXn/N1RZuykhkrWDB
Vhs8yKQS5zYZMb/Zi9V7qM7Q1vkswBXWO/UsIFgEbn0McIHZZ6gn70j5B4vMzWRR0mf0T+MUqORI
rsoqZfW4XYdn71r1gcnW5oczuJo0Htkrr5rIH2kgsSKfRMZseXSf9yttZPEwXv9JezXZ0et5LwTA
RAmu6g8QjIbDvf71ADG6KojsrSOxoWWJS2KT9J2MEtMzSe/oLOuccznz788R8l3OmnNZlkoaepYJ
NtegqeWdVuwPmWPe2EynO0e5GBztl0L2i4UsHzfApEb0hmrh+fRX2XPpzoByQUutkR3T3JOgEhjQ
SMQMZxbie7h9z6aBIrfryZf/7WlkDq+YkzVGeZUt7hO7Ebt+7MEz255AA14TiURMaQ3bKnad6Xtv
lpKMk+pE9cWLHhvI9IW507t/rKcDhsvSQfS+PO2/jSlxxnYUHFlAoe60xoR8yE13sGwK/9mlsAV/
ECD9wDsIzaeObfoBGoMWpyD9f06D5OjTcti5HE5GBB4tDOdufcZ6CzH9sxZEeSd0iL4WZrSjH2FP
5OGNzPzzUx683t0ajKbkFR8jiepKTzfuVwgnuIbh3KN7SDXZVCByiFCFWPetjOQVgZaPgOgVxU17
gkDni4e4no0PVEItT85evKoW4koPKLgJqkBS1nUzkusUDhiU4VlNolNQZxyoGXDD4X+wqpiclJei
i0eUeEKPwfKgaxthdcE12XyLAhWUIsKMMOn4m85rzJkV2PezC39zgo82OiTHkWEiTS9tanW7GvkQ
BfM/5ZoKOaBSdP1ydj15HpiJWLlQNruChjSPfXCXVOQ6WrrTuReOtprVSDErcOfzAA8BYE0cTHkh
8jYo4Yt93C+RJ5k/TVvmGdBSOizEv4Cq0R0dEfG8yMttdhSXaRXDmWhNnM111Zdl1CnyuhWZJ8aB
K/U47qoyR7Nzmebc+KuIs42z9/KAnfJv+7Z9UG4YKQKWBbkXt0phyMlxLxCBzNZejVPmIyuw4DjT
FU5VfHuZeHoBfWHky3xkp+xchDBzhNn1EZhPtjq5MdlGpfVpuIxm0Oy/klOmzurXzYwmTS8AoC3o
2t4oVawO1vI1KsMtX2NaxIFydgcOnWvgB1AVk9CqP3HPrIBcQTY45XQccOrZSUDgpp+zzR+LDdxV
eqDDnny8Tof40XyH2+f5+PU+oOYuaf3KrLPNbztxwxQPMD0Rg9KqP6pKSW6BK0DTMyWgE6FxqxKj
34Lyxaj4xedOPaiPniKsMfEE1I9nmUOOGCSr9E5UH/68+ZjUo0QXSwQJGFsI2q+kwl2LkN9hzlI6
2+4ebE9Oe9t9XWyumP/xJLeKmvYS5NGwxNA67PtjciamhegqwZo0LtQK5i/QqAKGjF/rmYe7rdvs
XMw2iAOo1DOR7ylYLgf9qwZAVOoGFj6S6W/ml1G28kDzatKzkP3R6c6j6qVNY3o0tJmobKlVlsLl
3Zmci54+aK7PU21mvMOsDEWPUTR0kRBx9ufrAg+7FOIwUGPGecyIB5sX82bo4bko/5LGOS1wDnMc
faJ9DXkYgkXm6/1PGD7yF1LCTpPHzUq4UjOWJAZazA+5/MtmG8lUEA3KUvbySs197rWmY0lr+DYX
y5uADTNLWa6rxMtRzh6dDndgm7EWSY1NZilEhFTsTEfyplYmsnAw+EXyu3a8GMOXjbh2G/znCHE4
6OpV2sW05OlI8gr4DgXlt1oaG/WqKBQ/DX1JRs7hyxK2JcXUf2RJintK//U26q1ZsyV89vU1ZSxV
3ziRSAs0w/cQmfjSxxdyK3/tq0INOCscurgMpVDYt3t1nGw+YyEShQqNjq5WKZyImPjDeX5/baFJ
+C8Dt+ZiLtaW49rulLXqVbf/JJBbXsK22oaOSfERcTB173LslFPYQCm/unDBVbdmQim2Ur5TEjUn
tPBPiXsf1vt3uKcXDmheIT2xnKSOFaFYY06AectOQL2rB5fyrs252D1vgJTH+MmXmakIJDHw1JTr
VKWCqDfK/ZVCuwgaAPrBvi2DBrMWjoSreU/uaWUKeOu4eFNPWo46DqGtnFXPKEDxnXD5Zrqzg+fW
IDQyhfQKeRnvdeNNmz2W+23Kc0+SoHyc4WWIGbBEup5GB6q7uMeP5GmKoMk/wjLX4kymXjzwlCsQ
n9pIdOBMkKh7WIG9LH2FyVJM1ZpK5DCC5Y2SelY2hGOGm+9ov5JIRd2Y7E1/3N+nlz1EAf49WHih
FUwK5nEKcYe1+A+GMFB6hrjg+Oq7IziPkj/96Je/XK/j+sGXJ2Cfw2UXTppNBoq3p526ztniJd/+
h0BmmZNAq4O7SMaXQGEOHATtEcPj5Oji8acbsdovV3lwHht55iFNNY98x3KNYS6lXiTLBNvM5uZg
oWTtNfdp5vFetERQCUl+hTaQCutZfWT13eEdmorTq2UEOYpWCCbGWLiqRPOdhylUrS58LKrKBbuq
iA1xF4UJarmICgCcDVBmS7SLGnUJ1MjmarKi/qVetfKPtnFj+Qb5TXnYHOarpJuhQFgJtnFzWIHH
yde48fsP9l6xDRDKQlcAuZk0VYh7Mndp9urP2mMx96buHzuftwjsMj1VrYRgOPl6i6fZbcKeK+b1
G/OoXSK2Kxh3a8cL6nya17Z6FuceaaBU9nmrKnDZzO+9RAAKCipBC+NBR3TNlNxkCGZqUA1ucWyy
R78H20eUlqMO7uk9qkvtgDAnqa3LZnpcrqb63ZjBORsHqktMmQVnfp6OYtuUDuWjc1jN/QXlfhvu
0JWle0SgwbnqWGgpuQv3rXOhHmiLMvbLHzCyTkZIvytlX1XChqE6vy6zIC/zQUQfBRkKNhOUnXxy
sV1jbfm/kXr9dB0JwH05md78rv5vaRqi01rte62/pFV1OetkQQriswhyGb16hplvPPE6kTe7ecG0
I0BV4LWP4iePeASaEshHg3SKQ/HFFDjGWGohAUWGvDN+fTCqoe86KBBWGejyF/YrW7bhISnctxze
G82/GO02uif6FsSjIA2mFnGKuiJRmqbjW+J3Q9T8KkW8m1yg5Tvm/Nhvys5MxEa4+OZsX1nXLYRV
Ab+7CO9GyFk9XYbc3MPjTbA5JsA82LCvPNte4k8Y9yJD7ZT5rQt7r0bOCYBc0sRGgron6sGPRm3t
tmLYvMa9gHZZB1FDakYb60nMMRueAGOaHWORzd1owojB7CZ01u+mjzGcfLRfBXmW/nwjezZ4myKd
m2RNDHB4ReLSTWSH11BWT5X/gaSKfv7kIyPACP/6SsX1QMMFG/kpRo6XMtZ72qyvcGPC0b1l9GMz
EHaOqEJ3zwlDAkMohV7Q/iUbd/4MLS39h/BW64xDkDjgc916l99bdRKXAXOmMAQ03z5vexsoRz3Y
Ms+iLcnYqg72p4i7bEMXdbkvHsHMT5TeE0d1bj71dp8RLiFtaFXnSaJB+3szpLNP9my0hWKYFxgq
NJCitT6ItNxtQ49weG3NlG8v5idK2jU8OaKAmk85DRmvCsWQtltc1noM/RrXwS0RpWCtjdPkpIMQ
EtCW4ZBZa7udo5eHC8BLZspfIkDiaYsMaOjwiXER7GgG86tWu5xjFM0rSIqovGDkkZxjXFJZqkF4
iigMJLbTTZmK2Jl2j4ThGwjiKfdZt9wRR+xGPgAFvpvlJfiNxlEpNMryr+VU3W8yrj/+Y17i1UGX
la4b2fRwZ4TbJ6Y6vlcIW7wUJ2J/QvWZZg/WzLvC/Y9xnBKO064j6lfizZoSfpwSWY8J8Qw05L88
wr3qrV46z8W8XbffOK6c5fWtVfkeIrqSByMBnfd2l2jcnxjTPLPjGOz67s3uJdif+fvfBw0VK5DY
SSehDhavdq1uVP8JGrDh5uO3jWYDB5qMUu65yP+H8E1O3Ckq/dBRxWe5oCLBfiR+m408EwFlhIHR
GX3KjPktLPzlQA9QPoj1WEVYqpWxH+jl90ZV+e7XkGrChvdojbDR/F7o5JIwf23mSDo5TuvSVI1P
CsZajLA8JDYfi91rDo55ZVaz5WPMslcHFJPN/sZZW121eaiAmRIiTmGkuOOKJ2T2sTf2RqJMPOry
mJgfUZMK/Zx/X5yTVS898j09HnSUZYTfLBGXUILpaX/8Dp/mOEMIo2sA34LgBE0jrv55FBw60t40
fLMuZCvMjkgPb606kq+Qsrsk4fwvdvDIgtagaGreNSD5F8NnIxOPQqO2fD5iRmXvIgQNKskCKv5+
Pu9tkP4E1+g0ZJ1dUYFWnZUwk+vjpnwYfBLttotjZCOmaH0iRa4x/otHeLKcwVM5MDtuzdUbesqU
3NWbVgPId29UKFOK3KOffZMN6ZbzFw3caRWLwArbVGICynIAnCdj6GpVZjxwgBWECfeOqBKJHBNL
pOKZQoY2PTe/8af0qjnLGW91Sb3aZC+KPaXayanKkukksZlfzRhk7gGHrjmw8MkU1SB9BFZh6Z+0
Ovbr1FVG4WSB/gPJ8+sdSzRsvKyBaCXZ+bUGsmCfp/pJrK/O1gBm1biv367y0aAeoEc30frO+aJu
vr4LGBUioyhbAixcx/IK7T/3zwx9QyHK53sndp7weRq4kgChuEhk+f6ci6nPcNhmtgu4dyoSvOt+
BNGOTOW5bg8zO3IOqD2AqAXnvPN9URCwZ1UNLnkmNo/C3CIqCfdKRJB5wB32GvV6eVr5S9E5D/TJ
UtB/DEPIGB0dSCTOq9czSnw//JXubIVowjvRQYsPcwxPAnBWgwJBzHFSpX1pmIWoFyierNS9ZRxe
sEo8/sExiouuAhoI+1nCoK8TrTHXVM1iqrupCesy62rrahHu+T0eHoh1TKlX9ww587X9T/WtBIrk
+MtFRwnmcy6CwGmC0X9zKfxlw6dWlj+G4oonTx0L7fNjqONQPbCC5Sol5KwVnKUyRbI6FGy3zSoj
hITBWs0LffxiYkyQiDqoPA9NYF6iFZY2xbB0Dflsnj2Nf7A9vFfqYYS3LL4YkN4F0SSC+LdVPQ7S
7iAwCIQJolvgU5Z3UXquEOHFPGSQw+PqmzH2iSxFxQiTk8kcYg0iZ5NzmKiOXN4sC3l8OefC8jen
LipVSmSXq9/SSvonba/OSYoEQH/Np7swHPfQAKJT+tuXzDSVxBm1SAk3c8zsb4lzHO/oojMovCcQ
x0dE713y3Pt2O8rvl0wzGviFYiiBU4XVlZp6KcuqqyobmDS2xoUe5lXOuJkk+sbk3SWaCQblTZek
aPDbYc5FPJ3cAwF8pNg+Q2vwkWQPrw0PFWmMVMsiAweDN1MtO07jkTssoSlDU683Ol2YBlsdNhsK
ykvsDf3OY60w/I31bvtp0mkt7JHHy0iNCXC1zh3GElbo7ESI58ghgvuBz4jZFrXypAz1mmjm6jaP
qQPYjk1GtA0+tWoENkGPo2e95bzrH2sTGqPHZQH+X/pRQhPjryNwxNCF1ED2yxpRblq6Y7Nyl2ug
QZeQK/+ss6gcw3uW8WzOa8mssqhg1wvgUD1wiXOuODhk1UtdWjp+ANJ57CTz+7Bfi3nHzcV3Nq8M
6Jcws/9Fp9cgDmrKknOEKiQpqecmsfjNwJ9Ka3uUyP/OaVfaok/eyovNIGDGBhz4JlU/gkFSHvaZ
4qWywqBtXeGdln3yhdPGYYWNN1N6CdZ7+7nrdPQ8Kx6NJ6V+cSqI0Az7ds6KRO+alBBPAilwR6sg
vot4VQEQGbzJ0UFdl9kAa58i6Lx4bu2NKSWD6kpEEcxZS1W/ItVnxBT35vNSrHZt64AtRPbfJQMV
AI5NEVCCpF6AmI7HJL7igz//nCKM8BUmOGcSU/ZHtd1qDcsYV0BFKrMGF1fc6MsQ/tVBZrWo/NBk
P/MScMIR4uFBpCpDdziVvGP3vNrmqLK1orKg3T0UxdaK2tL0gpA4On7yG6tC46s22cIfHCCNCURX
u0AbV6SbwUGEahcRLD1Yl3mNsPnYzkCmIVwkvDc2+TqnfQtmu/kaGAmTUGd0CXDY+YCf7vIbCLWj
TKFRaSQ9O4BZmPLDZFJM6v439GiTnLWmS6zX4SzX02CRyI/lDeSMXtHqWQtX4lMS+MEUPQ/i3n+z
Ht9r1TlbyGVyCcC5+5DgQhAbOyEeJd2VdtbzQPxTeL2kYzXRYqvnEry8ePxN7sdtfwSYz7rJrBUA
XEIsU6gBE1LZj+PcZt6fUzAKDWDECF1D3J027rfZhCWqd/JUN3iCFVHfW6pTuSraZ4A2G7fug34x
FwMqR5bgZ6fNirmiAOOuPYTH0lbJ/pRZHZ4DDbwLbrzImzwGulpm2NaOgPvqaqQyxwp2DK2958Ph
aJOGR6y1ZV9O20v9TAafxGA+tdNK+8paFqiGtZ2m+Mu+tRRrHRBipB16ZwXicvCzHtuvHwvmH/Tw
vpg2XCXcxSkd2ZH2rYxmkKbavvWQixh4XiF4L8PfLiI5+qpQ0u7cOExecraj4V4hWOP5ANG1uqyL
rbQzZX1rqiLy6ZI+s8GFTWQUlBDCL7OtlYqhG9DtQnGUKlsSbzQs+cdqdBh1WohfUECO6aAoq7zz
4FlazXHyCpkL2+xrtufvozqFO787aZvroiozThQBCasKa7BSRalVakZtr+lCbot1/UYQzKDQZUcH
RVs2vGA6I2gl4q/Dl5wxw7Mj2bKqC9AZ8Ox631p0o7D7SVSS8OFA+zoX4PRSyv/4XBXPQHBPvzle
DLByOcVDseHXiOX4tOjMJp0w+2u3a/rpgb2RoqSO+pjQH9zCu9oUbUdl5Zc8oUahQ1Opvtc3RQwd
r86eAih4H0TwXbirq4FHcdzgvP5O1zp8Y7D0xUy6IMKbNmRH8U3Xu7si2Md12lI7qiqX6FSgsB1j
NohTbwnGyJtbnhB0kg++d1INCF95bP+/GC8/Xj6TWuuBb//DP+0ytZqQZEeigjwGKzf0lm1DtzZy
NrZfRw/qyQpLPt/uf+4o2rrWe/6FsbYfA1j7rDd6oW7IPzr1QvWzKDYwuKbWc4u0hPkqP408vJdD
LtBUosrZsODu4W6SOuuqSzueeJ9sR1v/AtUiFOXL4PNmiWl7aL1qcY3j1SNL3uvkGKJpnLMYALxM
q/Jza+ombYCDA9CfFOdcwMnd5fw+MSvSKe3G2QxgAsRuNrJhyglMgoF/PTULImKuGa9hlXdSXPWx
bdXQaLsIcQxKg17YdfkwYSYBra2tIWcPLXKIrTLfh7sHSFZ+lsA6WOCxmrO9PhqviRQlaREaB9wN
7NfQwuLqVPJvwfgIHTs/hvnkkuRmt0w1BRYjTLGgOQHN2FfalW0OLVkLZ7bisXnZGM1296i8BrkU
3BJ93Wgkoc5YrP3ofzaDfCZGVdmRaustmWGs/1qoSkQq3Zw8Op9yISxvevwMzLgep6LfrARiFgsv
ogVL7J86gLpL37UMtUyX37KZTAvLVCfbxM1nS845LOACDYTdmyjj0wr50dkaxRQ1hsqT3sIfwXmn
MfAntamzpUSAoydpVwULu4YNLWUpmKcsiwF1frUe5W8t3G6pAqkhf8cT4gP5o6yCgg2Vgj+0ks8p
H174yNp2AAm/QR72um+ZPiiQttJG6L62BRbQ9mAwPHXswTt0ER1xekfxd4eAMcpp+ZTbg77xcdHw
k8ybTgto3dEQSs1LC18VdftogSKi9WfzIup9KxdyyENDk8wkCF6E3WfU+EvfQ9DwwUu9RG1br2wa
UBrk1AXQ4FwbkGrfNa12E8/lF/eXWbCDJfSRqHalVDgqkPuUgQLZm6o/cnj/iHGNLy6xk58v1Sa2
k3a4dHbPT6Vv/IDwWvWGWCjsYEyhAoBwEkynb+I3KEwthFZC5EC/092+YbBffUaFN/o7SgwlfTJG
cqdZ5XV0OrMbLn/QZYj+Fw3KTaAs6T2Yyf4t9JwJIghoog57fD1gKRrC+0DIP+3Q8BbeGC6QhiWv
AtbGGWG5Py2/hbhDe8/Tg3A/Aj7sl4p/rj4NqLVO90TGpcPYxNw8t1JMnyAkJzbPWVi5Tu8TVjn0
7MxVqcHGLZogYH7+F0l6PbjGBgYd0NIxxjWPFILVmOIvyAfqNDAzquWLFkZ2VEZBjZ0VFVhbHYTz
qe8GRRIYLm2rb6kuj0Tfuealr589bKM9BBHTaMcUW4voPCkpTNZKsxHBV5PzQdjnhSI5Q2CyCKjY
lG9vRmreuVYzmB60FmKjL8/Cn7msWj4AicPxV01Qd22QYrEiqMjoHPDsK95AaaSa5hRgUmBkTxfl
yntL8s1SKJSW3fCz9pA7hXB6bxcfU6MO44vQHPbSSPXENFrOGf24hyePA6GYXFns98iBGehJq8Hm
Bic61fDkI4aPfaPsCvCCKRw7aWi3idpPzy6MWqyBwtC2Aik/S8JZXXcoPSHSN6ZiheMNWxv/MPEU
cjjjAgfNlNHOGpJv/Kmyj1dC77hN8/kHBLd1f6FRKDWt2as64/K9hBz/FQvihNka3HwvJfZhg7AY
gVsr22IdaHgkJGftDHG+q77xIzJYDL8H24wzNcMF+b8vADHjUoQaPMKQFfBPHC1mqKH1MGfElo3B
M4URMsSDG28cqKhlxmQqNGMrpKeiIYqQ3rUHIy84ufEOmPafiBwg3Qke+FMzLWjbTL1PfrsiMS0j
wdBHNs/097lG6hYWceCDbMzA2QVcThi6SgVHt8kpRYJbovSVh+JZninGx2e3YNKUiFxSwSmh1DlR
GcOZUcicTiXfm5Mo9OlQUQAZfM/mHI+Yg970RNP4aR/6tnS/XQxgAfWyapxadnQJI7FJzDHqQGxy
Nv9VMOGoNkCf7CBTLZTiD6TJg/WQLkKiO+7jSlPLwMo3bOkccqcwWqrAuLgEaU1UwAvT6BsLEMGH
OGnYKa7EuHNMI/LYjC+j6aDmkp6nJ+nF16q7ZUt8Zin4gD+fDGT3N8raIaIBJmlj0HLk8qVY+ZNo
A4BA8TENl+cmqOWwQPExaNULcvJ6aRAlfjAAyELjQQVhtLM0nqokP9nlsRkyBk5SjMFz3UfZjpRI
08o7uyFh9VoJdwT+BXMh/mYXM2U2WrnISj3xO+prsjRcBlQs8Rxp9q3Obtn1QkGeO/t7eweM5xP9
LPgxvcUkhC4RTsPvN0MG8rvB3m97xQuemo+3D+1Z/9T1jTPUjbsjDPXtGm3DPFXjX78fdUz+Aof3
3eNRp3pH/tWqM6BHS37F/UQ1ynHrKrEjNuV2vBv/TF1eNcPIyW3SEO8cfkLUZWdp+BhXxJ4IA8DB
AwSO7iXWc1PiFCUnjmC8yhCaFnfGANFA/OsejftAfFIJx9f+2r90QaypA6aLyKAb8HmMXNlco6MH
SUOhXRmi1TNJw735DGjHD//BGl98I6DU/oalNk42JWxxaC0pFgsKy6H8+YpL82LQP44S/QK6+sGp
fBDgVHkYcvXiqtVHRkjbBd3lNedt+z0N97k3OLEXO8dA/L3m1InYJsxezKNzhBXCPfPRpIU9Sl27
n1p5WEzyhNsbHdZmuOv/bVRnjWkmDZzb64aUY0iL9ze+XisLwES+5ibxY2zhe57ErR/gGtED8/oR
9Rr0cADnuVzLfqQaJpXLsees6Rbjfb1AGZoY9nKmU4Xz2Vk+gfap1xnpNnggZdFNbwf0fQp2B87m
WeUZZPaGKaJ3Wlffsfftoi3ZSo7S7AMlQdi5FgcR2rbTMz2b68/VfC+UJHt/gphvJmNJTmLVZHQi
dG3M4vpHcOGofuQfDVqO3+D+VZaY1m3eqMHlEwpyd+0iOngdt6SGxP8v14md+Txegp4Ct+u5rTn1
si5UaBKNF09SxdNTqE+Ib0qEVPdQ9kKEbqv323rm9DrQuJqZYCtrV6+4TNvUESaDYgHEilXnQqKu
jgMbx+hFBEjgtu35qj2E5pBoAaJszRtS3Bl2+1ICtwTJaWjkkGAWHoVBlZ/4CQMwSPMIVqNOJ9CY
zHJQhCKFljAReZfeM0TyDClMQ4YCvKB0ZpwuQDDX8+ZLMGdXaTW1d5s8Sv8W4WmW8s5Q1sfS5HmW
/bZELu/ruix6uLvwMFVLWvQuLLcAT0WREBg369VDAG1ZSfF8Cak9bNJ+JdCBn0oLjCdxF+xrTIUs
iyTVvh6QFq8yPQjg3YTdoabih3kKIHbbyJd4Zw7STj1ab+aFqONMY9RD749vMoJvKIFeW9s2hqPH
lWOUdmr7R05+e+pCgzTgxb8YoK+JRXzYuCJXfL4qiisaS2GgLSpfDFLckEN9sjLNqYMDWlfuQMkx
spmBW+VP0VKoKDA9/Aoekx8GQvakwTWn8Q7dGUpcjJBrTtAmPDILw1j30n4bYNHlOrOBJwWVEQNI
ceBpFwMrwltnCt47X2BOdHEBRFMTIjjDgrER9Fo0JR1Z28Zm9vBhIk7FJDoVMOKMFHIEwxeEkN6w
SQk8JivQXkV5nntiX4M6zfJ9XBf9KL4Ju0CUtxVSUiM+BO9rC2lQ89eB+sHFGMiC5bQ2d8HgPEtr
HD66rTNBlii/Czq91y4uFOD1AahtZffTuWKaJ2ldkDw6XXxT1Jy9XSLGeVa6x8UTqyP6ACfgM1sZ
FkjtpYH6Q6tK0E6VxCYiGOa9kAyAWuv/46hQ42Kt33wJ+CaFN6Q/8sS7TGlijkEa3uvbRC+9cP+/
5BNy25RAH271hV6j6g8dduxvgc22+fUpPCJ/MR66uKe/vfkEBDwLdMiT3TtU2Ha2NA/qK4BmXMar
2BGLsHzval5BBu2fa3KIjlT6oG7iX/pDbKmZjMV7+D3ggw8LRrahJunA/aQ186gwpoDulyW2xphv
6ODD3qML1oRt+p9wS0OrixpYH9fbWn2Wp8XVKE+uqMSlzOkZmzp6lPKKFwkBNXGptmZiAOXTS+V7
ZAuoPuESdhzr07NEFxKL/qfN+Xsmju9gH8/S6spI8ZzmT4jYaRyPu9qHzKfNZEFb9bAaQkfjUA4N
41Hn67atxGso/mxY+8jKgrikPhZwKARdHRmdbp1Vat7IvTJN/cCiV27FqWhL0ImyvyjnJOp/8/Ji
1NK5g4yYG8+SjTl4fc8opi1nlBfjXHZ6TqWT9aSBDI2ThR3nyT9lH/TzNc0mewoKRruUaPk+3SF1
HAZPcaSfIu+ixkagXJS0SXwwQGhgRpMNRfmUrjJ3lJTNtUVj5hERw/co6Bk10JgBJuitVH2ClnZq
plIf07h3tu1IHZteUAg5EZdK7d2y2fhOmQ2UO5MsfVHjrsTXycd/yPPxWZ41iZQg3BPK6SczTOBt
IfOQNBrVLWY6mJpdp8U9uxGTIsMfaOvZ16l6C2QQHsdRtKqrUYtlE4Z2zOagEwbVbLf0p2eZe0DP
+ZPo3YG6evNR81p0rD6bXd7dMl27rEcMqWhnYrSg46UsF044Wy3/LSFddjoIz/py7ZYGZC2o5OPz
0FeYdZ39bf6EBiY6FPJ96p5ga4FbOGBK43K1NZbpvauRLbvWcN50vwhzKJDxWaLhu4patt5kC8k7
X/4447pufEamT/pKPs1c3/upTjho6mKCpqH+N6KBhetFWW/p15PC416a53Ll3QHKrtY3Ik+xVR+D
1nT+UIxodZA7vrx0rXu6Hu14Kcy83com9lv5bSreFdTDe8jwJD7WWjTOj9MPS6BW7B4JV5/jvQAV
rGc1/tJURnLh10SpAMkutRRx/CH06KKoVpz3QXwuVTYc48aULaI0Vd63b/b+z9L6WrdoTj37TtVd
jHwlL+eyxulpayYrX0fTmw8JPKrmY9Xx7BZKrjay3id9ngzcKDNUKXSYI4XMGA2CmgmcP7B+tcNr
o1lVhIoENZAfl+CnZtSkQIY74o9HAQ7QGnTrkVnwoISMxuvBk3VET/oO7WLvrBBRrFz+ztzub82Q
lf6pFs4+VblHolm55dAdmHPOWgyKm3qPyJBnBbXDQgK2ccadNj86o1Edim2tzfh1lSbGR2iwM0tp
XVi6J3LS/FuEZU8miT5yca9zzWwIJJO3d/JCB5OfkZakcUUl+Gyh4QFCGmC/jpLq0oam+Fpfj9Gg
h522Ldt44RFQzGZgGlUNpFy4bCwKpPzsebkoQ9Rte3Yz1iISD2+mliHkbQG4XjoRJfIvB8y8hMt9
sgSugJiKn8zVEey7d9Mwyg8GZPjCHdo4GSasXdExfgcLJ/5JiTR6vjEcJbU1Zwn3BE1BbRT1+wSj
6AWzLPR4+sZbmFji6O1XyPklzhEWxyeSmQzAmKopv4Iq2e1kek8vS1OLgj7XtyZGjAWraJFcF2pc
mNXgt2pCe5DeZICebzhdpSd82WUy72XvdGYdq/jaFyIJvSFrrVujTYT14x0S7NxEWJKme+jJTI51
hVh7eIAYGF5EC+OIGs8ZBfjBGJ4Du6+zsOWKCcMkHSTS9TrDGrVZRTfzmnd+ri4gSja5Pm3Btd4Y
AZLMjTsUGNqKaXvefhuR443qYuBesCyaFczdVdXh1eszxaFa1hwfXlxmo1t4y/9E3q8CraQn5eUS
WnEdqK+73z4LxK5JguG55qkzSliUi3joFX2YSirJ4lH8d330uj2YGmLBfNIsVC13rGVAXVWANqYf
1AH0j6zGhhfpHj2CGFmwSOjXyMQsAC8+Ue/WEWS6kBoDLhN2ltLi4N/qiMx/dj1U7cYRk4bPgvDt
P7pTOVH52kV8U60GdiQzG/RkltjeaVQCs7OC6lqp7jjAFucAzjcOMePDzi/wSpPZlJdazaNR672l
XyH/0aXQqB0SRWbsoeJqqtMceoM18DRjWm/d6sr5/S1S5HpNRMFj3EfejGI4v4Ll51IajFDqLoGZ
zoN9r/MS8Sn0+hAlQSbt5GCRgzi/sy34nn4TXsu/iwWBdKazOWb4sWZTlxZKDYlWTo43M8YYI8J5
ul8tY705WqDokEvCYTaq7XhQ1qwTm3Za4P/aYzJw/GgsrdZ3/vytEk9vWxORnkghTY/Q9CoU0GpX
7SMvbYL9hf3BdJxGMa4N135FX7usaD9Ep2Bjb0/AA7GN/EiyIEV2sdXLODB8eZCFlCkSlQGWIo3G
HdRM/nAVepDQUMYBn3SUhguXmEhH1GwGsyT6ic6T/Vr5iHCSBcyQLlVgIdABLBBCE2s+90B7MpZ7
hTUzclglFY0VcD+6KXXvBzPbggC+LWZ54INXkgYJddicXig5WCvEt09dQertIrHxmQgDdEBF5PND
IkryCVRKvfYT1G/SL/ZuwIbvnMzxLij3RPOTp/lO5riQchvymOXxwgrklteIpXAEx2LJBuIoICEJ
Wco+DR1ujaLr86PV2K1qjqj3JsozQqIH9KFw/o1vKgK0rqesS8qO4jOWo1OK5m1lBPjYHM+ctgkU
RdNUjzSynP9hsiN/xXI9AFZ0AGOjxVZInq5AxMmVZ4BdMo5AzCWZCeHAhJYu2nXiwz1mkoQPhC4Q
6jLYIfMrewVOmnKTXqDeovnHqx4Z50w2ginAhGHeLX7dHm877B6WM5UDaYtW/htqQVQEuYSA02CT
dcWW/6evz+LHwdRrpDBq0TX5RH1q6GFuAUraInm6ZOPTgK24HdO3vcJHY+iAPoGhJr9c10PpDYcW
ICQtZjJozhO1gaUOYbT6EEQHSqx1Xjru8yyodjQ1G/z4pfvZjgsd/5c3A53eYHeAdUpcvY3CjJu+
Fj2pAKal44qc0mIHVWUWe1LClMfoHJK84ohiZa93x+Nt8diGCfyud1YWQ8RwOgDaZ20j+B1DMkZS
6QlQ1236w200yZ8wPK99AZddPKnjwvNfmwLCOALrb1rtOraDsZIhXcutHtKeZVY3d0iz1XtgzO5r
BTebVff2+wm0uG2sC4q3Tj04asHzOjYscrGmI99Ito/C248dnUS/gGGx+McvJodBQ7/xb0HLlqiV
B1kxkAxBRPk13775yT4Ur1zeupCvyRbZS3xyqRSMjaH/dT9AJEYEqo3RTP9c/Sw9I8gwrwS9tAaR
BJadNFvIdOv5SEE6DjT+gyS6tU0so0SoBZ0Y1zaOclJENtv2kgGy+A4RpIiww51/7P+hnie1crFA
dF3kevENCPXonMHzjn7aDStc+sXpyo9ECsgfqMLVrN1JfBe2T8x6eLEaIXgq9Ut4nwRIBvC967st
I5vrYub1MUKfpCFaYgM4ACc+VFotF3uX2BGbnDLuwJtHeRPbcRbozMwyC2v1d9IcQWilacQCTJAk
eWvMUADpXW8MfNO4a8azofe+If8p+yl/mtLAb3Sq/dGONb+4gkhD44UAuXhfvqQNZ1qjxpUmqkSS
u+eVt1EWoBMZp00P+6YLUSv4h/40KkiBoRPEkFbfQO/cI/sSvcV+mE69+R6prlW4nXRwJOJ0EMQn
SoRT1vKtDMutMytptQd46cpF3m/tqe6YfqBiJtzLsi8O8EoOo89eX7XeLelGySV1t4lrjjUXJwwg
n5TpSvM8QhE3bR1szXcMuavc6k55ZrnoUgzZS7U/9PcQyxY0Jq0Slbe8FAGp0qYoqUkUVes9i9yM
dv8jYMD9uk3wRBJXS8MLgQboY+kP/zhf4DxOeVZZ+pqortMYGegQzHldKcnVpUxgbpzsS52opb8N
JjZ+iMucWn3qXjeX8KYhcpFzRBZBXrS5F0j825VEzQZg92KFYkselj8/ueUZDKfqsri2jvbeOglc
OP2u+qntjOqSNE/SDvAsT/21aIwCQzVdw180jSDBdTurchEPWi1Kb9V/4JVadLUJKWG6JhHZEQmZ
EvG3I6tXr9uVGLFtE8tN8xDNhRO29BwfJqVxnJIBw48bVhNfm/700LQEf8PRZmsB/N0a8BkGAbwn
O/DYS8A8OiyIs/JdakTEAW2nKpBq+OIi/qCu0SUpLZBsnYr0Mai+DY2zuJ++xH3b820llcyqOs8w
36qxnCBXRDVOrbSKKwd4rVzlafoLZ4ZmrhPRa7pkRTEM45TYHz5eV/dmqc+NRiXpoCrl0ptXUoQm
WPU6mQCj0VzloGp+x2HGPF2mX2MYzyfI3nJgX5VfmY2J2JpBqd9RBNTVFK2EYmNuuiEFqqUXuFws
4InDEX+cQl3PAzTdILrqDPOmJcRUnNH0CyHxdLwWnul6aLOSDxa7nOI5Vb7eALot8me6orXYwKTj
SHkOVzbCeBV9HpjpCpKsCBa39tBvu9EICfhgBkY4cLU9S5nRd8O/Fv3GSL7u92IDlzkb29UazU1m
nvDSNxI2z1m7Y6aISFsjyCzy+gPdVamK8qcLCuba8trsNP4U+DD3pmVO9Wefk44H2ZJf2ZID7/Dr
WT44/3j0rW5NiOdok1D/CmKs8FHWoOp0sUOIkuC4sdHLt3ZSe26cDJLwQB065FHij5zRFq6bad2/
va/yUGT9gCcQJXgt/pB4RIIK/rSyXDAfVzrtxHqCoHtVGqtQ5cMu3AVsEt8MBsR+eTTczaY9HPOA
an5CFvE3MAJ8rUa94AVnbbWiQe5y+mnn3HBUbEDfm3IjS9LQTxW79i104J7FoM7byb5km/UYvDXb
nJs3qhw94c4kbzXQSzj3EJ/P5qDFUi/7fkv8SIVUJQEPWP3SS2vwlUoCj6v3grXJ3nxvusCPn85u
VILyhHJalGxvPTW4rvKyZOre/7tZH+VQ5c5RUEC/KC0z7x+rS3OeqvlzZAWjNLgUcx90SVuA1E6H
nNK5V3nQt+6ZPZGlZMnOTbbQelF+829KWyTukR4jk+wNdL2lffyUXYIU5qMGhrBR8Qa4pWxMkKPp
TGMaxwT/yeeuRWJ/sM8nhydtxZwrQ+DyoS2gP1d7rIV334luOdphl1tD0kcpjprY+nkFZlcuNA5I
8XaI5rki8mRglb4h7CLBIEjxiEAN+3JlfSzD2MPxP9T0SDitsfSx5qVlTUspeXMxzWA6SkCH7rwy
jcprx3PmBzHecj4O+Ec+pcbPX8E3FFQnSr0IzICvJkV3NqvzyAsoIWsJxZieE4DhnKiXsjqwSIaS
419Y50Rb6Jng2vHLuHW5H+TiLAiAzh0cyoTlBCOaIR0Z9I9fR1g+Q6LZWFZDW+2aLCflgKz/TINw
26h7lWBoWSvNlppq9Dm6CQL9Pc5meZS5MctnkFCBWWavF2WP6nCTwhuXiwzMy4pgduZ6HsYXo+GI
CaI70ClKQaO8e7wOfcBpuBWL8+pBPHh4GAssas61xg9UKLbvaAxDao5ltaiQwUjwIJ1mYpYyiwbF
4YB8cw+SYyacsvhHYvo0zDivUphYWZ0vwjc7LI3kUEEYYxp6pni0sA6iUaC/GS8CpwjTa/kJM2CV
0NqSLBa0Bfd2yD3BeLMxJHRWoDsjobRFw0gfmT0danv9k6kbaAEIjxBZHcGzwVfZQHHZ+Fo4FI4Y
JIPudjwtjM62Q+JQo/4IXCf3EScgJW7KJwPMEiAB8u9VXK2XSVImW975OYFQm/CEVuahwMOujt2N
T+Ri0+QoRg2LTQAeyKuV2R4s+d62c70Gq9t+IO+t9I1736e4BVbUxGa+NjTlVo4bNL8lyNKGqAQW
k15AALaTZSIpGqF1ppcLp2jSDLdr0+dfInCfHdfjsYM8Ad53JBib9yFHDKmH9FN9KQ0riRFnieql
72ccH38NGhrfMAnSF5AFZqU5DzIYOqMboHrmzYkv2bzmi2A/w16WHH7GAEg62DPuAOIy0vZswV2N
zvCX7EEsUjN4IpfPCr2zSstASuow0si4PM8X25OMenI5Yz4VaK4NuxrAMN1FwTI69JlJBqCq4QhB
sMItzwL08O10VM6d7aqhRIKgTNOaqMUrck3Y5WSfA1jUTfw8703+s8J35n7x4QwA800ys/w4pXp0
dU/OLuq9guh+nK2Glny1cNVTuKNdD0pqU4OQzlVmlzAg6TQIkUMt+R8N0r6sfeqpDvfebFcpmcYy
bJ70W5EgBsuQrNbPQE6+svesh5cr75f1cH3I/jVC3p5AAsQlQ5VLFuxXgeH9ewM1kxBE3WSPW38L
/ocouOTosAnlDCDE1rthb1+jehTQQwFxPYFn52obrWe+hryqxuZlqa/3sE6VXLBGNa3HUlRSNhQW
Ja+MlmrFV0+rIVeMcOqwyqMtOD62/Dr0IJx47kmOCs2picxHcsaHXxBX2PdKqEB1Pg6g0Cvh1adh
Lp/z6tLbJVNQX9cxkTijtAuvcaZ+akKwn2v4YkbjPdV4FZ6R+PBUAQwORxs6TVNs5aKqXIkzHtzj
UdhSkLo21cZgyDJEKxD8kg1EeY/4OGcfWAsiXQfZWDLscRNbUtfLyCDv7abAwgrDeJ4lB5k3GW8S
3ryqLzGOPoRVyfjdKLXOOI5PnL3AnVeYMAqVsNUqRCea37ybnUSCTI8Oj1p86E/73yTszRmk+Ijk
N7G+g7aS7WmDos+zMyVzqxHRwhT83Z1qS1/QpL22zrgfZALeXVyLcwE1s9Ygc/aEl9I4spPcvm6I
IyQFXusQxQXNulnoyouJ4/TGNR+gIpbDNPDMQQdGUcXzD2HqJRwe1Y2c9U2P1CvGe9SopZa885PQ
qiXYqcn3f3c0a//ETCkRcPkm0NfTip4wPftrQD2KHsf5QqZHqOMnKvS7mO0qAl98Yp6NotNkxoYW
fHvO1Hx4CF29BJPv4s7s2LLFSfXiWx1VKPmcGUkmMjVZJXP3qkKd4byhNg3vAP3KL7mqeMoexE09
lEvBlAsFfZUfe+Y9AwZnwz9TttvCMwBLKNLQEibAExvXA+eJQ7n5qqazHixJIBtDbtXNZPMJKAb8
CIMr2ZSM6R8FUKokGDfj9LvCmLsDM8Gdk3XE8DNInnk+MlPB4GxSCnctHlOtvdBML0pUK3eacGOf
bX2gsPrRGQ9V8L9gjkn1oWGU4I+lKuuzYqkHOFiH6JZ3256J1JtZAcgAImlEy3abThxFLwdy/ZEW
2HUpmhFmh7fKu+v6hGjCOO+2qZXxuwHQow3uMtNrgAqX64S98P4aYdZsJ8muWDSequcqJ1BFL0/0
ZzAZ5UucflwbUZsBJYY6IQYiY1G0jsswuj0/4JWhUtaN31JzCea2uUSHAdrhf3Pho2vBMPE3dUQX
iQpj+UxUxcADBCW7NA2IoCfWsrsybXlXsa5DNb0IkM07Pebrqb4gpqlzxAkCxc/J7aVMY+kt34Vm
5sCi6t8qZLPgZ/inzICja1LY3TlEnKbUImCquT81qVtkgQYysbXOOfH4IpF8wE09n8gqAqtc9JWc
4zsmhSX+W/3LBcGSSm3VcYB9ea+LZA0V3MhJkNQGPwiFAplWA6p+423y0ZxPyhBNN1HMpcrBFsc6
kwZZvAxvveCxwEt1VHGWdQHVcW3j1WVHbLYGmTCkLW6z50s/ykDq3/a+Xx+ukct0gNPKsTwGtiFa
dju/ddMjtHt6f88vl8m4kVN+ewkGvX47vITiu6uLYf4ItxjnfjB5V+9dMa+96680Po/GJTT2xNat
hy0uzM7AXWnwAtE7PeLURnhto8R8S84ECviCMd11VWx5fb2q7oRO6i6tG+kjwziToyCMVGqKDM1s
szQBwChd2lqun07VfTGs7NdUX4ENeCgSc1Hb3ZwSIDRe4DRHc8TQKW+CoYJDMR5C9KThzmdJaCeY
HloOrVLjoN0kmmq7TiX/IsaGqYNw6a0iRN5sf5IVwi5xYutZqjUTRspdOVStJYfi2S6SjTynFWNI
zbCw39S07VFcZiR30xcMEtAF6rw9G3O00H6Cf0EcSMKS4RCy2TUrNK3oL/U7Rm5dY/JQ5wc0ki1i
Jx73urLAcWqfrqQKHQWBQS+tj66RxETYfzAA6mjRvZufdXgrJv9S+jZQX7pOuJRJJwQqAew817hV
g8W4o0RfeS61Ogl25yBPT0OfeUoF73G0YsZmyg2Rr2WgwZScEx/LkQA07Im7a+KT+2rSQgd+Zflu
9K8a/Qug7tXhnDpoq2vOcRsYreIFE6lvzIqfOGb8XpyxdIEp7SWbhpZLGvoifUFsL8kgIeFryPo/
eweRUNGiQDHe4o3OfNgkW/dTDVh1tN2tSuMiPxq67kB+SsWZ//vtS7ktW0sS/TyF/KZaP79Tyvri
lZZN0ajwRbwFngJU15HodaBMSiBtLC7l6r8mI00wbUKGPikMUUzPSb3FgGPl/PerHEJ0aHcLVJ2c
sqdsKBHIPsi496VTFhgnoV4Y2szQYqQTLSoguDSvOGHnhLZyOxtbkM1YA65EaI+/SkBrXaXPxLP/
82hrd9L+KA22tVfDORVn/Ydv3xDN3ZrUu8aWj2KzSjuuEGlhTx/WnDQJ4Rkopd+qcykvOYi6mbUC
6/juT8UjSUQY4Uei+6eXtXO2o2pjZNjezAMgHOvb7GKsBR5BY6YoaGWvLQC1TILtDZGbgpY/W4uJ
pFH3VO8IHO783zbqk5bJGVmBx0h7gRHi6C/Zt1Eh86NdiN3DtabrZg47dboajZVHQ+WqzQvoiYH1
E3b3/FiPiX+hhLr6ROxCiqH2Vw86bH2ChXa5MMa/bsxE+QJVyzlEP4of90IU/Axi9dbndT0HT4Qy
kww6i1CqnidA/HOcRC3FApNgK3Q9+h5Kv1X9XB1oQonpJjsG1W8I7iY4hTMIcbebgADB4s7hdA97
F+fStw7Tve1Nk8CpZGJvFeBxSuALp8vkZmParoreSAKg9g2U6llBFujICRsqkUAlmzhdaU1lY6UN
T6SNECdoIpfzor2lzSGecHoed1xfcX/YrR5kWP4CJeJX/8SJJSbqgX9oJEAc/+J/O9REZQVOQF/F
MTk1hPI/Ip7XVUIfsmpK1q8w1xaHAuzbTKE4JPAhasFB6Fa+FAFng55tfhnq8e9MZpSyDduQS6Wu
Wz5jNyfF2rZrxqjwNt7e/7ZiFI0sb5wB6whzcLca8Zm+je9Mt3ScL5X18pmEZj8Qh9HdkcrG3k4S
/hbxsB4rmzqYBTCxaPiD1DQzHxo7YKmqQFjCO4Z5fr0SmEK58KlOJjL2Yh/dzByYJVge2UrHTjYV
NfabOwy5nH8qo7bmNfdHpdNgQsWDOPD4r8K3Jv4CDmyv2vp5QN3JTUZ6CqrH1mevtdAONhn6ac3D
g1B6p4S9wqpdBsZOa4CtqgyOxYzH5WKBzQv8UC0zMsnf4vXkO8oervp96s6AyRMLHT7oN34+z00Q
hgUek0eQ2aWxC1S34X4SRTetnhhUogbx3djk1Lj+CVdpkZFr2oWVWdUd9aC/WN4nqieL9LPNi5+I
bt+3NdCEVQpNMMEQxB1Bqr3L2k7Ye36NUWwrz4poyRMB7y1dQ0d4dRDbyw4b3q5YiCoWMAvn4tn5
2v8T8a3zzDVkW4bru234URXRjuGjWfxeXP6lfEMB2PpcJ8STBUEYr/lbhtJl6pYbB/u3/awkywGQ
bOwz5uxpQ5RoHD4xApNIxTksW8BPt/tG0L7gkpFMYlvNXGt0TXKMcVlMTQo95PSHAv8+qFT1n2Gm
+c/dD7fHkYJkfBAQeZivBhc98YnCLNHvbMtBNCBVbT2YjDc72AhFlt/OSwz61C0aJq+USKPxXwRU
y0zQBPM4w3kIYBcyRxPr42pPe7xTsLxO6dgYmpIB2knl3jLAKl2m3EknvWFEiR2yD3SC2E7JumCW
rVtg8v9uOkzAdp4x0wBnybcK1AWa+aVdChHRZDNAKqtTuYz9m1kYVYfhfc6rLfwVHMnNn4WYWv0m
opM/fYEHYQ8WSAX0HLEbY4x4Wnm93IoEUqUyzkYe8gfHIgJRRelURjQFry6VWXkwSqnD1k5dVavA
/2tJp6n215yxo8mdfod0UidfS9dBb2PkpC7KTBW2eWjtHI09dyakMnBmivwZGwtTTZe/M0l/a1UN
Q17b5DKoQHnPxW7isyPLzCHrxrTQnjHcroe4xxtA5+8ty0OngyFvZtTQPYIYCMUq7B/y6D8YCxvA
6p0WohQFvuzPkZOHopkoAI5owLAYkyYHw6tZtCGAl3jK1+nIzatvKibVHEeLWNcsMAlDo895yqyG
3/pzGOqRG14Dhmz1Hm1ZqkBtEOIy+g4NezLJXAOQO8f/28vR45RxleHoctRNsFlwiq7I7KpjnYgd
SvJ9icwUZxCFqT6dQJ/A26ZHRBAjviwFtUHuIP5ubqpnem/KaJAeQ6Y9Gh/R8Cslm3LDoUA0K4VP
FtU02axdkyJP9LdoggGHn22prI/lXoSElXBiqzYkymvuj/Xmy7IDbUQVfFPx/Eym/s6Ot7GuCXT3
e6jhqV6AzQ+Qa0GnpHmvCGMaI41MV6o45UDZuEUMetEHAoZGRTdNpDsdIcxFLe1ya+vuusQFamPl
4hHWVzHqc41Dl0CfRWKP1F0cKZxVsfACuoYzhRBQCSKPVDP6QdxBa8w+d0tkyHXE3Ik5oYCE8V/S
KgXqqI0EGFKwF5Vs323J5VkKDjbfX9lWAa1Y97T0IstHL8/WLS8XL4tTp7LoFGOLG8c3OK7wH1f9
hIDFDCmz18+cT/zr2oVTHdj1huTVF02Yd+4PNkIdgRs8zFIfbJWj0QsO47GO+4BTdGHirNum/D/3
0BsSm/kC5cjmeqBW4/w9kinaCd51tA9Gcszx8AXFI4/f5MsiXEycI8VQ9XuNgXv+PyYbA2M1vz2/
czGWw64jez++3VZEeFgVtvu4WMxHjrWhcryBc5twi6CDPp2zsg5BmRJuVNkbAj0tAPOpvj/qa1XX
HnGdzRdWnToyiFdBevPhhfZb95g8VJ3/Q3DipilkJZL9yX6uQ/Bs2V/ee6+DCPXyaf6I0wYzN8b0
fRzcUX/67PkrUDZ0BUw2JikX0X0e0XQWKvvpW7UyuAHN6xWaggeohU9QaGBx5s6wW9uywCwMMz19
wLcJ34J+6C2BBmn2Phzk3c0BSFiazHSU26tVkdJJi/sqYw3X4hHlRz3NvVhjKn6Njx5RgmQb+emV
tbjkdkIB109o4Jf2jUO/Zqe+ZmxC5ML3cg8v/uJpA0UOT8P2dD5cwLuxDn4sxQ5IaTbDUwKEtpJg
G6F8KqxYJkcW3Q7hMWJUFg8YNMBhTCrzMrKZGPQma6GIbm8m6EW3Bx1EgXM7ZzuflmDr/QRoQkPz
EDe/IXJCu9mXoE3jFuufC/PyXXOllDoaQ9LGt56whaqyPs34aoK6yNRjyIOSJGv/RSUPBqZZxdSu
JSP5obFtVjeL0p9b8WQDb7vYiA7gBVkwnjjal/Isv6xF0al43+sbwbEJMVamLQaonqANX5iF4+l+
UzwfQrxgn/Q4vN0bPex2LvXjAwltxmj1/R7CckqG4u9RsRhsLTExPNtmBM4Uepf3JT6AOvUzO8ZH
IKDX6Tbr+N/y90up4Evim5BV+9pCcKp61On8NQzt6Z749s3PGkMnSCHMt1ZoycALESr16Xy2qHZb
ZcEbmaqjydDtDEo4PJe98Yz5+SHjuwpyqzi7YnUs234f9NScpYh1Mp++zMX1KyyxMGlXUqiyCCMr
hm6nKJu0/5ioJtVSwRxL/mUYU8BKwpO2egmIIylcaK2W0np45fDXJOnmrgAz+KylJayPVOrqCHQx
JhWdRs2wxzWVISckwTFBrL8tpc1KgI2wyWXjQDRUxNqMzzzqpiEiPfMDGxQt1N5fxmErYC1KHPMC
HlwofjsylsNjh/Su21WC6M1/BpnuXVXp9+EIW1zsulRDiILHKI44j8oisyxp3HhOXWI1/k5oiLSk
YICuXkEdDuShO77v1pnNtuR6RTvlJvA+giFAhIRZopHTFtjjSqkltr9use4EC2qaK09cVB4YiVjX
SoKj9ccCbqQu4nyt6XsGY8V7mA/y8SvixyNIr2WYqDgeHt8CL5ZuvphNlDOJS41Ha5t21DuuLBMg
d/c+xGLKAQrdW1KXmAJWTCm6HFVKhFLWJas4d9uz0r4iiglGgl3ChgYHDqjAMXGxTsH+lJoLJTRO
xKj080hIAIQ6WoCzhS1AYRMIsj2pwr5lBmrH4FRhCnL6mMUz/1wHuqZGznZW01WgOXEz8A6oCQaN
QnSEhxZdCxOkF4Ya+CDvZyFwr1dX+EYQ5Q/RgesdPuCKVpNVsI7mIx53wu+lsJuTkiB5sYZdsJD2
Z9Tc91WWYitInNliKgKFVMMf8Z7bcH93pfMhb0nYOqfMbhB276z83reVVuCN3gAfZs2yS5cZofnE
f8tvn8eBoJBJK3VEgOQsF/oE4w3MKtFcj2fYvdA52UAyY8MAPOze7UJZ6F0fYpxuqQlA6Yight8I
gvIS/kibBgMiN7rZV4efzLcMtwtoN73ldpGLVQk2amCHKqz64X3Tv6TcpA3TznhZIlpb41kUHKmY
ESwPxGRuMIY4oqerOw9i7ZaYxuyo5T5cSV0x8W+DylUzSWZ4edS3jJmejNcp3esohrM2cXZ+wdvA
UqJNqNUr5gGHMYw+Hmg2qXT9FjumDAo1aliULLqYetVQnAqbY8ngiHN1o/SdbRQNIejQcFGuEteb
4eCgllSkf0I2bUDvYNo2IANA2f1t1N8Lp3yOmVUzYKSuFFHj/gOAtSPYQEBDtZpAapFG32lqitnR
2Om0QKq5SEmQV5tKSdq2NZI//WkVg6uhXVAu7WzfiRhyGBHlzWzWeWn7W0fmGDdJLVTsiWuLzzc6
vC5SYvJIZYEOTE3SGOrtvpPBxZoZLjsIHvIqKv+Q1AFjl1TqcIeEc+K8u51qenWjomLmY/yovSo8
20sgFmYjCIX0fhu4msUjjfkWfqowjKwueLi+mH1W5bSTzHik+4LHl44Tz+s+VszMANAvw7ZY1S4q
szraLNBI8pqlnQJS/XAMnPw8Hk8cIU7C2b/05I6heWY6Fg+HY/TYoKMXF2a1AgQEUMU3EhilOOmR
NFDkAl/0bGnGe8+sgsKfqDMif4oM8BOkyQvN7M1eVHACLIm9mqTA4xb2NVDdQGlmVxrUe+1kTtQw
CYCkdQ+LOGKTtumBoJY9EUBBMwNf55Dn+6kj/ciC/zfw219ln2wzG4ag+6NOncSZQ0Rks9pptSx+
xdMVYG//yHOIX4soJ/V5NARVjgMnfb+etawYcJ2C1nNJ1T9DTHk+yh10DFKRiqBpBNssrheobdtm
GnOuo+XhbdI1eOe7AJhjh3VKOlY6ZVjddPjHl8UL1rT8aftppBbQasNKCNNxW6Tjwrh7WRI2Mv3U
WyqENczfcWlXldMbv9SkwelgJOsXP6eNfq9qEXv5mUkKv5VBddcssKxPzMb2ErUGfuO8BiWXgrh4
yfDwyer4s8c2/wch0jn4aqBRKUXUlVZPUrSEqvHEfxiJy+x5KnYFndXih24svLqgtdPToIN9sGWu
JhOSyKj/GzwURyZ7Cem2ZL24m9yXNQF+ztwRMjRdk74UPFhEWiLHzjl5rZ9L8T3DuzIiJwA84cRt
8SjoXaEVMNt+RmK0A3fpsiuNx096nN6EJyDel2q9Myks5nBacxRGLmRjlD8uXigu+yl0I9BtAshx
I6P6ePONJedGKpAbDe+ufYYGz1AMeXbKG7eTn0IbAbJkRyPOf/RjLXfpyFe4hZlmTp5JOe4cwlwh
SlLK1VtICBYpPxOhy4EG4cAl+AO8OLkwy8KYD+Kp2R96wM4uT+lgDt6V2zK2iKKwwtlVaBsN0VDU
ZkfBaZRkwnsID2BiWbbM6R172smeRGY9/fw+iLbJElIzhdjgI0HRADZJr7aB/3w5HX2PVNZwaPtU
KviMEQW4Fq1fpTGmqDxEaLwfdW89n+GAEB++1LY+xeJAH//2+CvnVSPWamzkXG6BZWHtTwYotkDg
Ia618sFfkECZmWzQIJjwPuahS0WDvO3+rOK0OoRo3g6yitzREMfWxV7CmoRP8NJ8xetA0vypicrF
JSaDvq2NfsvbCB64Nx/HFQdwePurLLH6J3mNpZYlKhWHgrMV1aiOI+mFDEETE9qV3vgOoR40o+KW
6PvTIcnY0BLj8EO1z7T7O+HBZdYLGNpLElqjjx/qRqqKkRzTaquENbT1X+GBBjwaxUu5yAegfHfR
dXwSnLz20roP9DURDLzAa5lYtvmnq7PmCb/aA5g5AMReigXUrC8Zv/D4e+JyE2STo2lKIgyKbvF5
+G9cq8SoYpFuJM4/jc1ViwnquNHC+eYoN34OXFhXJ/Xrnb1J4G01q1+L2P4cV9Z6Q4BylBDo1aTv
Gv80FHHeLLdU4mRcjniB1FMiZGaIQtKzrNvcVape3zfKkKmBV7eaI6YdxvOhb8vY1ufWeZNhwkH0
zd4SYUlF2/MrPXj/08RT7rjYc9hAFADiH6VFnw+1OaMpFAikTT1yZDaYs86BmX7mRPZpHn3k4kpV
rIv8eCSpqoZW+nUZlygnjZKdz7comjzbUSE4wdRVFUIeyARU9S8l9WNxD9S0Hrhlo1Ra2cVmTJeF
bEVIN3XpujYpP4IIVznW0SNnNi8gW91/umjFxUM1AhDPW+9XCwCm8xla7phfY++bbsD3NnJVc/JR
xLytdvNOi3iHhnNxLTl4L+UL0jRj+MDwckKxOgTA5BtqkTCJak3BFbSZhSvKhlaooqfE95+rE0ib
I5wN6n82LhjUF1p1FqA8tr7F+6sCctIBdaC/ie0DQLc473LsjLf7+wp9wjuoxr1e7/ontfPJmYEG
5dJnsfxC8jLUNcezvWudPpYTL6NiWIh2kGuP5uIM1wC60YIFDtU/HUa/pn1eq8FXztHnBlJEgHLy
Opg1sCuhHEBbXnXZasUKS/Yz0mgiEme4u+47ECY+KatLTQ7u0NmU1/TY4QtBzW1cGwVeyu97tVhT
i1HGYK4p/IFLX6Jj4Ibl3C5bX1rAyrlcuOVu2RbIA0IJpHmcri2wil6Jdn/k0FPyQDi2KLbAFw46
oi9r6BeCjEVbRS0RdBIlPqOZg7ZmpYmZRukmw3j/PwskAbApYrLnwtHx0P9EvzrWPshWkUScgCq9
PVrkpfX0sMZttmD9orUeCm5UJo/sVi/0b5f02A3T2Wqou5SChsvn1x2gsP0mD3GRuWRL/Mma8Icx
hjq6b5y8eLqFz2K71FBON29TLrDO7Qx9TITqZSi3bN7PgfeFhniTO6WiRUB3ZGstLVzmvyPhDUnA
HvN9sa/ApO1A/3GWfyMrCgAjSkJnAh9TwifFdLlUmd4kgyS8CbHj8jxEefD2xVgMOtpWKA8NAZAH
BnS3E2IazmYDC9yjpCcnILxHJtE68/s9GVVquIUplstszys+0LYR2PKnVtUfMrDrMeGgfxA3P6LL
9DeZRIKCgz1cnNCyGoRckSPxOYu1svipQD+g5sWFfqYBWbvYSowaxNz3UAUlAFdy/IJi5azn6ODw
mvCEmb9TYSY+toCGAJZeX0BncQHzm+BHsmbIaf6Sk9CubTYXo22KPcvIZqaJ635vuGSCFtu1k0tD
FRtJ68zvlDSFhj3V8gFgMWRa7lYs9+ahBg/4akEe/vuYr4+hH3X6UXjpzNn6RqZpXMNZCyO0w2z5
Bq42D9g7oUNHPphudwO/7PGmIy/dhjacM4zltXWMHjK08sQTIe6+yP67jtU6A2ZTnskyS7Pi5/h/
QrhXPoHRzcHUv5nYmsED8I0fXIxwIdtH1CUvtXVoXYGZoSFJ07ngQoa9PLKRzhJOGGH+NG8yobdA
Im3UzdDTQlMEFB0s4WsI8XTb+9O2CDHrdPK4E7OP6uI2ZfPdnRGYalROu1zYFHMdaVZZzvcfC8pZ
NEsG6urF428y9ux4OqqQY0y5Xo7cn3TFSzScTCIE9TkSWtupW8cxtlK3YX37pTnx090Oq9tLeE1p
qyHSE2M+izgAGV7wXK0ubnmvQ+nGOaoluQOugZ07XufQRuZ1/K1cPXw4CTBztcMcg1+nGNnYooZ5
7H/mgolf36cJOUamZzHFa9H4kukP0jgB0SWqrqbKAj912eCZ6gANMPEC5p0gfaImiVjZEGQ50KDM
9h4R3IPcoWwdk7hB2zx3qxNg7tQapv0yhI2r725KPxYeONxZI9vyt+VNWep/5/e4juEgFuP+WEv1
H6w5ywiOsV2sBuyggesGCuXyjhFiCCR9XP+VHVrGpPVHrQP5SM2172hZ/33AEKmF6cqwwrro+QMx
W6Qvb+5Nr2HZwNRnqx3TZsqcBl6EEBT6BCEpJG2gtPS6y6zFzRDvfPVYng8NAx99neGE2ukulRsA
dkZJAMv0yNgEa7r0cMjTE+lz26G1qbd6EW38DL5Bq4gPDo27Oe0jcOPC8qK7ng76ouz3xmkwEQR6
JLhh6Kk1GN2tHtvhjumpHom7xU/37YVutG0vh2vQ6nlLwkM7DgxDBuIXBsf85ExydSRgpJYuxcvu
hbg7zROhAW3L6/0m+7cadCQ9O53OcWra4f73hnFPoTzrhHNPzgCdzzwTmXxoj4Vr1vKKoJYf9cHr
Wp/1axNhb3HXoG7yP04ZoPTLuF1E1STKNp+t5F6JdWRE4Rw9FurUMUEVumK0I4PhVkctvPl2vvA9
kCossImThq2CqGMjUI1zo2mHcy4/4RB21ZUibPi7nlsHjB7Kgs2XmIqnj3EfVc1dPHh9TMsfsKUg
mnIB46mnnBOg0QuZHQ1MFgO5pSjARBQoSepiA15ab8yCFXRdiZTTrGU9dri3LgEecIjDnAICrpp4
PizES4kA+sz6vnLz5ceEGYBd/FjFgSBtaKYfD9hTfJBU/1RIb1FIJkYRNHRiPO3urwdKbLvMhcJ5
MIBmqJ6YUIfwc0iWvtsM/HJWNQpHDfz+gay3YkPQ8Ms7ZkDm+BJHu8sNe8izquG4vZezg85dMX4C
ui25aT7fOKTgIl+Wj5Roy9pSiX+vI7b3/TG4lE2Hn52oO7E3YlEXTXraXBcW0HkPBYooFWjMGXDH
ZaZ8kg7usccFS9WK9hcydMAbtdqYSmqXQ15RjKM/MK06ABqJVMjfyFPjHgX12qXxQ34DnjXXKnEF
6jXoIKvBb1e2RbEhYqc0kwtXVKUuFlV8WhN43kBmY+nhNFcVnUbVgOeot5oZb3knv6//DfEsTXSz
uSvufcZggOJKBYJrkG1MQTYydfziW3qzI0lFBlxf+Ev7BhaMHNTcHgkBDAGe7Ww0lHkGUtbtQoZT
pISkOqvGO0AIBk6rKNcEPYFJ9Ve3AlHXvoZdHMIVYgJvncLWRopHCE2q5tOs1XFAtQCaJLP6W+gq
4b7T2y1eAEGTWlm3EYy7z8I7b/DENSqteMrfV8FuzmE39UCK3W9iqHrFWrMxqssHV4gsf7Argr1y
NfvXz1MAvoYlh0DtbSBMoCqbyeGGW07Se+D9ucJAbp6wnoBHMkOQ5r8Gg06tFXnWqCht1rid+Zuk
GOBzf55O1oAX23dT47TiiY4jbKacbAdJ9Gx/I05hf1/PnYDezs9brCmIn2VgAReRkmDumIRTzL5O
WaPLylNJ/AZMfGHDQrTT0O7oSuVpcYdLyB1iNVpc/YNNiWmQaFsD38gZyd8ZO8Oqb5yzFCp/6YrO
OLS44UnLhfpOPTluFsTh5kUqV7F4pbPG2VTDmxt6EHASU0r4oQh+NY3SB0sLrRg+nlmn2M6evKeM
HcY5TlxGmZ760rrzHCIIQiB/HeMyaOU8Ba+J9R5JYWS0ocbgnVIv86vusrTM5dElujlIPftY3dho
2FeU5PylsocdAFVqbHJfJAr/vCE8u7G0mPtARp0fVRRgU7LGX+kJ/QIciY12hSl2miz1aHGQxl56
urzf7wtLX1+ZG/UprSXtRJOt48om01k4Si60sSJHt11WVCuJUcAGZtYAFYtIXEOwlrhuXMlfM4et
yMSXePFUPTnCgHLiIQyLpSErj+E8D+F+3s9tnskkDVb2YzRhhVBZipeBU8XhWnwQl1S705cYIfDk
UQ5bKYwQRDLkWCjIvxLq0nwc83RWMMDwmGzU6JK05sd0+spYlCFXgh24AYLkvypVP55nqB/hge3Y
SF+kTX4z4XuQx8+37nySifeOcAIT+QEXfbApIlN/HTem3fp6+xazM31G5SDMRvHebSVOvOtgCzOU
ZjXvCB7jJXfrxl8DZVfiQJFqQHiIMQjK+S1yN7N7lOyJ8b88Tk3vS2T+OLa/pYsbUOyVOf8VoD+r
gXxjQwEpiT22FYaIoK52uQ1WjekVKLPjMQRV4Gkx7A1VhjCAcD+MgHaXRBy98UgmU3aiLsYS4/94
mViymZlRKQR3IvyZ4mAMnSzttl9uUnnfCQAYymL+UIxSpspW6nja3u/XktisgtNEmwgL+J8kDcAg
ZQz9mdGao3iAn/XYnGPyZR52Oqb9hinY8f/SdQkTKgsGbl/BkXpLny0K7b5NcMDs4l8PPtUDysKU
9sY+s8nd2uMjEUamUxlAlxnkwPfNurUxMb8cjaMGsF2my7ApN5+RXnE14KnJ1QW3cY7oj444aP9Z
u/PB/di7I5IHus0tGgLX5GlUJvjmyjjMT3cSJj4J+x9EcsB3LmTfr19WQbU2Wu1KV5HX9jiKifB2
pF//vHzH77Ta/1q3KYIaJT8Wi7/gG2ieunw7bE9k8GmJX/YEAV9obHWXN0u1J32y8IXVZ/BVI9JG
AdQIt6EZQQsVseMG+QCHfWF9rOWre88jkQlwiy6DJLY6bR1wM/vN0G48G7y6z16xFD7j2hinkvQD
YdGAnjVfffv/SUzSqvxQX7xU+tGJ/gEc0YtmASN8ptyxxdwu25YrnM6/Dn8FNhzc/2QW41AflkCs
mtgISzRNQsqnjMBaPfhIyX1+yBkedOT7ECefD6nt/k5BwKbnx1BvtP1dSuY09JSSH3quXvFvhkjJ
HIfT/5fGjDnvFv7y/V34+hFYBynFWHaMeUoTbxSblXAkww8dcr0sMEICg1O/zDph4kXd93yuRAuY
s11Tf7UgaUJwQ57+A4pkCc2T0Zq4/kc9CmHQ5NjRjbp2Z7pvO3yIHfzjPoBhhk+FUET0w7HQHcbS
Qi/Yb6zfuUhNP7f1ZbzOelfL2svlXPY12KTXGeUiepwD5qZPSiuxiOyWYqlN1iT+IQRgzVALYb04
3tD6X8uE+dePWuYsodgKLomjhvhW9wXmQAvv9665mM9tTbNbrPoBX9DJJk+OF0dkskLsWwAn5ubE
AJiZEekUiSsU6FrlbzA1uMpOozEOTV9Ei4Smiovi0B1D04r8eXcYv+HO3+Cgc5SeYG3r2bltLNgp
m5Rc/1nCKuu5YMIXNH49PveSWqdjzDmoiZX7IqMq+2KTS01ekpFwyY7rJa68Fck+j0BJLKl3PhWb
ArEKHuKqLIM9XyAdn4fWzRCdM5vQcVeK+SiIDy5cRm14N1z0e2uGnt8T1BXap9NfnzRLP9fU/KXJ
nB8bA98WHqXSx48K5CwdJQXDzwqRnrorVGwX25knN4GTfs8do62nQBmFYXuxcLA+3/3JHunbe+5V
9qam/wBggHhJKzUY894BuM076MGnmD1IO3NjHRX8AayKacNZ6m2wCac11YznaD/8Oyu3GH2gpvoX
/JCVbXU5IFQg1wJ0BHi+VY/QZYf/aBIPwHza56KKBsVgOM8hRDTk2ZzZTm98IofQEizCZBz4tHR6
e3NsIy/Gl9gukwRkNSHmXkEsFUvgIe9OCTyhG9h077NuFVTq9Krfb3NubTQtEGryMsC5eHTuI5Qd
SeFrUDZdkdi90SQ+7UoTcyPrdiXz2j+5zgltPTKV0ZNItS/gy6KiJIBaMlpbHveyTIb0uz3HW2fs
YvAQqOlMD/5iRDMProeDcSXfxb9ktDqgebzXU+dbIb/l928tn9pAQpzpDFLBHPQlU2LOLj/kZ8za
JHJZmkTc4Owylepjzry/VyxkTAGRPR9QvxHR6vJQM4xQAMNs6U49nHP9adzPNssOYB9zZwGcda2D
uGhT56xbj+H1TBtv7pe1R8U6PGzODG88ieQpznPI8jB1oESMSeMY4/asbdJsmhDfOxKVv8Dku1hE
ywT4MUzH+EbybRWL4uF1r31GDbQ2GeI2UvC/pm8tfWAbNtGj/hhVkXQxS5ZdU400rmV1UC3Me+vp
0uquSTuceuJALdyy4/d4gFCdBA+/4z0/ZiBPfKOs21X12IDXE6ukWBVy/DmFdnY9HEl7YFW8hnIr
YdWVYYuxaINMYvtjCXwnL/eQ9YhUEVjMCMms4pefpftdYqBWZ8AqSKnrgEs4JJ6y7EWcf7wkxaHr
bdDosnyetHx40orzbLukEKpV9eVXyuCNqzO834r3Jkgo/8khS+doYZ8whLb5aZHxF9ONWiFBq4Xa
/QLH0X9zQxLPHoDeVo+veIfIz6KduweQ08aqvVBBtKQPQaI/KgxfvwhoR50k8BW881s+cXESRFBl
SLMug5r5GqrhM01zrxyShQ+Zys07K18whJw1Pv0fwjvSyY1H0EAQ5gEYLKcN7ja9fjM8KYeGISGs
pLm5ItAtENfMGjLXkq49JaZnJ/WBGw0tq0NV7a12O+OsX5QMH8QCyIqpaVImhNaVAIpYBbuIjgPH
aPbyTPAlBJIS0SITwWta+vkcS0B/LojQyMhLj2m/UYREXy1qgNo4naIEkHH0+hxbd1V3jOpSN7LJ
OT3FklUzdSaHqSsJw2jN2pcMiEiDZAqSbFWMvGv4Pp7nhv5GDq8qke6Z4ONUXttkHXNrd/VbTDNj
zQ88/A4fxs3s5aHfw3plfYrBZQ5mw3xF9vH49JEiXhFc5Bq1Nx+siHBahYkmofgSp7J6RHmywe0q
Fd7TYqzVQW5NPHcd3D8UYEdwAcgAf2pB81smyBVEvuTY1bltF9qk6aMfA/i4UHrQIEsS5RGk1BJi
8/Om61aCrij8GGEsyHbo0vqPijsWgFIP3INywtDWd4JIElA/VgUi7q6E+kn9ed8hACX8+jL5d0au
2Opd1jwZMu7+GdcaLXmp57T8u+7U66unNDdOPMOhX9uAmGqRTJsCwnUvegLwmC2/Bwa77nSoHpCN
A787/19xJNwP4DwS1yNA/ns6GQbm2mzdPed/DpwLj4xkfGuCk0xPMbD7H5XuZViAWB3FqDtcFDGY
sgEv3VMdTlPSQ4bpUV503Fc3MaS7szlC5fi1xnYNpDQwo3WSqmzqfxfEFutsKNe20l/riyVuSbEK
W0W+H8aEAKXfCDvhnsIszGOWLSPMCLWUB4yKwYtJ/tccyWiuf6b1zNBZwOpFvgFjJkM0kUYIGb4/
YE8N224h5RB/OQ7xQK8hBm/eG5K6SiHmTiVEo75tgcvfXQ/ReLxlVBtH1OeePve0uhtzbdvowRO+
V/erU7+s5m9z4QSdWkAcHeTNtZImmSVfGaXw9RsXO83wx1eWDdAreMFIZk/82Y17VdsjbEs/0NF8
ZTrlJAKtbNbEB6pfH6seRS9qFqV3H1p6liG8Ek1zT3wseJpECsgxgowtncEXOXf3RhZN6ouUvYQg
VRf0fIkVRHCSf8YBHjmND1kHJRJz7SxKNNKsKsJM4G42zAFaqIaS3BfoGm4guMUyPKWV+MKRF4rg
AUGtCh88HchWCUz88wE8Ur1Rqz18TzCABhQ4FnNTg85pclYxonQ1K8ceBdGbaoRIgKNSHejQ3TyF
tZPQiCHPEkdAQmxYFxxVheaLU2K0yX2Ds7cz9bgflcW7P5vKwl4OplGJz9pFj82yVPIBYGmDpcGO
Nqsbjm0UGd8xsZ2hbisBW4eDZc2jLRKiEwBZ67jx1yrvrrpL/Y5HFjgcb1Tom64H71H7BCK/vkPp
/fqtCXoVAMzjzu2Fx7uMWw6AM7FE7GPCMsxKiifIBF1g/5GK+ghFgPCAgpgAZhebQ68z7BKtuK9A
8g7KfEbHIe30bXrDadnC84CWotqb5WXK8O1xhWkC7zr7mFVHZOBhbN8jIWnNTMCNuCctPJDa09h9
qN90EHvUSwvIbtZ/1wxtrH2zKMltrdFfafbaJrrvuaJLgg5Mpnpruxe+oEBKe0nqbseoYUsQrh4c
52R+1FoOpfZIRXHcFL1SJqYHMN1kXEhortj7kXA4fDerFv0uW3pgvDQk4HcZerg5EyrH0Yb2Sa/7
PpfJO1zKecsdiWkH26OWymZ4N/rY4FIu8XCxrHYINSqCw9uy+59WVkKRMRxmhkYqhggtmBpkRidE
Q7rDd3raEY/5V5HYfV4q61Xnl+81jPowyhTFfovoxiUGHtGDNNus+ANY7rv0+Tg2krFfc+rKdoF3
+bEnd6mHMRs5AtWjrFVMVM9BXUnlZvi2ON8BOWRqJrfoA90tej5HHbHKAPNBQndmTKVqtO2wpNwv
kKBqiN/Kizpa44GQeExujuZLU7/rgzmX1Pzu0z7Iz5cbuKxbMHR0f9vFGXutZGA5bB2t/RBNe+lk
94lsfjYnkijgvQGLHYnZ5C4Lavhr47vOiHh2HwyZZj8Snq8Q35CYLuASKuZMJ+zL05Av3NX9gcOG
3+M3FAhrptViZmagn7GSeqNz5RvpfpzeUr7Mq2SPb7y0XnJwL7S9DZOcGqF5z5VMbM5BQAg+2aSL
C2We2GGFlqCxLnhJnp9eOxu83Ptcu5EBWOXvbqGBzPJBOPN4l1VV54tC/ZT/oYwgCwdMoOC7nFVn
rMNILnwULpnnbgSZ2bSY/jGG4TSzX4uNm1SeMnvaH08+qlleyRXjdeckPr0VJFYzKesCpKHokuWp
V7Ruws8uHupll2LTC6ghCdiCAK5xTjQ9CAXO09KCT1y4tHdPdq+8GNLdkidzB8sL5f6xOkptZ76F
Q0Hbh9UsXaVIhvUvnyi4pJfVulxZ7NOCy2IgaBNurLaxSXgI3aYJrIq9gSb1viVsFqpvXF1i0qMc
kbE99isJxRK1m3a8hg4wDq9AJVogHoBduuqxnoUwTUB0YSaPLeEhIi9/XAliwrJ5WMHVJNNZCq2D
L/eZ3iq9T18ochIEx0F3VidzX5HFHT4cdpFdMS0B/PYtqJqm734N9qmE/ZxwfQFw8FuEzou9grM6
WvkaYfoFzwTYsn13r+dof5iWfrjzBnOp78rZzmze7UXWk203nkP2OhtR7ucPmmVKW795S8rw3w4w
+mJKz2ILciEte0SAYz5pJsm9lHjI9dsHNDwLqujs/d7lS42KBDndSjYVtLbta/j2835Gpd/j0pZN
ajoJ5m/srbBtcZEOGFKW/nfcBzpZiVj2HTgUzgNfbGjYd0kl+J1sPWtzlKsYyOkJdq1yemTgejec
VBKWcEexfSX1EgoQsNZ+IhvhI2y3ilcAeKzFGkkVfELvIkcq0VSNe0KfSkPnGGHmJq9BjVnkoLNt
7p2PYroDkWY0qdmkobWcvMUCNU4vDIaor4uVnDfqDdkGA28RTAj3FlFX6pHdxueaiEbcnVorKIG1
NyTDdAN3zwVot5qxojlwCCAjsMm+srO0tXvTfCL67U9pU2pGT6h1+wS4AxO5t0wSwYO7PD6+N8hU
jHvfMkdkLsXpRG7EDX/0wKD4Oo0bHQfjtIyAizlWJFQi3mW0VJzHeHvn72g1S4o+MdQUBNQKT+qM
si1mV06iqVYXB17U9hb5P6j20PGr7vSj+FX0LjUpej54X8ag0KCfXRoVWrwyOk42geZfy/96u3y8
yTNP3MYAfQ+vqB5QllACLJ9ASxEzaaqWTYUQdBa9H5NcHRcasZW9VZHFlJ7bM3ZvpoEosh80RxGZ
WOKcdsGPR5WtOtmsRm70xhCOHXMOJvqOSB17BBRyzsUt7tasEWhlcPjJ4GuQ6Vq8sVvpDH6z8npW
qMlSiWGmKYIV3bL0Z+NXM0KN6xY0ZQsbO3FkgQRruJLRXHp8o+G2V2gUBfvWnThNcqB3/AH/YiIW
evosYhW6i9w9En6zhy/4/GaxzQHh9eVxKUF08gk8SaLhe683UigyKf8aXeMQHdWEtCvjrARhuCAI
f4ERQrBfaW1/0ES7GwZtqv/oMvCvNDS8k+sDMFCs0jUAP9J63L2rstewu/BIO8Y0NI8fJq1iI1Iz
LW4fVIXpFTBdZ+UMpphV4Z0zvh/R6fameT3A551L9kgmV8mG5WeN8KgMO1TGVoneyguip0SsXjuU
2xS0yQ2hLOFDKkvMqkS36JRgEBwlVMkRX2CUbUQnDbDuw+dTT1lv5goNkebHYmTby2fR76vp+/Eu
3RBF2FPK0Zzr8EeQt3plD08pYlEdJ+MSyE9mr42iqSO5yB6MjkuMU6GqQzRIaI8V47iTtoyhEMTf
4+tKrpNftCdmPbOBsmghNSqBYjoFHeTw1fBIwZpFZkYT3Z36GieLeuwPIEtmEzyWvdHecE3GVZki
KF6/Na7UxxI/ZVFwXQ5103z6Eoj1xsZyWoTLCCpRvz86J/G15vskkBMRvUuc9w0wO7KcmXHRg1Ur
3TWVfGZFqlocti+zbLfGAv6/B/NhYpuQuptKRvHXUEtzaCuxLv6KszZZrhFkxrK5KAK0WTSChuhu
JZVE5XTPYUx0gFRICrM8J6enXXT3DdQszQHHRs5hkp2AxR8z5SKhZ0s+yafvnpXibmKR4bkqO416
BFdH0IzQ+LdeFIeErrKmQjaB9TGj3M5BEQiw4y2Mucz6b9Di1b6ztHUbsgyrvslEVGtxcuuGyyDJ
ICD4om9SAptt2XX4mOajKQqkT8H4ep161jNmsahKC8uhIMldi2zFktoBDzfJRVp02E/FcBfs9umq
EQ/xk35A8juiHdCLehkrRV0mJ0NrSLQhyq6uuDl3MI4LNmHbnc6zcL/lK7hztFuHChU4yhQ2ZylM
x8X2p+hyftKaELomDnWE5GcORZI0AKGesLLcstVmgzsRXxHf5ma+XetsBJrZuV97QOHXIvwGsnnv
Kh2IaoxYPoNPx03TUIAQsbfBZXqmqN1+6PfMVV7bwR6bCG4Nl5z2Gp0vDVRGa5rJVh5LNx51ddE4
5/Ay4G6lNeVJctVllyl7fFGnlE5XfICqT7UrizghhL1WP3BOGX3ri/buQLBY5liGZvZjEX4T3eTq
T5zoUwtbGDKmzH3x7vH3vzXQRztX8uqxs1hah0jXQ7kBvyzAc0+078OAX4Zupr6vH9woozDrlIvM
Cts2LBg+2rVp7tJrX+xF0AL3ATy7uv+jZsNL5jkK6hAgptPZ5VcCwmPJisqdGxS20JPVH0DPQOPS
c7UNLE5+yfTmKKwdHuzMn3ESYK5ff9Sz7DOziTBYsmdKNURkcWrOOr4lQ7GgKHpCQzLcy6BSMuvn
+Y/Be2HzWb/atngHOAyW4SsanyVIC/gdktKyloZVgy5i2Amuw41E8joxRelgO30s9ZhoPFkKpT6E
Gd4TTFv66g8QhC2iNIP4Ng0LKvbiQ6AM6Gh8vrpTgNy3UeREKQKOLaZrZefqjyZE53v95zj7x5qQ
AyZq9ab8mMS5fGh+Oozgdo2HRQJ2j4zN5T2XvkFRO266Lmz3v1najExz0u6SkQPGlelyO+mnxHnx
ggrzUYdzFwn2vuAWruysVP+IWQg8XT497ktBIgrpAnmC8QReGWjlywFhbnkVnNdBEIZOnrUgFffw
++dgmytHZs/fMDPlskYnlrs32BeZ7R6gjSkKS+c/kC6rHAjP+n4sKkXyFec6CCYI/KMV62yaNfoC
+lyHNCq5IILCu8CDUJ8JTsocoAxiJjLUw+BVonoCuk8bCfoVScJHgwkkxcmFjpRKEgSvluWWnVdW
WAP5Nr0seKOYPpaUfprgR3atKRrFMvLpRfulJalTct60LLH8MRI+Fa+AKUpZeM3OY5NLxZnPDD4A
eZJgcO7GZ/enYSULE0HERiKUEW14n3fqciwMU7Vxdh16GyD7lGLjiM8yWDUUiIxlHzP3OmG0r48R
KFnSqyudTpF4XVmNq6NQbWqPXIXZ8YhDtGxxqZlI6KMvvbA0Vp1tq3Lq0hc5KU5LHL5s4InzmOhk
grP1camR+Lz8RAGjQ5zBK+x5PZXbO4vJJfpd6mrI5LMpo4KZkqqJ47gg95YUN5nLDY7Bypsa1E6Y
zcIAYJXBWpUT+03O29fmwLn4LEophZIJHq0JlzukrKh4MRyoeZgZadwk0/z1W91M7euAsfsb9coB
8B+1olhVlSqwxJhlPZpdjsI6e1yq33QbPxHpKoePSjm8rSOTPWBe8ou0aAH2tbRJ1Sst2oezrJ5S
s5MWp24/ckm3JT+MM5Yy1TQSpMPhok3WgXJJNKiqcOgYyVkGUE1tuqwV8JHGmRfvIBed/QDeIhLj
Jl/HHWDP5qLqcYA5sK+L00gAKH9CfME4IMAk27wnU9bLsQx4m/RWveSQXlDXCCUvmeiMGmAFmV8T
YmX3Duh0Aakk6Lm3tFsVn9inDgrQSOdiHUrdNZx7gvn6UL/8fwc9QjJSqJPWar+jabJOXPLyD/8F
zoaTokNscVXYL2v/IXx2p6c7blsyX+V27VGKO6XYwulb8R7t2kxt51ftRfp9Oo+g4bJ+qqZQRd0n
vcYJ+ncIFjAnSxPJT9L0MS9vVikKbQwytYqrGRtaHkgUee1nXL69HzdpfiPuZFwbfOvNdr6/Wgh7
44ZRxMF5zK8UKIOa+0/6dPKz2lB3oCj0ylZMttT8YAQOkJ/D/8viy9+tpqmzLKn0REFiiS61YiCQ
9r+yFOSpLQqxSu1j0ykboOmYkvNNFuOoMbzpoLIJUr+4AImXcCRq3zv4nhgisv/3o3SYPN3ZceHX
MYoOvi80c35j9mC54BAX6IrjPUQH+T0gXwCB8+53agRSr0mXhIJO0b5fQ5nupJxBKfNAR9nXweRu
if/CLnfwTB4Y0nstf7XDO8bmjU2AqkW3sd+EoTJ9dOMOqkH6HwJs31KfwUgCx5Z01Pc0jsCDD+2T
CsooYtyrEiecIDHprwT8a5kkcR89+yFzrE4PTYqlVlLExr012zd+8CJkh7F4DU0W9HQuRhDQ+TOK
YmeZ8owcNXk3aLTefkowkO3QvyrKfpJubQo3q0MT6BO5+lRC+vtH6zUoO+LKS7Xd8os0fJsb2rtZ
Kq0DaO+b0NLlU2K3K4A1Np25UOnWg9BlxacG3WXJt7Rh6oY3KwRlMJ3Wstgk6NNFlPYYEPG4HCzc
LZnn0OSQNu2DVNpZPJaWgKGqFM1gGzpBToE1QUPqc6zJ9RwQxupErsEkJjiwLbl9a5j8ndBtR2A5
Sfkg8jpFoxPA6kIr2SvmD++f+/DxNHH8oZt0psH5ASrVjH7cg+eN8vlbYHTC8xMjyen8D0IAzwUM
Sy1Z8lrRLxtGLWSWa0fIafIID9apsKXZ9cKTgI05gbTimpNwzkUGt4QqbBB2BsIFAnz2xfjD6yRR
Jum/F538+bNRg8WGDCKfkGJuBELEzwMzuFksys5vHvHJyLa8UUdXRm7MMWbyxxo9NDF2aCikpshr
ni/5WUNKVX77/hUe+aeQSwKs/uh/WzBcgeW/KBmVMAhNO/S5vb36LBv6LCuXvp8+SpE6jbFUNEE5
t4rx8TGslh5Z168YmBOj6qeu6x6F3tQP+bq7Vw54fEzGE4+3PJ9fDHS9Jg1Yr75Dll7gIsVNmAq6
KAOmj0TOVBhKS6lzd+PNRDdGoZ26siv3rIcB4UwOBgf7Z9RBtDrUOLtGaC6CgYeYg4AGt3iYW3dJ
lkJd4sEJ2icyoHvawomKJQOA4k1N2de6CJOxxU3Aq6Q8zwE57cD+LOHKK9du3dimRP/JlhTsbwmd
2c9iTMqVmASsxSuk4T8qg//SxL6WOXTEvxiOfuGQe73FByQwW8AAEAdZ5GRUVHXDBZ9qTJ5DwgTR
amM+Vwu2ORizZfXsYtNfGwlrEWnKbQUWs3jmZjWwgMYZUkZnRxHG3bUFtzV40YWLZzKBWD3FAHKo
/WvtWhHryC1Y2WnxAXHuwwpf1IgnL9Eyqqkvw/JD/Hex5bz8AhPXFWU/91k5GHs/DRKW2QhTuuog
09aAPT5uZ4JfClMwu+xWwIjLyYNEStSlT1DBAsZKhtLqhsOIe5bXzhSbywcjlZgpqiwrnAtY/qZi
PS9BxaoCwy8lThFQVFTtFpQovH8xoHM1JcA1mwrGlFEYNXwV+InocN2xQnQh3NTjp0OUUGNwAyL9
WDGWm0D3c+Qv79+Ih7bvdSnA5aiqvf5Gqd8OarPI6PRJ12JYmDwaJGb0tD0/cNjsJCEDUCxNuJC1
BkCSErWTlhjm0dc3Q3sK0G4r8pQ/Tj+WACUsjTw+kSHaOtunD6KWRhqy5adLbKKGKH/BakbPYcpZ
RTFDXA60VatZlLNreIPpNqJZUh6wtn3IcjkSyeFhmZRXyx5jojkvrz1xBKz5j9iEZKc0atEyRijC
IuoENVPjuEPzDSHVNL3QxZjEH5cFdwPkdhthJterGtmO6H6j3be3Ls4UTxbESlZYkBI4dZDw4Gi+
QwKsc8+tGESX+qnHTnXil9VWeF0uUFtyUSy1uQmwiyeIi8rr8eZCZQDAOeXfKzdNH5ldFLlzuL0k
WMf+FR1npVizgca3YSx2sMZdg7rA9G+sJzwC2ncy9Yy3Fp0Lu7xruAPTPt9ot+m25f2EZdptngZH
L9ke/hn4NLi+DblQ/3vZ67Q2cmPJJ8kHDHmIRG4vM0u49LY3HcBRv0TpzephQsEQPUJodJOS+/u6
/uSxxPKL7a5AhtM7SiSjxIVkNLQe2auKTC+tYxEgXPvG03nOckj7Xi6/JvbqQ85TaKKQlM8rOSbD
KWK2Y98WRe70RmMWXA3smpFs5Xqlf+baxD4pkaUqQNRmC+A09Z2OkHoJU0bVIJHGirMOnsr1AAjs
N/p4cIoLUj+LRUsmtGInxDWj97BRDbdDXCqCq1c42hrdSWh00s8Sqw4Kk3vec2qgXOTGJi2U/9sU
KTligpH3Jg/PYU5t7SZ8ncHYeCsTY05LaOTrx+fb1Wfi9gFKUZqPQvuvjbY7A/KIPC0NBf9RzRdv
gvCNp7VK7Qh8ReAue2qBruiuJfboFMsp+O3Twt9OQyeST8GuWRFXQ1JoFMyH6mG+fpNItEYmJBBu
wAg85c5bvZEeXzK8BiUOZUxaLZvMOW/sPxiJ3sNLT1wj42jVAQo1R/6mkZGEnTAoCyF2RnZV1UA6
qC8hrxqEX5Uyfh3cP1/1vWtUX7Zgewzed2UfKAsLJrV421uX7uSMxP1l+GD++m0WYlrpcAptMCTz
pZ5vstHFrZ1GGKLwtEhVq18DVsXDnbWOl0ivcgganMmNmZUeZgvMtNLbNGPs7deG3m580l7UxIjg
r2f2VH78Rz3qrAPBZB6K3nTp6Za1QemMemXqQGwbHuuKrV5gTl5K9sc53fOgjHlgh9z3kQgQqIiT
35QoupD5HMWF3oz8UbMq334Covavv0SBQzDP00YakvG01fAnCp0QV8Iw/YUkhO+stFBThCGV3MDj
1tSazQ3QpdZRdShPF/L9/1oA/c6G3RmAlB9S//2BS6ng/liecXT98y4WqY4KWd+lTvKjvGfvWUzg
iBij1yyyqAHHUBwL1dbHfxjI4jOBMKZbp+isjG5Y2i0Hxba8XVO3/KeirtVLrvzB1qYSrs1+Pm5J
lEPUeac6tLoG2Mxv+c7tu9O+lVp7d9RJ5cJ3U/ym1oLlVd2c97O4e/pnbaMC9c7Ui1R8Ow9/atky
vIh+nt7cJQqoQ0MXVcRdH4yVjawaKvNJfanBsQ5sKyCE3UYO8iGo1ZWPf7wKLHXt6aubkS97CYjn
eAUKpYvVc6+xkg4K7ESMRbdWFEcAIIogJb54kiJJl8tb6y2RtkB2Lxv/XJHi61RPI7S5hBeo6SAL
W+PNmVWk4rCgJuzTkyB2ufD5XRRXrY7NzjARAW9dU9stPQhUFaRLTG3LDgrjACCan6sbZMdqNg4/
cc6DXZYsOZJ5XldOT3P/tm5WTe0CnjSHqEWFq/xWfzUEeVz2cK/oESqdwiV0uT0xlXIfpJIGVuxp
jW/xttlX0YPbBiP++z9hOgLffGBel3KNJkM5mtCZHe43a4aIK4IMnb+aZpoaUm6s5iZVfCIVVvTn
e5pPKDDRs9VmcTwld5VSMghZ0TchwzA/smXsnZunkZh99Vwzlnk5tSOJflnn34uR2oNfSt1UP6g5
TVy2/EAFqgQi+JSQr2loPHnuWRQjc7g8uK54vwCFas6JJMkORiM2NzNF6a/aHd1llwVvta8pcR4q
S9lsZJaV0RXTYbdV9xxO4OAAajy1zuGGpudZa8yEl07FgO/uOpWS0ENTAssmUxwm6C+mJENkoFOM
nJq7WWaUVL8M8l5hVPm96ufjO6Lkynx4h/l5cPfOMJ3MiK/s3uutqMnvlB+jnVxXp52NskGGUF/Q
AGXYwuEg6NQk+NP2d4vqFOy28L0SEqSFtRTD3HATACBSPSO6mt1/gaFvV0L4TUcJ6eqlQOyOkci4
Grm1brKN4zXOGhImr/pDPL8lyyAoUG7D7tEs+zMgbzUxULMg5J6/D+Hohszz3la1QNW1lp3U4n7R
mILgQjaEaGi4VVd/pGfLy+sGs3OrV1deRRie1qq2fNxlKaLLJP3NYexHJESANnqnZWMWqVEXwF4i
8JyQnoBOQgGiQT3dby13mcksrKG2FWNtc2HsyOVCs2COHq0oaHMKNkFcMkZ/TdPbYMV8KNB1CrZJ
Gq4m7jS4FXnWJ49NY5Ce+FUFXfS7Lmdpxtpr4oIEWR90sI7P+dgY9pmW+1ytuweyFpf1AA1SSHLi
dBu5qTr9pxRgAwM5jXni4YnfDYtjO05OaHu9y10liSug1dc13daE2kF6v9074J+NFeK3XxNJfGQH
haKWksdrLv1amBIsrUaLjyBbkYO2MPlMMFdGpvIuqWSoBAb+Sw8SOPPeRiRzq183c0TW2K0fRV77
mZVRqMujB7hqBORo4m6Rt43KB8eiKFE7GI7AuJqgbA98jlTH/9nr1JF8oOvk1tBafTeOY/t4a7do
VvjK13qT71FXPL/WmNSPNJgMKlwVa3XztXWVJ6i6u3n2jT0+DWoS5tf9lTFln6gbQnCGyFiLYEAj
EEe5CESlkqLx3y4IdLe7C3L40+K7es87gsx4m8oCg+0KNGZsQair6Y51bj3w7CdeyjmEglnBvS4H
oKqyBzKkogFcDZHGksQiEPK3SbLpGW3ur+EAb2IzJzs2nS61vfxYf8F4MpYM8w1Va51J9RNFCxou
paH88lURV7QFROah15zUwGDzqRigUEQ5Mkjal3iFPg6sTY3qYG63YO0hEvaH3r14r09Ss3bGJ1bv
WOt6g41RIJSdgwP8/eM2Hy7DLkPZ+MzlgQwcKGYQHhqKLvdZDe533s2EUhr/ED8SgdizRiLEIdjz
E1mtyjM2FhZRfrMgJfoO9txqT/hc0x0fBh0/es0w0jcl4Gqv2yLBjjuWBass6DLGC9OC+YWDoSCt
j9KqX3zh9xgvTF5IMwwreVOUvsCi0lHT2sWSTYc8/YAcs0GGbaZcnw93eHeMGXYZi9rJLFi46XK7
hDJ0xZmR2wwdjyiS1cpcfYBjmo9Ke8BIjQ/wXOr+HNKsXHQRelas+Q1L/WaYvCN+VUpK9al27smh
PFHws4f9gYtLRb76u6I1YT0z513FSnpzP8jdQnU4OctxCCRrFK1XjmWWOTCdcOk4qxuDJFQdXEKL
YU6LL+FqEofhEmRzw6uZLRfLjNB7/yWRhpAcelCbqZHU5YZpxmvGjAHT1/DFw24dOBrLN33wrDYS
unG2f1FzrL7yU5tbK+81Hhc61SesykSR9yqF9EsWKm0stfr3nz+jdJ9NxuiyK3XQYVaKTe/j0dyT
HrUfn+KzZQR7EORFO149MU9Mu9uJiTZWtykDgTFYf4PEm2V6EanKH6sdF3aYvmZ1nbm7hGvudCTX
f0FngUdmawcYLiodUUB2MWkM05b4Ww9E/vVY1cjzqQCLp6UKqIn2ZZ2euYYgZFIwhxLmOqPuadts
62MXb8vXCl0ne13PsPjzcy3Ral4ml7MBWkSFXx5EOxEKzA0XuBP62iVeZqQ9uewbtoVdpD4WlVdw
vwsij9y4wgXgnL6Yq8ezWDoPc5D5C0KHPQse+VQH2+PYprnraXsDqcA5eTuY6hV9CvIbal+tNna+
CCxDH833Xo6Lctzc4JrMDKxUBmH7yk9nzAlxsUtj8ThA9m2fhFkdNUsmO/hNcBlqWvtRooqqJ56d
5Bo5jJNL5APqhyei7gaywu+S9Rwyy2F8YHsoZvC9oDhLrJ7Hb+/tmFOblbpeZHV8YVy/JCKe2Dkv
6PRpz15Ej1wpajW8OnSURt3kW274jBBRPE0KdG1nO7vt+g4Le9xFlCCwCIkkeywxZ55PUyPPPy1k
xTmM50M/GcnwSIBF6CQrOuCvUkdg8HgFmOt1ItLgOHRXi3If+Hrk/TCPCjEpm8KOo4Ly6Vjd3qin
1Ko/2NV2ff9Pq2u/HtprnirugM/qaME0NvpPWZAhOOP7aVK6DDjx4PgCJZRWJ8DsX79xln2fdT+j
M4AS0+1E+ramjgW7RKTa7owbnGwryDjLf68XaMLPOBFSHuJA+WoneD/y95nl6BOwb3/5/C5eTqx2
i42uU3m2JYn4gm1/ap2WShEMkA2oQ5UdnaZSMZGj/1a+JyW/B+GhdLYc9A0Z7Kl8STL/Sr3gVrb+
fb0g+7JBpAHuvluS2nNhx9Ml53f/oHaAzcm3mwPVMvLtvtPd+9dWmr+rJA0206Ht5XzyBuEPy4bh
mJyERXE1vn81BAl+QTfo7PiWEV6CzLoEKrgPGqyXldAVjHHLU0rN+R1zZg9J4GQFRggMq7xKwpjw
bBbPAJmLW1QS2u+2iioYRYDunw+c8jbJ6DJFY5AqNaDgXrFkIW8B35Xy+eJ2waqMMhsAXmIp0I7j
wbmHUgVVcTa2IXe67SE7jl7kP4+Z0ICUIPDz0vh5pox1Xb8haGAS/IcwER9W11Ibf3OWscffAodc
ucvw1leyuvg+61O+IuW1pAQLKZXDSznIGnklsgEH88xGIOS5uVOcFpS5NdaL2X0NTye3yFWax3t8
jUPaOzBpZ3kA6mLYtAucUJTeMn/2XSl3EJrkKYohUGCAi50f1cmUjnLEZKw1SWOQcAryJfb1PDLJ
i24xH8WqeT2f/Cn8SfAmS2f6UYnzKj8Dxob3EzK6fF+vkXesCNxyPLwr6fzv6+nDRnIXOye6i7Of
xd7ZW67EZ6pPUklyYzZA2IHcwl4Of7UpUWsaTuBGZsemGj2OwfddMmSkbff15Ioq5BLOsfOYJiwv
Jv9ScHEBEMcBO9vyxOL345XGnt246ELH/JC23ThTYKrDmfR13OOKhc4669er6nfUAOlWRWpF9kNA
a3EXqgpj5LCXO/+LSmHuuWL8v21TqPJjYmFu86N98V+oJWI5awBoeWWL5jlmzaQLpMNc6rYww6wM
yAy3/koYTVrn1XfVZUSUPX0HGbti2lFpTrGL8CwtAy7/QQnxiad8BESi3100cABjd8NQdcKq/3Px
OGCe7A4QqrSU3oF6mVGXtotvfYrelTlFwEoriSMRZsmpAYba4XR1gWxtrJrAdUa+ET3XUr16OyNE
lMedU59zZ1NW8Tcm9Mj6jYZuRhV6rWHpk5JYPRQ9Ro/1Gdi6HJF9ob2RLDynwPWLCQQegGKv7rmB
EnsEV2LQk5YeFzySzz7SRgd0yY1rafdko+BkuYW1X/sjxrKPgjABQMynJ11wPbFo9/jP/VNF8tkK
POGjCL8zTFGzMLH3TtWbLb4z/ncW/aw57Hbpu6fE5T6qYv7I0DpCdblyq/D8iiXIyamsgtZTBQqR
blKejD0FaPeGAFJ+BXbX7+ZwrVeYbqQSCsdzdCHf0pOl62wdd6MwN4husrn7wDUVvpOvWdu1OZnZ
ui+Jw8NgLBvyvojRKiV+FvWLQgiB6FvPsPev/GwfIiLBKMuCgsdnYt0u+IQSgCfXANFLIm1cLW7M
lv5jSdDn4t99ghq3mnftCt2QgQ3M7HCOuxNbnpEG6iW+FTF1QLnXXCvDUNMlKLE4eQihi5EXAOj2
l7ugMXchuwHBanwKKjMOp/qTAWoEGQYrB/lsCreGS/qa+STy04g2aPBkYjgl1pkxLcFX9ixCRGa4
Nz8VJ9NqLY1wkhFLwLllbr1HxeFt0C4Pjh8FqwS50SHL45IS/2t2TWe7hjw4UF2QB9Z2fEjyZnQs
YIutexGQFMjTHPoWJZsStTI5lDL4RS6e6FzIt/tibt1CoHaU5scv71b7Ea10T7agb/rDziJ8Hk9t
grB1TKUmjRBog5SSE5gzN5nk67SzfQcxA0a2a9RDGSm+fU8zPvCucO/QXu9BS6qplH9ESRVn5ROj
yuLLRzoEit4Urg9h26BOawUzf7T/pjhKtiziQvS5HKZy0MaNXzkbR6BjuL9qc9tus506QoFPFpLN
5ya3JlepGM/ZJNcAokdv0c+zmiI7nvZ0cTgLOKOQTsZthBSvCQvsF6F5pb8Uo+nmscAxrdLxKET7
CRPIK3xO3v6H+8zMGY/tgtOhU0gf0d4yEmyzrzp8GCUZCGlx8oUYmgRyXNSnSwjQVkOZMLFlWANg
NTJ6XAtUA3wWsFOFRbPZBIMKnqWPnkYya1cGuw6tb046Q5weROAzVBedkwcD8RP7HdeV63xng6RH
pVSsrc4R1a9BtL0Bk7rbn2I+3GkRVyXBb6sKpJRQ6wBH8w7oFQOTRHqge3RxC0JDClt+Xu2zc2no
s+IFVRLDct14O33Enx1PCeJf4Ccodfrd8ElpXE+IJVZGb3JclgKEcRBMstj7nsqFT65bDxVYru75
lGXRveHnmPYprFvbJOghkAVXaSjbqOsmwthifDPGHN8NjUAoZDPLMpZREMxdvg7I9X064ta+18CK
YxzDX8AEe7zCqOGSMl3wzwUToQjiOZSKN2q7atle+JbiPuM2hgUmxkBOtUuT35eMgzpTH3P+/3zR
ESNuG8O016gt5GYvRuogAx57q144kDYlDaLR06p7fmt4MvlwV+E9CyDxzj417GsUiaqV8kUNY02h
n87Pw+nseusxQAWc1rAa0xcO0923ZOYkq+5sZK5hl5bS6YBzBFmyNZ2nnBMbXvgTZCBcaNezGkql
ozQzpxhB8eL3gNT4xiaInBKB/llMl3/bX3vf+9tPt7TS+Gf6RJrBSnjsQEB5+G2Q+vnnSAHwVdn+
dxCpyxZPU0LeOF/ngNCu8enVmvpDYWMTgPp6khkZF+VecHAFaUSzKKlWqa1ttscQwToFMIVFpIrF
koSvNVHscnnuOeRyGkgLAVJkr45kWK05MeSBxbS1Ljw7xcqe2241DiF1+/FYEY102kZMXehRbCoV
xViD53xmlrW/CGxNgcTl8mqzG0ZbPiifKCoAGajTxue8T5Zaj/oFNUSUGuXjFMUTxx1e6kgr124O
wHg45JEpb7RoJIN2JuhjlJsWB6v6GdKqxCPsWuTpLXXpCXaoLFXQ1bYQifdPxyOtbe0WCFdvS+v6
wWXVBZGiV144gkd3kvlDxDlWuUW+7u5nQkxFlp5mD8PeWdqB1iyKoZD3V8LLujU4ENWBYoJc7BsY
gwfGaWsAGsRHrUHfoDhokFLi/UA231G9nSAhA2d/I1vcGnEjdPk9WPXKzFYfXhKocrukDk67En50
gCN4E86R/MnjcCp8gbCXxWiTr+uZRoMh/xlbOX9cr2IKSEdaEaJ0Tc9Vj7qZf+mbFFIC4aMPbl0a
ros8akXODn7dVjcaaD1fJZOxeVNoxuyajd+WbsMgoewNAC5JR0VE1dj4Qeubau31WvZ+qP0wmbHV
BQMHCI/CWQvlcoGBsNqEuVz9rDt6YaFodif/eFjgoBSF6wobCOg1ovjWv/dCuHGwo/d1w+pGHTlh
y9YCIB4M3WFk+/mkTsZnbQuLLG5afa3OYQAapMIF20whH24YXl4Yq/0VwrAseHdW0SvpdzFk+Zmj
mUT2hS7C5Skfd0Nz/5GBSuiLdW3BljiV0H6A18rQIWiFpORXTis3+IFnV/Zt1qme+fi1odu+5/yn
c+LNOKsOhXbC/8CWRTDS7fst+HJ28kEA58mJ3Y88P+xLmtIMzKFVOCHJaeTOKAAiYLy7kJSwQ8xt
d7Y7mu0PFVwwZtxLQ6lwcV1YNs+EjSweu574Mn03ft4x357CQMgrPDpqRuQ2wGg3bCuEycMDbyqJ
fNIMm3lxyfsUWi5qnHl22E43CUrS3NRYYmpY9QF4Dy/KMmLFdRGsB0liaAGb93Zcwe5eFzycBgqv
AUoon7Au1qU+RsYveJIKXMWrUouXQb6E6U9Kw3/i895fVTouFxPXLYfXbLPkR90Qbwt69MpX+kkH
gCJapbLAadNhnIka/e+mOUA2iBdO4WstmfMDj7JGa1m7Thkr4LPT+0SVuy3C5zJcZbWwDqY8m76n
Zpw6Q1pQoq6uDX0bQ2BLkoDMsGSUqAfIOrsLh+/p0ZTGi33mhAopzyH15qbMjfB5rTbKbO6Bx0Bb
DFEe5zqgLsB/IXztYGnkMf+oKp3vrw1b90NBVdyltAcPbSZ7EU+MUpde5Uprp4fk5scyH2ox/HV2
m7erAukjIbEpXixXFErlCoh+aSKgK2Pn9Z81YGDwHX4qvbCvExiq1ZODapXIwdRVvlMMmUW5oznO
bDY7/tGzpbaLE4WopC9/1lQgnV4qWvdlrWfyYDGip+KZxTfuCHJgKpTZ37nN5MuZwITblolUjSwr
7IY+7L5QmYDEmzZT1C3tljPyTANTXeIo/pRCQAh4cpMO7n3VudREPLBTu+TyspUJWQGmfFJs0s4H
GmTG428Qkmwa+PIeujiWoTlhY0J+eq4ulNLgruwB0oAKKzbbdI68KPvdQ0182OmKf0sc8WMFcDaN
WsoF5FnwirTJw6jlKLV+JW2v07WNFnlkgBTAsiMeciY1tXmI2ac4VAh8QlZi8VPzDDlY7rDpDEc4
x6MBvHcB/VCZe9saOUweLp9foEfK1LoFosGq+nd60Lm9oZo4UB8USPvuEqEg8/DYdC0eWIBy68Tv
Q0CD2pK5fQsAYz6K8ujL100t9Q+ZV5ScDzrH0n4TxfbZVB35V1bOapOFf/kg0245Oy68DomRFnz/
/ZjMjxhbdznwavQGqqgB/+Z5U4TOWQ3uS6kFGogAxgMp4M7S0DIngROCTJwhY9pBVX1Mn+8Cj9b5
pn7/QpWe72fquwAqxMN5nKwBVgTj1gWT08S82wllJhGmXyk+DDw9Zy/KGwJszRPaEyWEuXkeXxRo
K7nVp17nSUZkejn24VQZGx3/VC9YaQRTPX4g/eFnYt6rNIxUM4Pgu8rkLqouwAk2Nx44eJymzW7g
HYYUC7RZoLAK6qYeliRsjHroNeuFDhbYldSpMPd2jboBOsynCX7YjHlkZtuqmfXw/+ECZ9i+L+U1
cYX8Ox8FwgZs5Es/ph99Qpt/Qs3Gp9A53xKqD7VB1b7zcr+uy2mxGGdYx12e1uOqPkgRAtQnFHaA
mu/UIKs3+2rieauCXGx6w29Xob1i8j5H/tlXfJFcNkWg/a7E7yUCekgryUI5VBIGOa3tMapPTxBu
/pEoSqRYTLm0KInBnKi+zh7e9lxzTxKWL3pX5p4ZI/fXUI7f6YqXiahQtIAJWrbuZfBUT8PPKu5M
TYDG2IFSJn8D8WYScg6YbXmzvTNPUUNzLvwkhlUSUIaz/FJ3buLiXGJL+Opg6Q/+zASYYiMP/qqx
2bXnJHrBtdKrGhuBm/SYDuSfBQEEqkChTQoxqUGlMcClGv+3/7+JEcwAkaEKoxiupLg50ymDGaaI
c9eMV/wz124m5PuwAO40jyjXoSkWuEtnv1ZUXUcg/UdCnX6eBzHLtnaSpOnzdscMcxAoklYkf3V2
KYfDBZoBJjjirlt+9W6NaNG7AQ27LAVHvOxzFBzwlTRT9X8KRpsH79Lhnj+Oyxy+SJoCL4ZlnJy0
mhd7w+RhqWEpPOyoliBRjMlDOAIPoyouclt49lPgq6fHyd5aRY4siK2YuurL0dZWdGgejhyUq/TQ
4VGpIVxDh5mLqm/a+ISlozDMuTkIqRXag3c87i9j4HgOKKynCgLihqIkA059zBl6eoGbnN0Lw9eO
iBjQ6VWXh+toLbm9BMxFiBXVMawU5de1tezM2Y60TMbMig/ezVAywTMc2xw0ftnl6fxt+II8Cw3S
oXR3sTI9IzqiBIw8ZiV99RigCyNgtsAthibSch6xl7h+ijWH4s5r/Xcas0oMhztNb2LjKUz+Iob9
9x8rA+yNoG2aTQork7GQm+wmHAEAs3lNBx22XAa8mZhw6vxqSI7uJrtZu91LTgSucV1SpFZ3YB79
jqIe5KvmolBqGX6dHBwMEMIKh5OtMGk9JposndlqYMd9nlXsktDxYnINPCbx3r7z16E6lNFxOEwf
3Dvj2wIDDEErld1Q5ejnjljygdh3AdQycg8v4F1wPSFsm8IoUoUssYguP5VTbbJXamDE/v1YjUyI
qED/6FOHQOt2XlmbxSNj+C5iLp1dP/P8Mg3aJuIIHZ0P6vUoWJtql8CbtG9N4p43UaBPne/Po0V3
XvMGyipbHl7b/KbVaL2WIhcOLXoZC8L+g+S4IjMMSQiekAOIB6OqmnJWcQnVXb9hKj6qsbPcmABr
RKsVIs6A1pv03JFNVtVtvXuVM78IXa6lWieZU9FrnZBEm1MY+8dNTQGGIsNteXO8Ef9r1Vv0JrgX
FYH/PX1LBazCMSx2oezIFC38tESttUchbETcdDb2IKJVy51soIZ4xS0aLNxswxGnxXRng/m0Dxjs
JYDsq/NHoRcerp+X7gVhCY1WExPe8kT2Ox+Sd1W1vRWvaRVZFiD+GJfcy7HGgxJObcqxBPjf7b3I
lL75EyU+13hjt+HH6g38aox8Y9KHf3zH0aPwueekzoY21UHwCgNDC7ZZKvHLEvpHVaWp/kIFxOHY
xVvXucxLDpEoaV10BK0oN+rbx929RzykusjMGoLvguZcLLPZXA95sBJlc28BbPuCOUYoabk+tj6q
w0RNHKKo9CAANXLu9RsFj1+VlYQim6SugpepDUtzwr3QHjNAajM5KrDPr8tjrjRiBhZYmL5L7vRi
WvgTPkNWyhWV86IuThzx6KnFE4zo4imcBB1paCbXPlQ2RGUDwV08NoZ9pJhDt+n1ArOP3ulMOFwU
WRWAmzd2eDYk/9DmddiGjyqXbaruBW/xrrT9Q5PdseCNaTR0/B3FuTLzzMcgpN7y3EHtVOIqd+GN
x6ESQk6zht86jCNivzOITjN6RUhZa3tKsPU9bB5vml8l39fU164IkyJcCv+CgKYIzQZibxnckuK5
iVuH11fcPVLSfgqiz6tMa8MqK94wjXy9gBK0uiU+GeFznkuphi1FlBFq0m3ATbPX+OVMxD194UHZ
mEyGl7KKdn0OHs2ZmCIZM6xE/XZcdHZlm3IGERMB2Oyv/nveYYqF/PScIawbQBnux2gbDLLBPh0e
q4EEb9U9oDcACi/5oEWdQ2u/ObGfSrh0L5kY0OW8k8vJDY/HyWQWAoEiGODmZkm7wzFFqi8BclMd
4zBfhb3UGA26yRJ/6p50fea/nGrwj5tfTzibWVqUphPlwH0L+zhc1fxvrqLcu8fqcr7lWlsNonXE
Z7X6CIdhftd2P3NYBPkWgE2hJ+HdVo5W8H/s2e7sluwNEz+M2zwRj1kCpBeGa6z4HhVPIImi47/D
t+LyYHSGKzdMWIQ1R5Io9q8QHibErFn+QMAYzfg1FQeAIKelYGLsqlNloWhFXdAyM+7PR2GmjFue
EnAQJ4gTktO6XQ08IXyDHZ0VcLlYbugwRLb+4ImApcxiemkbxawoo2JVOgGDAYVEiKqLbKyHpX5F
X4Vt5modAIgyqiqubBusVBoKKUm/jTLUfmkplG0QcU3+g9b7zmJiXuinhYzf532zN/LnQ3RZfiEu
iqv2nhdl5iAouX3WZmKZRRmFtihf/iac3Hna85rErY8Ls6LZ0dgOAxEJvHR7F/MPShksZk6/f1OR
kRuhQpVYR9xHBcMqYUZnok7HebiMjkifNQDZvFWkqPwJKnHJuS0t0ZsWn2gB9PO+fb5FCEi+Vfgm
VIj7JaomvxU7yiiawSQQLi4gK5ZoXNIB8GpHOqIaOFe2R6hFQ3h90YH6pmoRRETF0Gzq+j4obqPM
yPoGJh6bIdvreAZCCg0ZHmDsCf6qw9u6b34SWxusakBaEmhKEcMwa6aRz4+gR32LvWjsuOd2d7DA
FZ6CxqhSiqEqyB32dWuDtMeEFVF4cEktIab4Qq9l4WjY27z5WE3on/jIvygocokRZFFsOfvTw/aY
zFWeiiVAjQXzcuuWjp2HEhI2PhMc3mYbFoFgCw1CDrsk/kGwWcB/DQhf/dku9ra03+Eg/6+EGiS4
bBcFVtVpyn4Ig5NWYKPoQc17/aWV70bpCBjOpuIVSjjnsISlHlix+mTZwEhMe+pS/znEHtdLWkpR
yDoq0nn/7j7+E4tTdI1YP1B8AfChamUMSaMIYBRIUAXZENFwp279j6iCcVzY3dds/EoXHDILNZ0+
fjI31PnZLIa0rqpF5KlNEn5vXezUmCSsDiFBiHHJTUxSHVCH8S9jP8ty9ibWL4+FHbQYGZjM+lfZ
9TQUe5on/vK9/VHZttW+jXGWi3Y5DFfXghMshgdJIqTU/+wlGBXLC7EIeX+lbXuzD/ea4nrMWnWi
Cwl1NauquQjpW35iiSr98plnw9nEk81ybLvDpndiR1Bo0S0zqXhHwF2sZHW365tO0UZSPIiA1qnJ
jOsW0LAv+DYdwooTd60NP9yd4vmoi5DqOsSWvnYBdt/63xtEpx+0wROqvLK5lTv+qV6V0WLRV/jF
eIU2d0PUd2M61tT8IsGaA4C/0nnYIyQ4tpak3+Ou3qmFenhz620oBgn/GgzFVtt6ibJfl6gWQDID
i+hNOeXTWxbSS6dmDBiu+us248YiQmuSBkNvBLQsn0l6heYDdKGcqxMAEg4AzwfyAW+EEOd5mj4K
+kCIa8LF/DLNWxeKbtsQPbEURAH40Kl6Cgtljo/Niyj4uW+FzYITWEXbXRK5KaPLHC39QIsSn7rX
+OaGRMFn0xT8h9Sg01riQPY2gDTwFBP4057OQ1FLMddWzCoaKP2ZBkPW0OxMCiAjhRSGAeuqhOrG
N3tdyhrBd5mV0IxwB6mIWdNq87xq2RYPit6vYDgk3ECkPtec7+iuRtqEylwjhzTeq0z9oaxCM2Zz
oAXS9xsNV3rfMP85AB+m9S23fb7a8B0WyDgPUv2KLf03j7NJzY1cVWS0U7z1REG3y4TPwsrIxKGH
aleHotxoakN+YOVlytP+8Nfi1L+LtfqsrSLIv7UgA1YmUWDeJpH0pRG/55dPFPv3Pe+ZxVM215Ge
XANZy1uYBfbEQhROcdbe7dmrc1UbPEJ2ZKPuGUVWzP1RKXSti49GnZQXGplzFLq35+5ds/3Suq+y
0zAbl819mhfdIkBILJEHwsA4jyH2Oz3yxTfZxBZkWS2RCri/4kiuscF2Acwo2zDiAarVspx7SqVe
uc43IIgdRoYGh5oDqxiHoPfP4Z9TkyQZIkvNOYRTGE1uW3d8lItvbEWCxYa78+FW4YnwAuS7Vm/C
cbATpP7wUoJg8boEQuZpm07V7lDlDbNhP1jmpRsnhHpxAUaqepGxMxvKElHKSHXbty+x2ZlDdR1/
VI8utZCpHTnn9SRsld4hkS+6PkfT5f0oUUTrZkQ8Vzr1fDBH2H+7Hq+MbpihiC27jzAq6/qCWBvp
lC2dJysOmA/dIvX1R7YSeujPy/jVR9tkrVsnWgovy3HZy8wWay9VXuY5Y+EO2F8bJ26Vo4hxzynw
zTPHVI2OylN+kUGzGZRRSZmxUPre1k4XXH7KD2PJrvX0zjpgoISNJSF9L9eBz2sRqibz8oQbcubR
1xmWx9xWi9x729yDvzaC7nm0RXBFVV2e4THlZlm88fNqKy0Eu3dNFcL4GN4GgZQn0Bigc+a0bC4S
RzTlx6O9NKkKiN71GeLoImRHV8n+s0gWCeIMvx/BcwFr7ksLonnkHqEiXOJw5aRqHcnAzZMaBKwM
4IJWPJKFRe61/Lyof729fWYa+0oPfemv11tWw29dcTGiFezzmeFl8r1SvEuEx0MAICFi3AdeHG5d
oS0TRKFiKJOIoJoqNGM3ssqVDfQEtiIwhwE0Z8EdY1rpv6TcaSBjQpkBhnde72bYIFpkiH3BStwN
NBsB/hPb6tyJF/XxBaRRb1TzolQ1W+2hzClgSSBNdlQcWUtoE6nWqADIipAMKI9Qq2W22nhbTHs1
qbsNL0o7tfF/YL0usD/zjxi0LtAQ4Fxp2kCqh33WJdSDWd8Ufq6kIujxX0Zbw2RPE0UnXro+0YgA
GhLYYDKqZUD5GJueVNV8QA3VmzychtxHgXg7nBMA6Nko8UkoDsF5p7Hg+4vViYY/dtWB7xYTSQc1
reZJA+jEYjrbIcfk8Y8Ju6hU9guVSY2CqOVYEqWKSehX2VMVxQ7CA+4+hofNHz+sZ1elIwqpXALO
S0RdYYguqhF1yKqVHtc8W5cLk8o96TmIDsvJ31u12nfG6iavGTEpZiBOi0xlCwavAB5NMW5qUf0w
Ao6AsyNkJjkgcr4fjoVf6kWnXZ85NUcDTpT1yYgILlKDdhxH+W6pPpnjFUcBjceRDUWvgRY4eaNA
ad/NTWFLuCiyur2zKgXaYa/vTwXyzmKn+8aPMi0ukNcLTZIr/hKIYgeq7/TUHvEY266IW5dlGyMp
F6SY2+7AkYLhwln+nzu7f4Q5Bf33ll9OyzC/mn+WxIftaI0s0a6w6U6Z64U9AwbjFTnnRphONe6c
uAybzzbpYqWPG/BzKlmPhE8Fksiuu4EKUC+ihe7EG3bYgt6aebA2agYw610wkqvH/n4naKe0VJLY
d3uCqfxEIp++hG+1eOLm7pTFeeZO8J7OO1BZIykyO+vDganQ1SNwYrWUW7Em3m7J7ZW15WTEZ4JR
eThunbLgNVj4clPw4hil0/U5pky/Qyeo9Qq6m80Qs/tyskNVZ+aMvDUUljAxC5qyPbNSzwjwHD8C
5N2r0GXUX3E7qJOsxncDGo+vWqIwT6pZsxJTWaGZGl2VEa3a653FA/ivjct2jpbagWVXCs3jRTUG
DL+gv6mawpFBQWIrUef+OhezekxEFk+iYvbj2GG/RkPQ+HJMAF60cz8ZrrzFUsMD9w11lwYF2D7M
vVtsaTxpBlMiXh6GbVTbKeAY8N8ujf/Q6zonK2MKNGtWZELj97wxpW1j4Dy6B1b1/XZViBn/XGxa
k0Zv41Z/zyiEv0UQks0smPrOxcW4JZicHXPephCkrQ6wm6z3YJoCNlKbjWHcUReCqg4V5K/IZQfN
dBjutCEnmvikpyN+S8xctfqjmtXXnybiiR7ZHAWFGlrhs3oAR5YpNB4/5XRjSemClWVZ/5zKT3IA
4zv+hx1+dNOzh/n8gOLnc6Fd/9Cqi89ICM5GyTtZWraYcaHS9SXkZWBNr5nqnmhUkKVQQEIyCGQo
yOkhXs3THA6WD+mLixuBZV+vbWWY6IcSu5t1dm4x2HytOjgnjneea6mCz6F/sJ/bBPw56rVHf9Bp
AeV5DV5bEWWDyLS3tmE0Ze1U8RHa6JmeUOuHDxJD2G6QkQIx2l8r9nnDtXWsnBMibbDdyloNh4//
GIu0UjN+5lFWBrCUwHzwlmth8l2Cigwg6mHrOibdC/em+aCTLYz61TCByGWvq/Em6N+kQXGjrLq2
6j0elUfxlTi/ilhc6NuoFZnxTi9/2K3SuZdt1+LgV5Snr73F52YwtSTuSIXbhTjI5HvOHO9IHrim
BXevGZV2zcW3MCZcLIj7NGU/oXtfwNZmq68GI6BAnSDRm6T7qlc18rqiUDp8Eit9K5O7+XoK/44D
VdXokJl27kfbhJwHkkFrFNPcRegoTJ4dPGWQx1QVFZUOspX++I1bI+rzcqTbP14fdxELlwkXHX3t
k52kDf8sRSSVMuDNpiJ+AJXYUKuTUgQTOC7qT5RxTZN3IiTvLGhdRbO8FVilHc578RKVgM22MX3D
c/o/kwMGUadLjaaF630OhZSKUhZxa3ucaPAuLQBV9m4Yu4MVuEtejSlDfv4D81YrGK6rUyIfhEvn
a4Q0JBBzFLWinubq9/5JatbrQGNP9oPUwxhV5sOar5zgedQzwi9Dpjjm3nRTmGbzfPDMnZ/zH99J
6rJCUHmzICdPZL42rGLDjEZRehUmtuRw0dN23ETEluOsSSPhVanwTcwwk4Px+cN5AfYFmIUEoybL
ZczVZgund5eQr9zdO6l+HXZT34TZn+8Cgq9Sv52Sf/KuXz0Zbi4uUezL8C5Z6TW7xS8T2s9PqNqP
IThYGTXnCCCqFTBmF+8Zm4EswGrKKAxvc5qecYGk1no+B50Kk7E0+yf1fhzz03AZd9bvmvZ031X/
9XWb3rVTn8WQf4bTiGDNO/emeZ8194V4ivFtDZelSnFhV5KfqxbcnIkILmrn9oCbs6mQs85k/ud4
QB7Q8oCZklyBhspfNsHM7EaiL5afKV3dPCFXW6KXWIoqb7f2aPZz3b5gprHvkYfAd7YCtGvGj/2s
ifsJIV/MZGImOxeLgzvc3LHsQWDah4i6+4f9Cag8OISDAVhqFyyGUjJMjOAXr3qGpiiCGQvU6MTA
52qcemWA4A7Ge4icHHQKMDnzdtlxHcDFyVqtLi+Td2yFtdx+IlfW3gxT6Wp5Yp4vO6kurV7mjOID
1n2WWwmFW5wUJUl0R05aCC8t6wFwXEBWqljAAAaD3j558ojGdBVx0EyA1aiMOVbJR/INo1SVykCg
fLkyXssJVpS4WfSucBG6tmHIn+Odt2wnUxm044Y1Jcf/zBYEA4AbPWPzTcxK97DXolvhP/0nJtjD
Wy4kBPTR2X8Wa1L0V+IHTaDfgiBDgiuDiaKAGKrr0qdrN3SvWnjvM/lK7cXJWq7eUYvtXdqDLCEU
9ljFqUidZYFvKob3XF53pP7xOxXagXM/9A9z7q1hJnytaMTk1iUeU/yXAARSTSF/d/I1tPKctvuF
u2++w/7t6J+RHTa+LMLdLFi/9Z5zouR1huhFArFliiRUzLN6+ma6lDgCGZtEDIOY0LxGZfDx81YC
jsvV17EjT0ZB/lRPVFkdA9TjyOqRv9+Tq7GuND4Cjt0X4taA7CzLXxZzrKMeKXwPonD9/YLz2Sbz
5bGJgXEsDYFfF8TNHe/OO+jJ+GYYWp2e9F9IcN6qX7gVSBgSIHKhdUlpMZom1pwbr9Afhm5m+lo7
FcuKr/zrFG09TRnALQAQHPpcbTgDpE14tSX2Y1peDIYam67Jym4ENOB3UXTNv18I/aFZo93nuh8y
yH5xLT3VwJniDZJ/GzzhftfOZ2aH87scsp36HcF8/xiR5PQskDuVKfnACtaQwK7lC511Ng2fqUbH
BVqtYZ/5ncqp3BqfYnbS9WK/T5uYYPXGvm78XPmu3Xb/pWgZaS69dJ6ut5ah6DMgER74JGwgsOgW
EtaCOAm947aYQkcyG0VmuNNDLY4wCrC3RLoqrBa2jAMoF3X5OJOmQLvGgLrW9BR2PKVk6lSCo/c1
SDRN7NZism2k3N2uFyRrodQr7Yr6Xz4FylneYffnqpbeezsxREoWPY3M3vGikZJKDB3Cq+hqkqA+
wzGBGKCkYrYj7gvozWnI3gO+foDkWXirtXvgcsZTmn9AXOAO107OvtuVTubE3vsp24k3cqrfDhfo
g4lNRhfpBS+LOm2Hxg0vtniTJwcjdd2YyEtyKE1hCL1jCoeyRRCCnZfq2O+2NyQ7dTprgd57LWLM
ObKUf0stkdtL0DO5Kx/Jf32RohlLw2xcQz4cYDkqHFci4zrSCEUDA+sP6B8m6vZsKWOm1vNebKvy
dR5dM0HJhy2PVG1fRrqQOOh41nozJ/mZ79N/BPmEmyAETUXLbv+B6/021IZIlusDU/PplOEH/LsJ
+6cY50fOTEpdfO7JcVvgK1XXcfQIhoiUyi3iW41OF4fCLw1MYpzfgMwnHGXUHrs028BL+4I55c7Q
tJBRTnzrQZ9PdnUIvk06Ud/RK6zzTh4brcp9dh4UBhZQcYYy+UX1tLuobhJQGpVXRoZrv/y0hNtA
GTlGfpEVIDpAvsJIGlRV4XOk/TNlFcZ68n3rJjiVOHJfIg6yLl2ArxEwe2MTe/zmOEAYCphNBpt/
+v6xkd9DR9ARd2G3mVskUfY/sNHBaz1qAv9DwCzpLs7KLleW49Ici4MHEb1pad4pH41cL5+Mniy8
2zle57zi2xZuDmIY16oTZ8kJ0j4f+sV1/8iXmhXeN4LfF6LaCf3D5yJCPuofYRN1fKaH8mKlGQf9
c0Ed+ssv2pnaKH+O3KwzBXbDqCC1XFkzu6VTuWkcZ3cvovXw41QWCxa7GZhNiBBnMnDiHjajUMJ6
ynmErUDgaPajEffALgWf7S2Kht9BkoXIRUQ+d5CGAuceS1fA+vCZfeJPqVGDyGlFvTuHekfo9Czc
Sz+vHUG36f/qZhCiIUtsi/8V9ILJO1EasJ8IPNP1HvaYuUTa77d1dHngQ+7wWH63iOWmCpNE+KfM
6eocIsH841VHwCpz7RiZ2KzO7HK2AnhX1VxSV8WQla7BWZqQ9OtHJHLeZuj+4DxRy4f/S4HtSwFc
aX2aSRONpxnGfuCKhiHhc89jOundEXg4qjhWUipEDoDIV1oTf6K6TCKQSnnQUire7CA0A6qBHfW/
O0UZ9KNhV1yvYwpU7vsaH+naOxIprnBYPeT9JBRzuV4f8ouIq46LocSlXktrNqHh6zNBbYsZ4bi+
dx8itcdF8kHHvzRBxmIQECBGHsvQHKcp4Urwma1HoTOBf45EZ8sMxW5PtBZ5tDz18CaPGVdsaib1
ANRnXs2U65gVUKEBDrkDzBSGA6IpdZKvGYHJ1g5fIdMZtUMsySgOkjEiVscw7h/9k34FVFHz9eXJ
MmWPediM+q/gZ/eVPWFKW+JgGpgJ91NoW70wuUaix3g81LS6TJKMMpGjOdfRqwDZlXwEm80cjZh4
cOyjQXsa+YD43lmANc29feg9T6evdgqKqJN0X9aN6RO87GceCJtyMX14EqHMVv9+2PlP5Hqyt07g
XhuxR78JGI+jTlVDOVHGpBcSehnESFS6hgjxT1VCIw41C6MH+8DKe+0QMoAYzJlVs7fmkK+70qs1
W3c9bZL2WhBFvrkVXcq8QKNczKgPeywUDl+2bS36jqUrz1/MgX86fiNId/qVwp8fu9fOzfOR+e9I
eQT6vQcmSOPPYICX2MFQpnDqneSkHlx/6LdF65RlMNrp3mO6tOAprYeghtQXV9bYcE8jCD7gwD4h
ZkViQlJT7xRITWApgqiui2sIKo7Qe5MBxJJScD7z73GFYhAeW1HtAn6UskBPEuqhbI+DFbd52WXL
DrxI+7raeQIFybQtOFAH4CicDarC8QXaCc41IoCg/PQ/lcvZQ5CZ7YSDHyJRfCRe8TG4zyMFSare
fnNByi+V+lzBIr2hyHtrya4dxpyH+bZGdExLTKeM2LcPd7v3LabfJ31h7KRaS7f1xqG/GqnBDkh0
SfV72WPnO8ITOeWvugsiTwhfH3iPwyRuI88XnS4SDYM8Ji7VnQ9Fa5w94od1QbJSyoargZile2JN
smKsMCvRpyRRXRjsKUmzxd6Y9LtzmTpHnMr6P6VoHu3xyiEusDPH0We/SsDw6KUQCJNCN/Gjw1sM
dXqiZlcYsSHRVs2MfuP2NnDTPPjsE4tLd4eAKNXhYn7+J8leEwYmfJ8y8DmLAal/JCajxx2pFWLY
M6uqwTnEaNTNtMtLffgpcZGUW/MZfXDjC+iME66CNUE33CxS89NO08N0v/u9qCkHJBsoPTqFzC39
3oRgnPlF5/Hr96bjsZeV6f0xUsEkD5BSgYV6GBE8jGj4umOiTfu6zngMlGZwlpgcn7kKNnQkiXPt
p0gvFArQ/bK2umOgzlZtnU9j5Qg3er5F/UXjP3/j1jvUSNRmYRA+GIwbZEDvvn6fsK3atE2w0tbn
+7JvWTMR5V4ScPAtjS6RulSNWE/E4kvJYLMnNZHWNp1B39kLisYIQUQo/V2pGswOzaFxn46SDhmw
lHui2+yxNWWGM5zGZ3hutdslz50B6pBXGLwXgslqnBZQ01cp68FHlUsjxjmFHL3g1zmYkJjZUbmL
GyoVtwCRcZDlXbUouLzcXvuLNtl+qb4JTnGSy5v5lVktqNAfTt/PdFHA7p6iBcnxmTFbv8B+gn3F
s495hQJj1NeYmFstFA1JEE24658zFt+5aqe1ooq++mKwl9L+Elny4bOe96N9uB0zOjpEpmdezIyA
VyM/kX3wL7XCuRd5+TUCRL5NUfL/6wkFwx+I3otxBVX94CRUA27XIx37FGbjlVT4Ro1sfg7aH/Gk
YOQCb54HiFDQ9qwH9R6YJvwonBlaePhjrITG6mgfSTPDC+L0qsPfGJhs3Y2xijAGGHKQ8be+0g2u
JvIFEdoTQiZZBio3BFsnZNJpwqsX2VMtsnLyrdA4WwugGfo9YgNWWL0AjS062X5kA/idTtHfx/BB
uoo5N0VfbIC7x6bWP8X64DhGSxekt0yTu5C2B6cL6ynoD5OwQFHwYzseZcTDBol1SsBVUvDFNkRb
Cm5aEKk6DDJjb/FLeGaP0T38zlIpo1JvVEV4JFsAyyDdumEc7uZArNN5m7LEjW0EDoD1DCGKmBHV
FBmY4SOMNMk1OwTwjdIRTzpYEn8aYU6CapI07hqwCZ5ye3WUT3eD0qw5+Jxu+w7DaIVnQIvtJZGM
uJjdOETBexnjl0qscsRzyJqVKFEQDs08UTRLosM1FoiDxwjUT5AVmAgauIzT1hRH9cBNFej4ev4X
ET/Euu4hUsoCRSdc2hj/05+78XSQVMVvetRiLy71CTw6lzu1uW55ZEXXHzJwpbZzkQIS7AZgLfo/
/soT+u2VsoYL75dm0+wofINStz80/jQg6v81722pEjbpL6IplaTRixCueJYjStNqZovU5K87XHze
i8aoYuilBioObdt+kOYyZQ9QvarTN9Rei8pztF5SR+iBZKqLtSMsgzjf+Px7IVWZU9uxWz/KcpSJ
KawkQKCNTphn06+ZGX3Bl+FkUPwipa6M1ic13F+xNO9L/+LpOk5xbhJleUTSGG5KB0nt7wHWk7Dj
sqrAiXyvNFVcNGNl3EAo2uv0d5TEIkSjDWmPhBhFna0UATra4DtDKB2Q8jlIVExu2Y+o50xnS3A2
cb3yuE848+BXcINwmVUfOpUrhfbovp7tUShrG9L5/l3lxE4g97+1tL/zORqTzEc6zZBfTMdE9o4i
kn9KDOuolnhfcI/nvDTrBqFhmMmzxtnUaN9Wp+DRK2+fTy3YgfWJ3zpTIeN4sAumMKhiWvJ7lzDp
Qb4VMFUUz4bXe5VyrnQNk7c/kB52c/Jo4Ie5e1tA6z9oxHk/NR5ZST61Wh/HITkhzfpbFoOx4zWV
ouRyqlm3DeIgG/br/A+gaIYxpzPxYO7uWi7WifsB5N6CKb+HPjEEW3YVh/4vv1yITkmSmQEXO9pL
+s4VjV7cVgnnV9A3/JjgEIYsdAWibK05MODSwFwCOmEWlgPjXU8ONrqrpsp5AtX4dfkyeepECK5E
12ZGHv5fqQkahAIydC7h9CGkCDNuh43fIelxxxKayLZ57pWclq4X5iW3DfeA8pX6eZKKRZCI3Oyt
3EOaF8Q4JWxvb/Q/DO79a6abnNi/sdZM27w3gU9IspCKpDXzei8Iha4V5BghYIWo+5oII0xB+vfC
gVMu/DxuRixvGMjDGnzB3urpD3Dm3CQvRky1g+83Q0opnsrpnND/FxdFXnJQ/9owbFc5uD9HHEwT
mDhRIJluFHFsKr/UMp11Byqr6nlOEXBkf00JF4UJx9y/lrHco0/RxfHjjiW+Ql1AObFdtio5ux1c
swL0Jmjo9IAjDvInjwKlpcuQc/EQmYsQNA1YEiobGG4YqPYPZhCzn4Jo+3zgg02cFYmGQYEk/COv
cQZtNIzToTv3KWF5Ruh3Z8wvf8PJtR9hbWJHIDBBBFxCVGXu74o4AL/l5vht1YKHIcomjKuCyKEF
6Fa8wIwqQNfQLFKE7Jdk0X+nLDYRGkRQ/1euEOu0GEcMp0YcM3LnVpOscJnJQcGpxhSFfLzR/oAG
J9IF7qNt0mkHrx/Qu4qM/kDRfHmWbkPBGVedu0TERTCqmgMt5+XRKJRJXnlY2vO+R+hS2gxahTpT
q4vKICdrhGZ84YKibeWSJEIrQ+EXwoSKGCnN3bBqvIlu6qjoprrL29FohEKzC0bS9P6mQDrkFStc
XY3BIJ54BvXooKXQD1lWrX3ne19pXhWKF6w+QIhU7cNHYsNHmrxsowcB2l38kdMPzKTX9jhDFhha
0XadmiIlww804xI1wUPluFzzNNa7N8Pwd6QSsfVj7sYqbNMEYtrRccTQHMHw6T96UpehZRj6Km39
wxZMhUCy953vp245LkwfR1rwCf6jBw/HTrZh9nkwtomkN3v8FPiQ3friSO0k2j/ZiWlELUm8YSsO
CwtyZ8kWqrzAtTn6Fhqty45ltqkUETWjtc2nJ1+iirgoZyIyjqi3S5A+bPZU67Rhn/3u4snqaQY0
Hd+x0vuGLEgeqNCRDVEqaPSaqLuu49aE74JpvNvrYXlrCRexkN2IOc8bqZD3w4i0K2EjT8fvQW2y
8bmC4wjwfywy5Mz2IZoVEzgCrjY48H4oJSHQSw0zRFWCLfjrcy8k9w42VQTKiyzqfMq+ai+WnNOe
HzEaRTTg5Bn1mNZFhIcsgC4uw86poYpa+BAcZm1nVR1F8ZxCxc7xQ42pqaEAVbDzU2mA3CF0nOo1
SNrC3SiLLczlpMJObAN0jsH8OMpfyCF41Qgb2qKtkfYgx07J7NHJNqUzXd1C2/ToZvg/9z+J3yDK
pVeoK3Z1ahO0xe02I18Xxtu+d+xCHYET3TZUhIrzyLvH1BFzQlNfndRNz3NMbqvcAouQ/Rf+kxCy
I5c/L4TQ1t0l2LYuvWpaNQ0JLz7+YJReAfI1ArMxR9KhaiwVaHdzh+KGJ8LUPM+jY3LQzr2gJ6bP
tOh03L5+NYz+drxmufXkFLAA0YVkzntq90NGXNZwthV1rxB4eNZP7yedTZFVd5JxyWvox7r5TiDl
pvhxep9Lb2c4osBqjPWILDQv288rLr8Wc1I1TssmJmzjTszkJpqP7kWiE/aKMf+QKdz2/l3U9x6G
vd4txa+KQ+owaFdq6qnFgrTF24RYWsJlSJN3uAl8CbbYce3phJtFilg7ygojHwfBu/aOCm9zt60i
eh7z/zwB48KMsvRP4jdE2FcH7OrkRxYoXP9ZNrneJiEKkvCRYhptonRgDQHiqGs8WoSAXqnRGWLj
j5EHw5Sp675Zr3PfpaqFfl/Hu2Sp26JzSf6kmb9OAea5pABYbS2M3yvl48gD+5vbN26jEer4lYdu
MMsu5xYwtv6d5u0V3VvUTKxRoQjnrqsbwQ6tOt2BpE4SiFsI9WMz4uRGEm46kjt+y1SIfGeji6xp
K0oC4s2QZ6nBaA6cW4jNbASLQJ66MGo2c0LzDg1PNlupjWWnwCncuAcNod7hwtz6RflwLG5D95Mz
//7fSlDdCRrL198mDnyDw0arBWdG4vrBYiV3EBmNX46NzRhfAeamaAsoG59DeN6DQoMcZTI0+xVo
bZVDBdCKyzFDI2D7wM53WVDKEiV2kOZOlmsu+a3dDsYmT7BGEN3biUhMJJeX4GCnwV9LL3V1HR7X
iUNfBTMaY4sWbU3ip+xzNUGY0xXp/mBmz5zZoK/4JfOb9nbyoAFHmhpqo/zPFeHSczOeiVkOu8YM
b2kH3jBIWCzCFpTTUoKqAjInfcNo/MvQxgVtakrIRgM9fbhrJvGu8OUo7fDqJT3evZcC/fNCaZDz
XVMnMdd4LTg5zZWsPFZYGj3vPxmMNhd69Wl4F3kXR2an12RQ6lBlhfJa6oNuwtHNupy8D5ufqvQo
p5tRv4AclavUjylFMechPNS0MwCSDI0Cvpf6qQ/9CxukoIzF5HE0cSxOau3CiN2Tw3b5Yq+fATbL
nH5ykrETufNAkEwOLqs6XtXsorvcdFAplWwq5h1jNz3Ea2VI+HZG/YbDTH98G8mkSNCF7nczXWa1
8IHY8uO0f2W0BypxEiSqvLx/zP5mj/1bRJ/qAbjClkurh74+on/PXVGxkTfvLFOt0KnygQO8ile7
642RbCZhZ8idALKI3dncHJ9mFlWK5i34QLvBg3yzwT0D8HOfJom9W7I+orb0TEJKpZFqxRq2KyGw
HNT7mg+/rfiVE8SFsDeeL5gu1AK2u7vVYQ+UQU5Tttks8yeyvhWJI5gMP0IQBTrR+KaRRsH1P+EX
ezboypfjEn9yvnu+0vjbUhChfoAFHx7Y7xUsErY0U69m9TIhifcbPguI9mtMX/hTAjiM2Qiw0OLH
XPIwCTBqg631/PAJ5EdEFnR8vCVtmYaw8wynT0k4dUQCTOjYIT3wq56483mme8YAHy5JR+alfG5E
wfyyDXjUzs2WDg36MXbnhWlpj8aznVpd2FCEZMsjNK2p8AXGu3x7KIV3Q4mhDNnh1hGfT1f7cVho
NVHznNiuGT/rFrKZjan/cxwFj9ySHVg+fIFF+VQBnjXTgDIqEkC+1bYtebFvc28lEeu3CkmeqvF9
Qj+jN+vZKXNpwgNlTlW4NOM2kwy0+ItBhlvdd4EcTilgGui0VRFfUXdLWgkzZM9uH+ucK4EkNCeT
LFcke06O/HyiPISLpWwUWSCXNgt85fI7pCz+g0o5IvQpqnM2hgANI/jD4v+pIjOxtualrg8XFRDs
bnf+5zW1jLZeZrS3ugrH5ZgHsssSUy2TZIC93tqHjMSpAMOXSaSZlegJJr3oQQbdappsel+/yjvE
7SeDea7LSOgXwrm5STA222gZ7uIcNqE3x68lPWz1GoEsmiCTsNli6clzpLlGSaVIEWBjfmDllIwO
2GJMWW9vs305UjwEA/8wSzHj35oK3ZfganTKBKRXKREsNQwNgNDx6J58KQRUZFhBEXgLq0kmOOpe
wxwSSZg+a69kCTjij6ndNeUJW5lxo5ggk+c0HsaATe84YA+bh/Hmqktmekvw/ezyhQbzfbenZq50
hILJ7mKS6/WvIAljXSMt8coT7LLyzv/4H9tyiOVM1UmcWLTKfhnzXuNxU5NMtSsV5E8T9bn6attv
+k63lKZ0ZY6IPrUyXE5HggArsvDkbL/ts1GVr2uMIljaqGMItmA0Po1s8EkZ48SLunlyv31808ja
o65FVv8tozxfZ1cYXzGI804JsOcDtIGf820/xEADaEEp+Lfmr2q9sp3je8oELEHRoLo4ZsRyuX69
b51OpeIjLajUV9EewZeYMOgzq3rSI8p7E+I0oNZcYAAP2/S8PcvL7k/cC5AUAT7po/BNb/GAhOwp
ZAduTGgWIvv6ZEEa94k6xIA1BZxdaaf/sCRJwL3C1w2RAJ2jQ9BO3qMRr3z8WyMYDWEQgmVPQh1C
E9eMDc27tzFhE7+TarkpUWlbWdDUXew4AoF/eQKw/CrRpCqpxxA+HBX8hI8RwyQ7tl9nCybK0SgB
+1KRCp/X1JHGLiyvW1nJ+vLrftg/t+ZdRBIzr22IZ//9DIhn91OjTNmXztzku2crZXK6rTNRBtlw
n8JT8rZODmCfRiiA9FIlluDGWFGXyHlbL3eBHy+l7NdSGNBammH9hQ7r4vgpuKBlUGGeQidCBe7V
KMiwymqXN1ijQIPZYQtkzsWrRKUiCbWXQMsHx9y6A85RrPEKrPNHWuAy94LL4PAXrkKsa8jO9AJe
o7y3RYePZc1U5sZMnMoKNhCHuCeeOvRAA1EHcMfuA3nAdcVYozm3g9vxhyRtOTJG4RtCL4oW4nM5
bE52mg5ktHjgn4KEww1OP0jrdlaS9U6ZdjLn9M/p7Soiv2i7yZHKidG2nq9iz2Mxz6cFHjsh5h51
E7hJm9Ks7jJOroRYBvez2kX38/zAzLNO3QoLdXWtZNBMSf87vsUYBEWhK2WBGOS6Kf6UTENd/TT3
O0D8EyxgqqZ7MSLw5HypMJ4LS0dwk2V/O8g++7mJMVaXHx3tfKOk/UcSSPSKZV0J+0uukXXVO+jn
LPCzSm2abZCGa9ETJRYibK1iqGnq6ktarVgKu4Hxx+RnXquZK+4oDFpgJfor1c/KTcWLsuVmKs7b
kXfgkWkL9uIUhE0cXbNue3l+l89mKmgVkR0fLcsiIE9q6jYaY3ZD9kqyKkCjBWalvT6PdHUzxi8j
2utIsqXEdIW0t6VLKtCegt+Zgwoag+B6t8tyrzsK7KZu3ASwJ2Qni3WejpI04MnCZTqI3hn87vsz
mGHBvFw1FNoilk5YFf7lYs7E0l6ZHXc3YjmQbnnMWZeIjb+vsMw94xIeFbMVYmqqnEejNTOtOFiu
cBPzwVAJM8QK/urbZPC7f3cgeQIZ/M5h1sBfC8s79nbzri/WmAh6vrHMroje5Nt+BsZnopgMU/3N
YqEYkbgpdsJ55R0rSoJ4VltrVtTSTsg3zOroD4VRBZzizAa6BC+ogpCafmpyOtlDuTjUJIKIOgO7
JMaN9BordMCk/JwThrULunKx7t7hdLkIUghrY2wAKzNwtinl6gCx68jHMMbdcPFUFZiK0FCDjVKe
Y2zHmpqBohkKajQYczS40wbxX8k2Q6keX4l44h+RHzVUML+2g49a64BoOYdgCLzl+qtMLa4mvJgH
BUXPZYDTYCKukp1kF7INqfF2kTz5zb3b7if/XM5OzqyhIRir4bkUaC042I/12xCx1I7jgBlKbzjd
ZLfF0tRSx10sau35ZwiDYxrcIBHg1QLd9NKdYZhhXOAR31uMJ+YnGxebLuZsPn2eH3tyvl6w/emN
NgSsrfyKIrwnJM43/zLehiuevdtpyE0EUe4zXXCK+yP/0feSHrZJ/sDvAsa1lKbnzoT+OmQBxpsN
Z+pAVeamQQaqA8xq26l10V04Vk+V10xfBYVw3WG7laTSrnM89iKEvrM221IdZSneiTiJkI/JSiJp
m6rg5cD3Ny74T/TFK4j4WpbcGpuPwyhP2Lr7ssJ5abo7UslYXrA6gBbCC18VijiVLy3Oa2bwUUP+
/f79IyMKZ8ezxYSzoV+LXbPCl+QrDnF+i319bqeWjm7kKHxN9O5KwwiZ4sZUrf+0bVpQRLEXRY30
7cynqOql693UxaEvZyW/xiG0Yco9iz8HhicdHNvIoW5OPi1ZyNnO9GRvsZGn3x2DU9Q9TKVLLd+c
8E1v3/G5wcxnbeYzFCW5ZgwKA91OmJFqyDefoJnMXwn3gjJMZtkZ2oklzsLt0o6MluQ4oRkeeCql
GRVwEQkuvRFPbyqFaWhHdmZZfMlUoFJxWjhvfeO/3sd9bWRJynNTsX2ojYDVrc3aNMZZym89Uze5
Ux3fVrojAgHzxMVzTTy54RKicIl7yQFfVg6Rl2ZK5ZMtteQthojOtCJjVEvEPIF1a99WI+tfVgWJ
DUGga8Qngh1+g1Ijiv/9MVslOeak/Uo2Tygx+AWI6RLjKFpMc7EYuMXqov97CwKHNJwqroOJqaEE
KHDlt5XV/Tb2zq3G0vftp5QWtZnDNt+vD3kpcNi0OCgMbsQc8tBqudDp98MI7JNiWeb/eZ2t5+nz
EXL6xtslqBIDaRUMa7K1Rlzu7S/vy+D1dn/aeKY/MaiEoir2FlaMY4iN//LDCmVZZGFt8kGUYAls
ENj8fDgJ84PWd2G3z1r1fI+PVSL4Bnnh1NVWHJwJn0kldLrOU8Agj2okhxdQKevioLS0STKR0sIB
M+vEK69NqVHtWN+zrR5WJ/tAnQlqXKhPpu66I1/mA5B6t4rolDBh9RKeVTgSjZFfZqLhorAtJnTD
Wtk1br9YjFLwqA5WmLYRBL964VtKjS9r5X0MOT7i9wew4CLdsJeoSH62VII0+/G1NUoRGCcWwxgJ
ObO9ClbbO9RGeQztP8kUb14UDseD/6UQMv2oW4TzFZic5l4DEXnKESKrgZXyR3WaC5damGI9G6uS
ikk0cY0/sZw4bN0MED8nYxgCtffkUivSeEf0ar5fI/c9XbrHQfed6FJIye3ZEMdAtuhp2LscYDMw
hXLjHE6rXXE8U3uQgmIhNGPOuvOKC1bQycwpIy0H9fzOhhS6cCn3wklbdwa7ztUlpjBaP8MWhs1t
fbWkfQvXyCSrtGnA91rSgz6vlFVK+T9clquJY0GnSwdskOQTq4G5aqLvwa3+KUKI58upGCA0cetF
jfqdQcrZqyPrl/wNLt5taWTP7vd5tpXP9e/TaCZQOQlodAQuXPjIsManJAkXAnDkRagu7MLxXDoN
hk1WPsxooqcUEcjNQM3tKcfAKRAByLzVHxRHg5s6vGoAVNVrfaJDO6TvcGc4e1CYgFxOUQ1SCXIL
mKsHM2tmVjWm5Blr8iwwwMA0Qof5EDjHn/NBx04g9S4WPhpBARypOWI1sEd3rzuEVh6qI/I/AO5o
/XUBKYu7tproHmeW1AEJAkBk3Cdsxg+CV67L3Y3qVyQ/qHgVdITH63goxvvLuVj3zBrUB+KivOye
ljv++oFly+nqL2dPBuCfjCxUp4AH8x0n5dMAn9KJFxs+J36YtNuRGar6BBP/FACZO6WiHcVPefZP
JFu0ZkHu0EqQEm8JKjcGSlOZmjP6avllcT8/owOJUjhB0lCk1A4lnjULdupAYVIh8NQrNfb1eHCc
Ey+ZXJ/ojGQ3mBjta4H4oRx+CKB2+4M8bTHQnTwh//yV7VuZ1Zlu1LbvD/vDvsiuOBHRy72BO8qX
EVO3nyVeAoD3XC3VF2lwkqmLqA4/LctmY4BOL0eaGbaCfhsF1cKp17HoEsN8zfZGPqHL5PglMK+M
fviD7aLFmEDqSyOoB+B4dN8Fts5OQI6RdVdIEUUcalPhSDG+RHiDvPeYDftlYY8m/CM02q9paLVn
/ADnPAWR5MlTqvK/K94VUkW0FVnhFV5Kz1/7IjzjahO3uyaWUdpEg9TbByrZGrMcgaLHWuV1WNa0
Cf8RK+HVjZ8t/pS09HzVXGR5xTHKryFdouBMAsKz+ZshMGJpOI57k8QINYugRHczNWEaunjsf7HY
ZDfanbqrolAV/X0IVaUd/BOZ5kRYJob839tgpEsDLuThvsF+/r1ijjZyYlgaOfTCCvQMdJzm06ux
3lElzN0Bj9WgjUO+uq1CzrOKcKRrxAvOgygJdMFpGGwsfN463l0De0oK4Srll+QOLndFkYbm7ntL
O5OuThqGPWewvGQqOnwKF9N0+VBfD95SXNeZxofRfhFwiysSnWwhhB54CaWHEgtN9dyGjzqUpvS2
abHl6eMoDhkhKNBleTsr85/iMBNWfM1uL4NuI/zidp5N+kjxzTMKWuJc21pHEL1SREfO2mKM9W8d
kG12mj8gefjZ7U+ITeiITzq0TQZmM2kHhOwgP5pKxXNkMjZdPAVAllihj4VMZJJjAGjB3QMOJEfF
F94Hn+yKNIPEnGkFz+pPxdWgX7YcByB+pqL9q09KkIxvYN0OQWg6IpRg0V71sfTs3sDKLC2tbzUc
vknque6JBgsbsRIYqEfd2JGeck64WqlYQ/QcG2rieF5DqnC5uDzzNUwv9bp7x+4hcBm7pGSEqWtH
VKhPeDu+zeJwEbs7a8ej6cliCeHW/QKkep5abqRbNYu+O1LLvNVv3TfHD6URElkRuZSUrG/if8EO
V/IyeqtwBcAexhpjJxlIDLqSTjNaJq4G4r9nRr/iiHbgPHzBNKVGOh/O6tOGEP+GQ2MHe2pb6jOp
PEXd5M9LxPq7Z1y6co89ZGtkYcZelS9uylKeoz4Q/BaYfEZpvO2L9P8bzeIAHhBYt8JbFPoNFJYq
q3PK73nngK+QdrufVA8YG1Tkx1v1gooZ0baqPdJIbE63MatSPQmeuKmEYvmo+gMDWgKElvdnqq72
bc2FUqlvAeX+3hyZIzCqBBfPwKF7lL4NAWWUOpeYZcbSox+zm3nK8lt9ClGrGaoIQtT/R1zXdfbl
GJp6RsrmUaYUDWF7jsAg7Xys7ao/v73ngUHeNe/++LHrv6aarNgGETKgimPvK+PSxQPbk/Hsxrrf
oN3zwkDpgv66a0w8bIHWkhwmzS+Vx6Rl+mLz5OLVu7sRqci9dmkqB58v2Jg4KbpVT25VVjPVeUw4
uii/ZhyAHsOk2w9gDOtrrsqNa/ob81u9g2xHoWHHzcl2Y+J4UomAA/oK0x7pNpUSY0cuBFpnaUrg
7rGbqNfBNUsNIeewH49ahKFhFebSJiiasWksD7je6p8R/hsKEAnDIiDRsh0KIoRQv9l89fep5Xi8
q0f7z/b3rWqCYcL/kM2Ez/bxC9MsMO1lwVLkt4WntAnScw5c1yu42aPd7iT+dSKKujAAXk775jrH
5GCJDZh+00rbpEPVkHpxk6GOlweW4DjSHpIy/0sP5squduc0SueTX+AjlMiG3q5p6aCSkm4v9L+j
1N48YDHm9taXNrUbbh9/Z0WwMqKo9Tyaa9xwL+kbVxf+N3cYcXIhx7jiAzww8ceq5eLzpdTTeJns
NuGhM2P78JrvLedGJQWSMmWsj6sca4ecA/6aQSnGZ3nIYF2tK1Gv7ICXZUzf7qOCwWCq2haZmVn/
e+mPa2565kmzw2KQ99KVsu7HJaoG208PmIrxeZqZssgbQWyOEGsRwi1CJfE5VJXlb87eW1OoGDAc
qhQt9KF/eDJE+ckS5AGw4X2vAflaz05QclbQ+89DlTD/+YTOCKg+WkN74rBCTK8kHxA6uwMvkhQZ
xlQvARsbP4FSNf++Ocyc+GsaypECJ9cwlHvwjuZOy4UdKgGdf9lketSCQgwdJlJS57RXp2VXdfnl
DEQMLR+c+SlnC0enrKoBYue23lfNSteflVkFF/PWjHhiPvOUxK1MydZqp+w83eyCEdNTnnSJHyDH
XD2Y1Exvo8U2pCbE21kyyt8Iof2KAP553WdSvTvIWmz/VgsAjdgFLS09Oe4pY8HnbKCuFhcVyFx1
HqrPa1CQhT1tBs6fj5NTG0zew3T1Ri4i8ytFg/Q+dy9xz3OzQHxNr+E1Blu8aL0qaa6UM48wwa8Z
7kAcGX4ljfm8NG+UCOLOjXGtA7x+gFDFCCjCc1+s/3vkVikE2Doe1cgT87tIq5lT7mjiTb8rGrf7
mlQd2bXzVYxFaE/D3OcAne7KIok3lYtB5oYBnNmuAvmObBl/pUHlH1mEo8jV/Fp0Jyb0K5FH+68d
1RyMJ8+km51CdNyO+whU9x70no+8LMSnZogaLq+G4wI9286zvnaQ1VTgN4rm+sfuF9vl6AnCbSof
znqCRH8voWflKysYThLXyd6zjhYDu3Z2bho6FeBe9CcRvM9FNyHDkMAKNPhzfubHJk5V7rWBa6eB
7YacRRIdW6ocBXQET1oasys8bjFTDaFfKiTxnI3xd0Lzt/YcjGFOQrhHfLZTxvMOJn60VC5iLslb
zWDD1eomPxMHENvh/AWeNOri4ZX8wS43xCQ5ynDnRqx71AloRDn9Ap1EK01xifqLQPvWPHs1yN/r
ok+Fm/AnHZvAeAsrcEbtAJmxpYPKBv1sPAUTWN5pQEQR1f/caFxKYhJgVznrDZQJZI1GDq7MqsK9
4qzrmnPmqCtLr0sRCeI+GuiZ9tmTgobKWbAd3lS9j+eFtPqNUMvx+Izzow7Ez2qo1K0E7xHz6naA
AKwYveZotm8Bt6KrF3ItX/kR3FDtQtQI1Fa0ML7uyNkYzyhj+llFXdnge5LD9jZcxyZsckV5ntGB
jN3+MmqngLlgzAleAZCf4vU0IsUYicZ/yQUxadGtVyyK4X1UGjXwdvYIjQqTyp2xMcGSYTpKaXLN
OlFgkUXDnTxhQW/liB21EdzEDiEgQs+jHR2Afr/eBrUQCQhEV6xv1BI51lEBSxtEb9B+hPIoe2Bs
+05W5OjitOvE1vi8P230titr+mF4rY4/K6W1HCb4VgNsecVhXBzpK0hXm+7xpy0cESz3l8Iqayku
7lJjPA6+WN2NrzGUyHxduoIjVPbyn2iHGD3beEAo6G7jfF391L2ivQH6TOKJUjmG1GHHxUaPDyoW
+cEYzKWsvW+htX/QzUd3XjDGz1doL4KTPIALMlU15Nokp2zyjRqbPFR9n8m/JMby19Y5t2TiaVcO
fKmq6D6XEAMky1ucngb300fNJvTU2E51tSzfHz7GsRK1o3YMdfUBpfrpWWkmIqhQqJ3vUg4Q5ZqO
zrZU5nlH6Z4nmAKoncTUoKxCdlOxJiEKc/NKWrBf+vynfmVRYwl05rPaLEkA4um6trTFvRlXH4/N
RrWOwmsxGdEgVlAHlJTlxpjUQow/0SPlhbTZlrJZQFnRpubdtA+hNQ8SNhb9jwB6Rev2Xie3hUZ8
EfOMbGDTavXPKBoRdcEq7RVfoHJzKCd4jRcq5gvV/qZuUPiiaH99/Q93M20oUWz9MzErbLcVeK3r
GOu9aEgNcBfWhFuivDFs4umyVy5z7pU1Q3JbtDl0Jqo4H1BYUuaop987ZN8XuyHQEv2RGk5Ktmsc
8dmX1QZRAztmhg6/jnCXNspcX8vIjU20BFPcvMdd+NNVkcvfb0Dqj34SXggCJUaNnohnHJkwG9Dg
poVZyoFa0x/P1rm5UNb8rBYCoxRBwV788LOKtKQUmfexkywXrkcZf3j3iMDBKv6rqb8ncF/cTL5B
MPfxm+k4QEsBXRxRtcF3NQg9ODyASsHSh4/9QR9DqZY84D+LZ88qwN60cVteIpz82Otw8O8sx2Eb
6m3liBdIjQ00jm5DUoK5wRYF24SNhVW0f3LCdwama7R3wjr14rRbt0eZdzJD9Q34j/ALBHBLRly+
NKenO92P3IVfzxLGy00P+yk4/kta2IXgifvcWSaLyQE3KwitbwnK4wwO59PJRMnb1ZgS35/vDquv
nCbfNP4DiXFDg6RXTpVgAsNrh3ihROYubr4IRhwnksqYmV1yF1afPheGzbiY94m3tLAcWW1qrvWi
NvNIbmfeiVassdS9tUmWhyv5Nm3CiCKGwsZF3AaC4F9mMuG0UHEU5OvzRf7XlCW4ZFJy84V/OOM1
VkOM2GJIZfIXKf8Pu8VWX3lR6hCMZX1+GV2z3kKSWlrIO7feAIPeoWaWHyPRoGme3hGW+A2Eq5IA
ACS8b6z79Q4xrtEQRSG2yZJmrFmMFGwxmSuaaT0Wz08jr8YcdYMhvr50wc6khBu6jPI+H9QrntEA
M+DbwntfLdXP9ovd1owMeLuzfKo6lgew3V/0oJb+cli7Yg6emLaCXyyvMaczaoymAgV3FJhET2ch
TNQz1cSkX7wCVyHNkqJHUCyYej+a/h1lvDlgbwikB1a7dFTJrohL7zFZhX20xgmDLCPyBoJf8u3q
35+Yln89LNVlK3Yct9xL5I1/Ws7qXpLeCcybA6O3a9wSggraYulNpoAYK73SpFE4/7oEMO4TqS1E
pMctM/PXzw6PZRmCutBfBe9RdldQBSRIjwyh4eXX9Zu1zkL7VYnDLe+wrT/KqKfpEAc9C/qr5Mrq
LeGRqPDlejQjR40Ehb8iiL45uCf/lVkGRZx/8ed2wRCOBK/IYqy0ErdsvJN+0Cjg2rMq6Y008WKa
DmYYG3f0CWd7UtJR6fXDgcGD8jB8hfo9pGVdp11jBnUnvmyZsGp5UkFrMI6U5dFnGZQjvX14Qp++
A7aN2JGKanSLn81lB0DPBt2zzG48cf9zIPX9klPTJuLsDWrJ2akg2Qhzyo6EZ+cVo4cmfD5HXrvz
TD/zbWUOePpt3AMmkreQLJytaJ+5w8EtcvSxV3tOg/HgjnI4/0P+tDwA9jCJVkDGObwX9xwva33u
OrmCp6uTVpYlhyrNP4aSW5tsjaJzrKQTR8BSl/3+EJ1ruh5ECXSyMyx9Uo/3Q2+iZZ5evbWsofF7
lkmqYXDzcsGqkvCZ7xccVqsHoIDXZVjcIH1hcY/1rdN69qr9uUiYUYY8hWiD5tTRa02PyDOe5LqR
0b9HZIeTXJT+flrGQobKUkC5rlwwepEJgSjPyKNULRZqtISXe3P+YhVEm1kU/sCcFc/iCa1BnvyE
SCcR3VJr1KrkcJD9tFnE7bE5BI3F1N8Jq1BgY6DaEir/E+rAiNYmEea78aH7BmaPsWsnLTHYQNeS
4B+3F72vmahMGiGSMHdQkQXe1yDvCHFoCHQFRspBvihwHdqaDL0j5dr69qXugT+awtgFomLw3U0N
D/e8lQWPogJccJtAoL05tCChchVyxrOPd1OK7UHaGazGKM8YfMWh4nUACipuwHv1o8ibG3dN/NmP
5ewX5vI960igZ5VyWbDv2U/W/X//VAEtQWm0bLy5Fex7uukgsdEs0cYpZXV+JulGkH4jS1FYlpT8
lWBDAKMlHulqnnf24uV+ir2tqYscIu/60rQb7fvSoqltMoH+WCObzm4zCClPMu3LTZLsJrOA/AME
w/s90DIny9BaKf8h3dNX6Y39J6OuEprSvHtar0fg7idaa1TUPGvRpSKDPm3cOqmLGGdZ/KzI+J3Y
N3TRt7vL59wLGaqKdcXKfmTj9WDKTW4gRk8T2J+bANsrpKku3NZZLC1PgLjtaknymw2wmA/A3y7a
14TSfjq59fp9f6BBvTzs74DoXDhO7IHq2C6sZU3JujZz+Wp0YmCJKq9c8ztA7lEJCGKgJ+cKEDDh
wUFNoKYZU0WM98HmyWZr3uoOH7PdieoyNJcRXQWZlNHDemjbHOu2C9mweRO4RuFa6Ydwi4ts1t5Z
VTpIQ+kKm/u4gCHZfqh0ngDZSbYrjvR9eTjzNZJQRVl8vzHuTQ8CnbHlvhj5w+cnnwOJaMZ3FRVb
DIOzH6jkCTnSW/GgBE1/e2IMdEmvDXWyayLXytuP5P774VAtCjQMprTzfhw5cy2YMWI3cCEYO3Wq
Vh+Q4ukz0xWueTwktTt3eRjxApmz0vYEry2+1XuVZ//HuKbz/sGejuHqK5g0kJxFaZsZ/+GHibi+
dxSqjIz3CBroQnhyVWFMBpVuIUJYpDmyMmct79pZchzKyNRovXZjr49Fd46AXbG5kKZyZlVFAkP6
mhQrASyqZRJJ2yTpMVt2u/cs6FC/zK7Mn9atoFQUQ1409IvIGbAM8qLNewLLYdFG8gp1RDX8H0HS
hNErIJcEPrg9Oo2qHlPE/nN3/CrsaenXTuRaY1bef6NtaLWjHBiwG4dDJVh/sCrYrh2Cdcn2NhMR
MH2k4nraHGGMbniOw/i8NX7NDzsuLyQ28ZCKETyyHDvcn8mrX6P9JpJ+91YsKlKYBupNobt3B23+
XxIYLld21jXetV9+ZVh/gfMsyJs8XM0eogjNLde1S8C3lBUHJutkYJIkZ9mh/ZJYc9sIkDk0ZtkV
ovXy5HWT9pPZ9XCaiUn9NTWJzJTEkznf5zgaeqqEfXIij0JV2gf+yLoCtiUvUkgmyQXNCtNmcUfd
QjIWmJQ/GPjbNsjktBzyLvmwc1JDAxq5wrj4nsjPIIutvGEA7C+0Ld3yVn2oByTAhb+FCPV0/obk
cjjhRXIrhmaLqcv9VhzBfyeyaoEEKd2wFZNu+Zqi0QCi1W/+YzIISR0rVlwMaVH0VxLupTykr1zU
2x2VWCM1vl4hg1yfikBqDgS7frUb/RbgQNYs8BXiFNhWoqCbHX9G+HmlgZRmfniUO4UrUQbt/FSl
VIdfVdZ6zCMXG2uNEHEFYSo4bqEXhpGnl5D4da0ZJ7+EDcZEdn103/Ux+J5bISVD+eQAn/SSU0fv
elN4+oSlqQXuTYWNSn2ipfEOplozD4xALGllIEdolXyMj4Cw7kYvBVhB/QEAPTAJJVFLBbWBjZYB
hIpOK02YQoHrmMeJx/TKE4bSVQWZbLYLcB58a5AtSLhuz87gmMYJveWHT4nbIs+OSEE/9yAAS5KD
0bAO6+YLNrPUUKzvI8BNpiBv5URtJKbIY3azhKZRHR+O8tRzqqiKXRe4Bgf6YFYw9nkEGJDJ1VKX
Th+IIUyg5/BM7TYtbGd0aL/ab/QN/Q6cpL0irfrMbLnxNX0mDx3etKeVP6rLdv4273U9u3twB6Af
WRAh3cEkBkHdQglRx7NDWjVsGxpLNthAbGbEua5hdJvvJrXu3bxH1kdiK6C0U3jQeJNMl51KYpV4
UnbS8tBt1W4pD0+KYXLrkvs9TvWS3zpTAarD48CvmZqToEMzg1VfQbxHTkB40R/hBpEjEM1H2S2A
465lSn501HLFSdYp/pab+Ib9ykX9dIMsq4DvK+KV/FYLjFQ+uhFk2TyMc/EddHY66ytZBRPb0inZ
PPGlG/MvmIGnecVZGOpbvZww/KDtuZ11naDfLBFkzq5FG/BAY13Ms3XE9EdL8xl4hBY8x3cyXRzj
V/Kc3NZW6mFbQWQPnIeE5eY/BdUZ7BVygp2EE1aHHw5UyEEMb5tU9RC7TeNLeGvY3VQtfZowMj3c
uJYmhLlo9ucnVSSf5OIP8EhiI9PEVS/Q+Pq+3+fQ/jFpJQfv4falzuoNFHh/GdZPQnpZY/JvtKJr
Q2RPLJIbTgBIVGidZQ8DatUziJVswC2BhqAhpfLVB/1DH2OYjHq+oRuapKPsEz0OoS2VmjuYOPLT
pG5CAQiSUBb/zF+GGKiYAY6hHMV00wiobX15KLFZ9D3aZllsYx9o4StRcSNOHibRjhHlxlqj7mXE
li9Sajr8rbW2rvunYhMbYQHPbm7BmrVfvfwiMy+BQtp/xqyQDIINtEOOjHFuFJWV7XIsM8rXLEzJ
WtSKF7X3iFXA/Wfe54uMau4g5Kcyq2jdKlGLMWoiigKf9ngtSJm0YojviCiF6WdK7oEUrnF9/mGi
+VGzlOTgNb8O/LnH57ZKFDXP6ENhg96Y0vVBHO4zw5+CxaD0i41UiOBJNs6bdXjulgGGHCMPtzDy
kGH1EpELbNLqU/s43v/ZICBCA2kpJ8yKz4r6bysnJS5fVts0MItV++SFOhuk0Hc46i1Z5wRjWKEA
BiVQtYHCuiKuK7ZttFYqdSzeX9rbErsOQCT7kId+my1dWZnJfHn8sEnza5j8eU4htgxgi/d6GaCt
qJ1448je3VI0PzAKp4rm2wCByeMuKdAq6AcMkWQBr5MOE5nlRX5zJ58YDHf+SK1aNKVmymm6E4fQ
4ZGJ9YTZOb8sAXqo9aAlmGvvUiZ52qNEAq/iCgQEjgQ1m8VEd+sam06nQP803Jq9eFEEw0TQtIzY
m0BcwcODSBm/n+a6qRBwLRscJz/BZ5WaF5Dxphdj0rrzWmUZthUypZyTUcqHcf72bUsI0EQL6WWi
7iNA1iKoMqoXV+IifX51oR5UZU/z6T7rMR3F+SEd7DG2XpEuJd4bPTXfOydMD9zXr1+VbNwCP+uf
ZQ39E09r0yT7n6ueI85ykzakDCtB4kuGpUm4OF/u2XEb7j26voo/zqtnY04t9Mwnfan9Ww0Fp+Mc
O9YgMU0PbhBRagcWcBIoHsdvL7iNWL6Dlbhqq178Tmoe+q1PyTvFLVBN9axEuEOht4c7YR3x184G
rRJBR7MEVdheXjrGuRUYbg7LQBW9VqETipICZd0cBW9WAbVA+Nr9rsX308/xul0C2CAF5iOKXSsy
4J7l6210AIXqd76hBOfYNTIjSSfKJTtCPVgfYpp52j6DnQW9GYQajKreirP/iN9rkqgVmdtVBhz8
tVXYXHJcaFwA2rBJX0Ja8Ep0w4WYxc0mToZS4a2sbDCmfMb1nAkmdTrIbs3uYjHD4DeJptD0CNOu
zXbWwhW+h1WjFlZkOzefKZh6lcLLGt3YuNnovf4xya3+1mgiiLWC7XMSg+sRFJByqiyI1m/IAGac
UNSeOq6v710H2gcxxjWMNi/PyCZCUzUngRDE2YNG96qf7DG/UbuKLtbdH8rg2bI5lKPqaXKLU7Wk
J61oCG93F5/sZwv+8oq9o/Txusm1nRTgX+R7kYBiqVCytkJiGOjKJWQK6/MV82oG7p1977WVWoGE
caGm/3QPwkBFEXWOAnDWESo0quTT+j7SQ1zIqOR2frw++qfy/mSHsQrfYtSuyN1VZsIjCecqB7Wn
IdeBmr3cLNC9Ko5D/9AEjf6wMY/y5z9Jw8YQCGWEO/wdSujRpyKvbxW/WLfOx/YBrAXZtNTQQAAG
+/AWSxU38q572bv/e9lT49WTce8M77NRTgsmQ5PivFZPJeHTCNbZUrDphkFLM733c7DyAXHpPIrH
4SsJw2uygUkKzYKpp1lo85R+45y2+oSv7rAkLrtaSrmPw/SjV/SiztHm9tU7U6U3l0QI+dx0hEMo
QomcEBhP4lxu+FykO0gcrjI+Jl/mEAxkRrB1h2iyB2S0qNEA/vyWu1jC874ixpVl2tPZqpcUN4Sd
iVAfc15lFTKbV1oWt63boQUTYmKuNkPW4MeJ1Bcf02FBZsKHGZKMQTnhxB04x7IYT1ncGy6HDCq2
1M12KZTpp1/HatMod39k8e1TBISUNDIqmSrNEohNYexIFqdMMl9rrGF5In8ZSPpHLhnFP1rnVLEq
7uBrOhvXoAYu4HUL+2Q98BZOYWDHQ+XhnXOKjIFqrE6k6Qf0UFdE1Y4aaAhaWiBjA3rrsVnDeIT4
ttHyktCuc+eG6kN0+AhYgI1xJtmZ+yP5hfulHuSRPSeRcHz+aUAZTe0Av8Jr52IKQA4P2szMQpQB
6UEYMkJ/ygpumEt5DZRKfgKIdqvNoi1zFiJFxMn0O0MhOltfSKu8tUei9qKHiyZldzO2hxaZCp+J
e8V4FKJDVxzNwqOIvM4svgjAv8qJnZ+lYZOyrxpI0a8XT5e+SxGt+3BNdF6RUfkYwnG2G6efbi6A
mK/5+I6dWLrEViB7gLy/D8fufzP0Ur2qP3JKTHsdJGGviu8pvJIvTX+0rt5nmI8XIyq0MTYZ1Yge
UGjyq/SCY9n60fz5NipYw9XHmKuzkT+nROnDzlh4XNswdhkoloY/aadgrheA1FI4a/uA2Bwi2lai
1bjpZdr9I4hOXEwBx3yjjDEezqiz2dK0KdqJ5IhjtbWDKSLD4LyyMXD8qcBzz9TRORShXJotRDuS
vRm3DzGwtip9pI1u2UeN9wraApA6crinEIkcG3rMrWwaw/NSlkQW7oMlOvxSjATliMTLe3zAHyCp
b0Dc80/lF42kqPs1zsi6RfzljkRBjEIQKIZRwrtE+9o+Fp+j2Z1IRo0veOn2v76cPBwpHvzL+oLm
RQeOrQyMWP//h8+OQ+iK1+J5uYu9ddt9ONQqzxIIyY0lFn7hXR1sTGs7yvajeG4hjhXXF41xmjem
cTAQS/rsTBOh4Wc3+M4V0pyIXokIF2ySBM3tVqGuaB9Hf2HFT2kZSOs6ISt451iPx/zYO1tJnEqr
0T6d0aRJ4bbXm4+P4J4u3fTmMJyWcSFuw2crlP31B2KATaelzTc9ljN4XW1xP62LkPPHWWz0ZyKK
wH0cHQ9PtHmDxWTRYcUrvRFH81brziRHczI92VZHhNIS1aBPxMqWbWcxF8ksGDN2V4pBs2Lgbm0M
ZtTrbZIPC83atNwk3xC7GNowzEPbbiFN0+jilCAoVqhywlALaW5t8n05foHbtXRHc0tHdULwsyD9
6nnLx4Gv/4cBDnTU1tL/mefjB7RxyghEUrFhaSUyDKbDEqu7dqOLZ34G5JG+fY0vjGra2/rt0wwE
cEmvDaUzqstPb5mdwlMbpFNOLAQlfnnpsax3AxA1Wl3y3XNyT1Kp+7xSh+L2+L5a0NgMc0qVFcXt
iJTuk+CoQK4EZGEGeHZvyxH8M20UVAWbG54LQwE0vRnqWVkhNAEGrCaeEBL3FMndaY3m7WzIe/sr
eoXQ/DmMS64D/BDRaqVNVTgILnExSmbIrvej9v4cOOW3fUud+J6gkwGZp2keJE61xYtSiQJKtakQ
ZiRJsDV+9ksQYD7K2HpxIW6CmsX/YFF+T0IcoFp09/p9nAZSpkalxW4g3pet8/QFU9UAm/ca2MPR
2masFjmVMys/5h8SXbWashF2MSa9miwGziIFAF6RUk/4f6ymtfsmuBdyyY/XB4pDUSJalQijbksT
+jCo+x1CQS40WA2tWXxbjXit/yt4/a23lgzdWHdcIsKRDTku5LW40vUa8dVlsofeNXjkQ9QnYmio
xWgTB6SN6flBuVq1Ot5f0lvyUdmFLFt9yJXjwaFvDUnY3eROFWZQ6HmC2cUvESyNOSnQRzkP8o5p
MkQUuNCcPUl3WJsSYbjw6xNF6yi+Bh/+6hkOgaEbhuD1acCv8e1Ps+eawZIcRSh5SlT4ZbSceFFX
lrPnHUNrF4YhzjKy4Ks+Ob3fUamSo2v61P5JEP/w1mktqc8qqILGZ/dxVUdSD1eT/nQxuRMqewmh
7YVynCMcfW051OlvkgvCw+bnQHF7YmMyZZbPn1Ar8ohvxkyBZM91V5Y/Zb8+jkiW/2CjLnN4o0Ed
nqCxQTYPg/oUEQiAsxS+iFUmXkwS2CCF9hyNB+Rj4ihFnpwvUVMtVY+pUKolSirpcanQjpnJ/YfF
hzh5LyqH6gCcGtdPWOqFPCoPMtqRlp8M13+1aFs3QyZw/UM2WGG1fDxRMSB3hsgxUPPyVsrEn/+S
6w2podxnQEMXQ5DarbKTnpGmmZ+Yxr1hBimj9mNl2ktQ0w3dbU9n+nZ9VjSOe5Rhu68Az1PrcNNj
dNlGDXbqAVOmrnGoF63wHLJv+iElgNZWz2aoE7szHGonl4J5RaRkH1XYhe+hAYr45SDysBdAyVFt
pSrCs9XR5S5BLc5m4U1CXKxnTMMi0tJcGZHND+LL+E4PeKWv63fn2EnNt0fASZYQwGijUqOdFcpM
604VQWuTnzddXKPLd0Vj3EWl1OIZIZG7P21gpCX8iDQ6xYHg8V2TL+NSbmIlVF3qqQvLKJZ4yr/x
BQ+BT3mFr7vNvzsGG4Sd+mqBu7afiMthlaD/S8e2d819DWldzLV5kjw8bdy1HjuBvAK0Jh4+QDDD
daqEwNEbyikUBbw8urbUy/0epmMkqQB0JZI2FvidmlsF3tAQ4GzNJ80KFizR10VYk45up4o6cgfO
iXlc5W2c3+BUe1v2WyrT30XAgnvgkeEgGG/wFoCbUA9cTYbmNI2Vqh9XzvmShXiMO7nSaTLm/7Tq
4hGdI9V9uTzCFDN3SYta+NvZNWUoM2UgDQWUFKc3+NsQ7y0+ElOx+1DCpZ4InSVdfNpkFXHF2Z0u
6FnFRBC8hIjhZGZwzeBzUHu/J5Zu7Wrfdj9t47uAYMcRC8CYpM8JVZD0GgZpnoI/UVyiR4hgb1Q6
YN7LPkdom/FCVG5rhqbV27laz50eAx0ukT7Jtm74y56Xga2xbTuhlj8oQXr8iFy4UZwlF1g5e+D6
KTTMLK2bEhLwU4guxngSwQZYggZSKoabMA+Et231KM6tLa2lfP/o9pDZURmYEmLEy4m52gzJyKiQ
FZsho98bIOyAYnsooSQC+qeve0Sk+Vayeffvnbq2lFGozV+g33EQpS4jxxvM4CZkhwf9166CdUll
kFJluUe3wia4eXO18rbUp9a3oLWidMDgh3mHqrSpMiyCCjrP971ZlqpuVl3zpRvGW6aZuOovhloG
AU56NnI3QywQbYnyX1BT+xIxIHpxvTM/kC7YbUC9H+9G9ajBhZC5eSMb4birMotEUgkqz/op/L15
GTJdSq+Beg6IF4yUp23oUI9tUmcMt1wNKiOdeYwwwT/gm8SDYGInb8lbcxeqicyzqk3Cnah4HV5O
gScdfZVHUBsgew/Hw20kUpU/2rmnyK3NTMmX/fthtOxqn2a/vrgw6YGHxRqaxqHbAQBMOlaz5nZd
+J6VjibuQ8ofPPepJtVmDFkc5vBKo3Z7PD5kEegYyb0iXtvaOSwj4f8TlttYr+//CeagVSt0Y0Fp
4gdrUyC3z1zyWdD3EI+X88xebARPhx7l14SIXVuN2SnpNlmEl/NgR/BzYs+Q0gPEjS6Ir6MACecS
6EPE/dtADf2yYYP7Z9zn/65hoIQGa9aAW3FJcsC42Ul2+UbGiSJs4toA3AKKiTEYc6SBmG9RI8Fb
OWS29MxOBDC+xO3LDptqz7CkvwExx1c+njmodWq2xtiaSromOECTMf/HEzVI9DLTw+o1mtfhu7t8
45nohmyq+/YP+kEB1TwoTZKRj/0gYV4ElIBrH1p5AmSDByCNOo1zwuApZsPh7eBVYVWhu1GpxxJ/
+imiW7L86bE5xNjkX3cq24Cdq1ivgEQZz+XOSwAcqNoLgTo2KMYgcNPSMNfXxAvdZ2OiqwZPtJgF
FY1hzGdkhrS9TbG9cv1GWnEe47IBXTTUi8OUuIihZHqKON2yK7l1SUDBsvzw6kse6yLKRbG+RJZP
mo/ELk6hYSIB1JdMCnbptIBlZGNabdRqF5ZmF340KtakG9deSRChPgkbzQ/fRiIUYVaM+PH/pfHX
iPMh3rF1uFq6NHQVzmSZ5wz54ZQlBCbk7kkPcSAYyTWJDHVji2QbsxB8RVlJSXS5GWhbizjpuXpF
Hkn5g4Ldo5DJSrOn4WjhdKksrcr0IC+7DftrkoO9KmAgSyKu/7p8ABj/FT4fCK3FnGO0G8as7QMT
JVm9LdVfJyiRIfl1iuuGreVYAUL7xGURK5O9FNQlakXhO4SpMehwsfuhzgg/cQl/+wurnLSaLKZY
0stUN4Qa7Wb0LjIIQbKJjQhMU6kxVyUhKSSHtyry0sJORlT3bAkcbu2W4ElTMBuWH3EQFsS/+B12
+yq9XSzHXGyJBSH8rHPsmJ84dxvcnFqLWUG6mnRCr1QgYpJnvSNTtgOvx79zxCHPRblqJwNJSpdG
HNm5jsAgJ9QVvZexyn+IEwmqcszJQa57+OEFJKIKSNmxd1OGWkikPCWPs0ZIDzhlO5oZam2nEuOY
uZpbm6gjdLDTftLUl0aOtGu9ALFMa8ELmnej6R605ulmTWhXNkqZwgVvliuJLe+0jmI6f8jFbtjG
9b0DWYa0XR14gWFGzHOXOBJTgk76Eafd7p2xMbf5N5wJjHNN8mvqFK5ulD1+OXLwQd+Y0ug6CO3x
PH4hyYc4hlAwVAJ/GcDdniqoYDgiqOjBZyUktjd1luTmJqRvwaIICSkfY3no02d05MpTF4qrVmFF
PIsCln1NGzMXwJX/cYhQPpLp4CyCqAB61ppr6tIi/QWvv3wxYEG9RsfMMnndyiwglnoOTl0fjtTj
oK00O3GmHeLqI2t/8hBT+eSQKNrpbhsQQ9h8Po3NchlloD/DDiipDCvPhg4r9E8vFPjpbE7dcbfX
8SCIcWNmVz58q9+DIr5xD4hNiQ9fg02o9gieYzjm/ZH3CTXNSnWv3JoSk1WpgL4WwNXTIjUw2uoC
6SUx0CmnEGv+gEYmjpdT+4wGuTaTncG4/ZNgFiOqoppBkHh9FVSnktEAy7qv95txw4LbDJfoaKQb
l9opF6LI3rDmfVyGG/4TJ4QhxQe4ZXts6lY49/px3gCzLr7c9/H3n2Y3S9HxpBY6cXiuiMOgqGjm
hYYv1jadjUG3X0t016eA9p/o22CCRlUcN8x8FxtxuyUuFSQ4jzeWmom+8O0XM5O2yUGeHP2oqHdL
ExM07miONCZA9vN86RTZ/6IckZf06apEcGU2n+jFpnK5lwAkj2EtJplYOj6O4YroyMPRxlfHW7Cg
s1RA5OMRiPIyxnEZr+ATquM0wNE5SsscPk7mkN2XQib11K/dOxukKNuw7i+6Ya1n8QzECciQYjVr
az3UIcOGy4sLsGU3E1tI49lWOiXFbyvdCRfffpG27Ng0/7itSy3gX+N7nDisYJh0n7s4FsLuobYY
bdHPKZep8qAbbd4mJVdwL9EmBNJH2MndZ2Lqe0YileskyZo3PwbnO9mJ8cjS0WMbEqSxUaNCVwPk
7NM8eJhoJL9fa4fCbCAEqr1Oc/Zyyp51pZy3AC5g0uiblnF2kCxzmxfiXbFig85Air+cP4mBpdgP
BIAsnLRrKnLSkem/9JwpIacRFGW1jBfooJNOIVTMVSdYIkfXa8DRRkqeytmVxVWBOuDA+o3+vbdw
5QUjmc5bJLXujW1/kUToaT9i7fawwU4MmE7N6QQhDmjW30Q+sgFlK4+uJ8MYM7UFikexSlqZFKWc
kO8hXYgpTMAUvtggLMsGUHzae228XauHLUQcHDyMiYUONYHu8F7xp5T2/RaMfZYs7rdTAO44r7zR
gPWPsD0Nq5iZM2r/KPiM5udYqu7LsyvLZPBgSIYys/wRJ4Ygn3LHyzpWc0l/WRq2cknYH0Ecvdd+
W6mgYacVYc/VyjYCyds8/MrVM7Ofg7PtIvriGTutFN3TUEurCELDZxc04xb79yuFs3/EnkM1ploO
ATvUVFeN2RW7O9wkz2dSwEMnaZFbLRnjP1eNh3E8Ke26s00m/ixSROC/ypmN9N1J142BuocNEqMe
keWwtYBXkCJ6CQqxr5mRkudoOLF73UzubyufOkS7PsLTwAGABa5528+W7RtwR2ym6RwhFD8L0aAO
GrhHnh02QyULSvmkahcW2OAo0MLzJjRsWMjb1NIv8cbrODGDS5S/bagA5VPDnrZCkw6ZDw0o46My
xM7hkYntE9SQok9AL0WH4SQub5egozGJjvKRGsyj0OVJppYL51vWHZ6dgzugV5e/xkdFGDHZ2w7D
9ja3sSm9In7KeZEjR0c8gmp3fUUXLjbv/pBg12gMG4iCdIZye8Cxcz0k+OS4fdcRixpWYBOz12G1
fgj76drSmwJfGhpy4EPOFhT2G/rG0QlyV2dkm4BgO/yjkRGKFxvdcbGyk/xJThgx3LNTSrt9HROD
aba93D3R+jzABk6HlcHhHHivLG9y5aIDNEa6ZI401FoU3cl17fFSIdK2s1VA4wF5fF11Dv3rt+y3
TwJgjfXYwvDyiQ69O9tsWqG6/m6EuM4BPfXpy3H4fqRq7owABdDWHzJkUD9zi9Tm76xanru9tnBw
T7WEXzjsCRWQp6aRr/Mh1illIU42N8n6fOyo7q2bfCCHK8ZQcrtB7Xsa5x6jmkLiSTxEo9ruKowb
6GEc5nKPsRjyZn3n795/VOQ0VdD5SWWrzhSayrbMeqnu59GgYrrYAsSiAyfnFclPf3lcrvYFxLaU
nMmhNqZx3KvCgx8lSfvIBgPvoZzRG35rgCNqx5s97wIP6B2EuU2Mf0O9enN1D/F6nKavqw4ajpyI
gwnWJYshVE3+fzv4bTBX2418wh5xLEDjomB40Dn70S5V7JxmljAE3lk7Vrzu0LQOJ5QkiZFyqYTW
30IOD7U2lhl9R2Fsdxu5dDmn6j46Qx/Liqn371s4U901TynLGfPkjdroF6tCIC2IMr6+McUsi83S
blEW3rrnl5gJ0837jDv10HmqLXyTRICcfgMzQOM36qgIkHk7Ww3VX9emuShrRll8BT8lM3+45t/y
CpU8lsr6QNDvGhD2CiN4iR+lBbHlWRLSqvmE0p1WL9OMjx+ItCTkXAWvaBYcLOFwI4s4NZ8+OUMN
HA5hRYtU9DQjG43FZiSLeu9AHkDeyk22Ai0N/g5Od8roueQd+8BrqYtdNTeueKYeCxFOi1L4PSe7
pjsXsdBaDR2C0GBYndYW66upw3EyEXdui2C/vYfnQS+Pi6jBH0Wv094TR94eNKYsUlXmL5mHd4Wv
Y4JNFmrTGMzkt+QwOAQcoi2sKAHmCxsddGWyLoehYjb00I22iMogGWcXtmjSwaiqVH1dtPscEGer
uWg+j0N3FD0ar077tdNRVAelM637IqaQGCA+Thx/J7M9IaW6qn19imqu/V594GkDJh959PjKDQ1u
8KRAN+s9DTW9gC4ZbHhzrFbqWXZawiUyxH8KT1fOwBYeypLJPgXV4y732WxS8sPzH3/PQ2C1prnp
A5PmlrcxyUv5vk/9jZ2Ld5w0AD2rYUW2DonPN2lEw4fpW6qMA3Dn0wtidw8Qkvv/X59STYWyXHxP
uOI+NDA1h6h4CI0WVbybUqBF68NJ9O5XGlfsZG+8aIMlfu5d/cs1mZNrJidTgCtlUDR1MxJbeSkC
fm3xsXrjUMDC/p9YA8Sxya4T3pU9usWXo0meD6bazKXDnqFAzndQ6WqQPp/qROEwmvfKC67ZlYIQ
cA5tr4puaav5iRQ4kz9+c0/Si5kD2gYWOPCIaer/gNv4eUF1z67uqzNfDXr0GICYOBS++4abHaft
aBcSbLme8VXQRgt+AwZhdqY0TD3DQXsWMZcyEaBz1SPgzBiiosOw8fEKkmdiodEXgaDegwirnJxG
zJpYX9GvHM6ed3BKUTfe+gPSOgFLkjrPyebZnc984XgKrrCZkImdgSvgT23qq0e103xL+eljho4l
uwrv3g5d6VPnYKxsPsJXNx3NAR835bfFLDzEecw9s8+JPqLDGZ4n7WRselx0Pbnt3qwZkt+Yy25N
eivWqYztVa2VVF/+kRbtbJdmYGIEU7cuKALhrybUEiuVIVxTXZ8TmHx6Xu3Ak4oZA9hIELhUv+Y1
Ei/HcYxL61i687g1yg8MU36vAa1rXpKRbdrMtV96zXZ2Zgn+3Zu6IQ6hym7Qx+U6Kofhbx+BAeeT
Clz1CbravxkeIaI5xKIju5rXpzE9AwaEjpr8LlNQbYzpLgw8iyhFII4l46JSQ3/6wduXjEJcpuhA
AlItX1aJ+awpjKpxLMniD50rEYWqMKB+dpt54Fuz50F8OIwyKkTj8CaPOL06yrg3qROwW7qg29Nf
soCH6ESShGPldC8NNP64+krwMSgxtmMMwFx86SpH8khLStpf2RWe1btSU7k7pKP5cqCIH2oUmkDZ
Y3jTcSxTf3qxEYlac5IkYVhl0gpZn5QE9b73g3O2EHboP34fNoWZYbKmc2QmZ4luN9C6EIsdY7eT
yvPPQp5j59Ju1YecsMzKCfXWxWAoByTp/K8nJNvSMKsxSihJEt41C1zBXLGL2POq6peiVolXw2Y3
zQksqtfaVDlEcz59jFHefeo5H3rqOuxoyKf6ZGEObE5XUio+6vQJcOD1LJRd0hsENOcUlKzVddf1
XrfqwwdkR5IRU/yLySgFxc57ptyzS0/213VbaJYfa8DJmYBoL3Uo6Qgj2rIA2uVUYaGrEb9G0ScV
46OK3ydktyV6euZfqy2+MGWsykDeQvS0H/OhZer+y7TMB8dESLNpgCl8cCmvl0nzWe0tWDUTaHK4
i2mnO5NnVD0k5JPoztFyrtVV3s4peuvO6fAb6WYa9CTem+YO3f6+UGVUlq/CuZapGVAIVc1bW4eJ
cQ73u2lxTTXXHQNKntgu5NiSSWecMGdeFprDzUQ6BZD/DmCuJ8oU2E0ef4KK+Qu+4xVZz+EX8DZm
+L1PjRxL9pOmzjprKvfKMZW9wQmZB65YOFMmcD3dCzGN0pvmn8G8Yzmggvgwlg5ZoQKWSBUDD2rD
nhNY+xaDP+1Y5DgcHEPo9Rmn1/5msYqa89t9SFbMbFJoOQncL0g7LyRyETx19fA+ujXqYd22JYB4
4a+J9voYbQkeHZ3PBK4S5i9VphiVyEHsGSXLo9uAvw4moDS+w4egi1lSz+4RmJ09IZL2lBoAOPOG
lMlWtGOr1V/15akaTokkrrDfLGO6aMJ9IrfRkPuS1uAbGP+pBza/nRtm9FfCIMhN98xTm1IOup9v
GJM60KdFOrOae2erwlW7NB2JL7ENHvtLc+dVcuwe/vRNv9eZYbllFyYYZCyDrp2TL4BdVvj6HKLS
BfrE1whapRalNEHrwVTo9KCq7WjhhVIVQu+tvgKDVTiC4/kRWUsv4I5Fwq2/9EdpxaMAdCrVeBv7
tj8ZoCl//CSmUN+ur+csOvx1FROaHkUgM4CVu7TbhNKVsHLieTfnwKH283RLZlZHdosAFCzTXoDQ
grGg8WCcEvuxKKPidc9KFAFdM6FZ8Bm8Ea0bIeEx5zJn6YBmJXB+vyQhZ6PGPQpgyTur+POmzHRm
fIujO2xmdbpAU7IkMo7XM9uLPBBQTY5Zg66lfIm4qRux2DhFT/iSphmHu4eACarpU/QFzp3tHR5k
RiBXloEPv+/fTWAa4d9cjRjr7lH+fEyzBPd6+toySUrQaLQaQEZHr7OIflOqWSjgE8lye+UHNJzU
17JS3EhGaDD7EbCV/1IXWQ9MBRc6lJMs4V0QSKLxKwsrkj4tJ0Jcv6FnrMz+P2rbUYJ3e8VUgEWd
tl82yDR2SaZWIA/5AAUsjeqgN/1cn7ZjtjOrbfqLYVsy/am8iaabBX1YZUREu2rFwk2goKHFTco3
HqRhR016jAYkzPvbltMXcFM3SvApVootdBpY0sneY7pAFBcxn+inn+FuHeGsSjX6nkl8CnVRn3CH
rwsaZV5LUglU8rY6XKuYlL0nwUYf+SdOjOKNz1MgI5nyboD84TffL3JIoT8jQf+eZHzkWoXkq5gT
1Wj9h72mqvoQQURMOm6xvo4nPZyuXKAfYjefNaFJUbLllTWSFO1Epyz/Yuf0F7iPIOTuXWQkRGvW
utN/gnVDUXDx+BcKG1HbDRMooP5bu5+9zMOwwyfp/h5bjco2zs3lL+QWQlHvPfNY/2Dn1/OQ18BR
aynJSggh2pxZKShK5OzwLbg2LVUZg8qnopx1MyAFDD80Fd3LHYwLDaR223wTT51X1nq+KrO0kyYi
c0grJ+Xbjh8gM/4T1B1FlFarm9f3C+lpTzeQaCT0vINKZlbMuwLfrHTJdJpxihZQI13Qjxe9OWgq
99Xr5bi6tf5oI0ztWX99GP12Bh1a1OdOwlk4rDaZP1dphWnIFV5Q6Jfh5cg5s3i/Ti7mNH3lZ2Np
R46gtq+vRQcwjK9xRt1J1BLvfdWEJh4tQJKYjM4JIXuUy1JEodn7TuEC1PlbkE7Gn8orqgdfy/oe
51OaFaeSpfcrLUK0KqdoCm40gS4z6LRxXyegHj1st2QnIXkFFD/6Mrjlp0eaJ2tfHvXq3sS9bbji
TlLdcVvegWD5AhqL6oTT1duG/tZ8D3kfk1Cc3FTwGe5oUIlnzmF741UpLSmDVR7NxjMDM5OjXPkz
Tc+Sg0b4EaW/sv7HIxw/jfsA6mUhNIpN+jyT8GBpZZTkPfMg8R7G8arHrI4FDBIT2ewVnFiOQbYi
yoZWyEAvePXCMqqqcAwGYsIGuE2kXQPG1LvsP/78ZBqXTmboJHcop1Guar9JlIb97ezYWVTQEswB
KIIp39Iq1CEt6lFFs3o1XO0hXiwoitIegs69TkR4wQntOTsZ9qbCExHxVPsQ/7gdZjgU9kPIKPPP
gYB065zw2qT9ho9/Kyefm3L4FEjrNFxXBNkIsbIE0Ym2CRphDDb5RPAdbnIuenbMlbQKG8wxJt52
REyRF8wi4BRenu9TM41mKlvUWvlKQctHRocwR1fV8jreDwlpxU6g1J7l6uR/ZfNF0HkjWFGj6HU4
QgBc+VPkjAhlR0Uc1jS07MKHeDAU5/8lpWCWK1ya3SiuA96uDqEsyNqH4D6SpdF9/y5nuR1bVwHs
vqNChtJkfZsAk+ghs+KusGyCJ88dCK/fL6VUwZMudWZCpDxLiNfHhXxBFcoPZu/GUXlEgUETgqbk
Y/jroQVJfGxqeyL5eo3z7ugCaogIigmVJ7XZs0lpI2wnTisKhHqK5Vzu5qovrqquPz1uKcYtx8cI
9iuzThGjnDmgwOLr7mDJk7B9S0i4FKFzF65KdqQS5R70je0XZFL4NUDYFDwaYyedkD7xCeA2ZZNX
e+nmIt97CxN8z9KfjhWrPLDkuU+1egwIstewKDj+gRD0v9J/YmbRpShxX9w7p23nUsuAnPBdC7be
RtDTc4WU8iHTno2xbQhiE6oEQ6UmPX0RBtPB0UDJsTa77awrkrprsmn7WH1kddP1U3DzVMBH2+wz
gvA9iCKaH7yQDtrElEtt87+PKgLn6pSragUMpYFhwJMgtpHcipIwxhxVB6LSS+od6oFPuEETvmVD
Z/WTsgbhwj5Zdfywz2R6mSIslKxOqGVPFmBMlfTvLk1d4DEKIfzw8ZN8BJbgDsPwQObnT/h75Nyc
a93FzOQjXvvejr+R6ZOWojgBMKgFjcxxbhJt4/rphPDO2GXvBZRFxdqd3JoQAhEmxabfJLrA1+Pr
gCWYCESLHheSp1RjkgGBfiNLz7vK3YCgWmy2xNtm2tg47yYTvGY9nZ2XMo/LviikDUTanm0+S67Y
Malx/kenp0sEUbmhkRSTZ/FLkeeOxIlPGEtEi+LUd5VWXsGlcc7/eb9DPqo3Pv8iut2YsDp4DlwC
x5c44LQmCjQdaNVZd9qQUX1WFrlzZZOp6lOrfmY+hETij6ek8tWEwUJ5uNQN/YLfHdBGONsY3eq6
dMDyMvTjKKuUj3NZwZqjIdCnozvHw5pUbF6Z4bT+1E1QinfCqjIt2ZEl3y+LJP4rC2fSmNd3cCy9
V6cEMKam0ME0i7NwQCCIWcbISsYW3buE9fBtmfFIrKQK1sW6Z7WFlOhV6kWmXixkHdSwV6ZAbuyM
vO63OIABA+CC+rWKeYjgNTmHMlwb4mk0x95VAPuJHEcNBtUJXTL9ycvmeyVKYLIPniN1hhv/mR0C
w6o060glo/PjwpuiErgh7s6okcSs9llx585ZTsK1qR8dkskz1+PzU3IgdhpStnX0mzqokJN9ql9Y
r5uOiMud8u9tomU4WB6HnxcqZUxjrwzxWzlxRPqH12bYldXB2shaAxZb8tof08rYZCzy4/ncG0eK
kedmzrraAgNV3ZOax3qzOntGSA1V3HMHG2KbsSx4znsZJ7xd4/oj8KgC0u2dtv0dRNGCIEcssW2w
lqnzgRGqPCZVpqvWWdNpqNZvbT/qBVopzgUdPOLnTcUBOg0HdKDrFNGBu5JD+R3Byo3H00zoZw6M
6wO8WOmgEN3HsXry+poZ1j0KLGq+rHuOacfsACuKDrIFzV8BHJjij/DQ3X/uM2m2Fld4ZGHC2psd
hbkT2OeMzCmLFzdrK+lUv8pPNB40JsIJB9Z9c9CXfLANOANyU6AXXaBj6gBHkv9eWlN6l2Qg33t6
b+VNtTrxjV1Ucg43OzffyHmv3CeUP5q33nmJnD1ox2JE7Luc3llq4cZSsEZJ4suHLmkIMUCqqpAb
0MC7qeI8GHPKQy3wtLJcT0tMi6uvo4/KL8Gk59uHYVc/Soh326847ncqxX22tMMZY4+le8J4oUek
KpHvAr145H7JzIhQ4ZEXEvr3ZKtObtX9AoS7ZRoTrxtLrZi6SVk1/owhdn7kPYQcJd3r5fp6ngjc
d0DlZ9Qy4btuV/RUolgCrsdvUdP6J3L8ZONUdaP3WX1xdVgjj8uVESkVOAfNLUL8C1Ccjvcvl7aU
53Y7WLwfvRvAa2DdrfoXESa9v8vkewel35uNZGcZ0GkObwbs31OokiG6wQ20XaDhPAEMLqoWdSEu
fmP/HXo+oyloisrgjlKdpre74CbajSecJx2Cg7KJcTSOncZEEYEJSiiWBKKEw19NReN/ZLhWtZP5
EeF4ZVJt74IVu4gpMbpROfB0gs+uuc293QVn+4BGBRCeAxNF6QSm+CNkt/HFA3/YCIZf6Famx21w
sl8J9FLeTBaF/EA7FVGyVVX464FHUcqr9IqV0Zyq0CikrjowtDXqLFhsia0pZWI7AhUg0k8bCQy+
InWJbzB/hSZOdlTDhdCR6DHi3sJNm6zg5kzeCZk3lemoUFGG+bE4Yu8AZO118bDADH2NPC7j/g/6
eYJsSuFxIpvoHCDry3F6HBoRlX1s5WYQjXFhEF7WVzevgMqlKN5V29yP1w0aHz1I7dUgzRORY2TV
ygFr2uqu6GqnqWVbBDQX0jaFJt2/pjEmF+qddse/Am/R4uSrvrqSN4bFFy+bDaNaElV+vWUI4RwX
e3k7OKJv34jkU0BKYTEhhEtFg2qKrgvVpycDNw+gr9hVcLCxzHf8BP2nZ+yCNy2X9aZdrqO7P0Dx
5XWZBaJspTaGH71YjNYURloMe8Zq1WmNhViqgIwse9ZQtc9yXgdi3LLYotBMW9+MfggOGjwdy2RF
sC8kf4y2SDBTS0cL6Fmtqc/QE7KGAkVx0qFPV7WmDbH6Kh9BTChy8Lry24noRM+ZK8llOKWeKhat
96yjbH676FPG2VoQev4d02ZlABsFGKfBWTsOE3uNOGuzrQM1l4Si38ROj0a2s2K/43Tt24JMMQfI
JtKsemIi7itHqBUVEGNuMKYzRSgpFJ8a9CA6skjbqSWPxAXdSkBT72QpE/QEMwCjlMgJBtauYoJB
POKxMczMyYqSRZCkztpZsiBv5gacZvDwryZtRZn4E9ndYFe95/ad/vwLVDeayHlmT8PBjv3ItOgX
BbsZcQ019nqRfOi3YEWsPrYlHIVczN6vvZk7zFi+cXhqOhze9CPiehj4ZjBkGsLzX2+XSO8BHCVv
IPkHQ3ie9h8tHkOdmV2M9a8RoH4ZrM+ke64IXM55VBE9OIrxEufNnbQTXTeINWtoliasGp4Tm+jP
NachZkmblnzt4pzQtsZNhNcnAmCEa5Z0XduiZtKnjXnhWLdijo+47awPr8f16r3nPvrFkaO5juEn
FuHwp6HXuoLflDs+/slPbt0I+9iGOi5kOhK6nQYyT/0FnP0N9w9Op01RgXLVrMIKpWhetZDjqqGG
qf/YV1ECnqSDdif6YGY0PTgFUAKUdZ3H8FrtibMvcd2kJJkYNqxq3HC5oMF0MFHRoQuMLdYkvPtu
g0uU59bg/v+B7NHI+x5nX3oYvLb8h0qD4CE3ZjpXBpsLAmnuvlm3O3AAwWB1qLw90pZ5OPof7XMl
Uh4EtGJPBHX7GfzZB6VX+Kd3qN6mrpF3VzexH4W6dIYLnHH52HHYC0Sl6dJ638Vuecq8i60HkcU0
pL8iqq6++AN6Owzupi8QhTu5SxbxwT0cNHnaK7zPcb7V2QShXj2HydY7F/sXaBs8EyJC+qmDqJ+5
U/SqQKZ48IH/g05dICXv+4/xee2uCEb3BLhefwtwzOeRFHxOFY+rZW4nwVziAWLZAfUaAnKfTRq3
6470eoejeXwlRrLAPpRZw9uU8rALUQshTKNBNtEkVFI3LShLyL0IWNECUnY+hC4U+OK8rgKX1T9r
EXCPMMKgKxIUFd3p0w1nC7CvvXP+OpDUKjFHGj3cXtHdMnifd+YdlO0yZ01iojvZAUfMyJP1JwCx
IcCI0EZeDxzVmB6tvOC5Ryc2zrFZsQiSvBfYAHyVv1Zpe2OtXL0yUWdKcCY6zFZdIDSRhadOfAwZ
GDTQNxHHP4+KnpWJ5uaNP3hLBxgSb+Q9keiKfI99HPhx4AOfSYxcXIWi6nkYHCF9tSxqLPmk9DwW
j+XvJrQBAcrEtmBgXRBwmL8f69SZDLnFyCUseXhIYbBdP2W80xVbigi+bjE10gw3yFN8C2PsE6jf
uDme8ctvz2HudgUrlIKUhdtKpsTpbHH6M8VLBdXhcyx3T1og7Fyga5vhwrFUfNFbZrCZzWnw1Zux
DWnVyUmrfZ93baLZ2mP7umDq4ZP8V7hYtYZQBvFCNJ5UaE1aYcerc7Efp7ZL0CS0FHAAqwLHJ0pV
lJoZeiYio0mAzL5JjDa+fvRQnhBun52PxwLlStPQHpYaDxwZcnHNu4WHnnDQ8SfWCOTDrAP8yzsq
6zAVWgcrb8HoLQuBumc5dHl3NbdtGwj/RJK3YHCdCQ2ZRrvaMP08nM5MD4GUAEQGC52ncGPldvUV
7v0x3s6l3QaWjxz6Wpsx4E0YhawNKZqZzlO9enXsuJVSg5GAtMQos+fdhY1Yi5bmY/0maGewdCsz
dEVPEq4eQPqH1TlI3Mkh5Ac90o5MWSQk/bWRGPefa7OYT1e1HuIXQd80YIq5+7yXLMKNIa/qd7Vn
BC02OVdBc4YuJPbA10gg5WLhYXyckDc9YAzDxPYj6/cE6Ud90vdaUsQlRlD5ot8Xv7FAvRdP5BLU
s6ABU1D4ovL3Rp6dLiq2MTiZAIj+A/Fu5pqiaQUANc6KzblRZceCu3qYusrSBHLI/u0e2l/gsmuF
ujeQg9SedW6I8Pc761DAyJRc/PJr+Aogiy9CF8Iou+/SjiCcfVb5sBDWj/hn7coipDTnbX3kVWfI
3fOjQnfNJ7Op0KmWu38HIKuvcJhUWKHrhdPS5zgAXk86DRK9pXqq7MWzQYA0YazO6jHjUnu1Ugd6
8BHrvTV3Ff0FZ6SVH1oKZwnXoWBgAMe2IBaS1T69zqpHBS0wEsKWrFXUlSrT2CUOnlT4/42DyyMk
fKaYzbSEH/hgH2ci7FQN4y+0xmbZUqbcXdgysh7a3mUofAcAGy2XCS0c1sXXM73abkvPlOi9fwdX
/7oEPLaDRDio+4LWX2JKVZxYV5eS8japhVZq6nrFD3ObbZtXZSZpsB+rscsQV2VJuV2RKUG7qTmV
OwjPAls03BSrTZ3OJVx8DqAiba0ezGnjWblGZ6TtBtX7X82m3s+53jWefGqqDO7WLJtLXIbL8muB
DtkYOss65Kmk098kolv69BzQcfZl8iGoV2LPYQnkj3hHx+T7E3XZmNnwy4NSkHrNV+CPYCaODTlp
ueDwubuIvxhBFsniFwnMhdTi2B/KzdIbAV3NlGyCrGTHzBDVLADCBFAk+m3r1uu6Qobd6hcGnviW
tnJtgjKABmLjSGP0V5NxDjzCqy6HH3eyBcj5DXByZQfheX3zsjd6A2AZNokylZh/h83gQSbCBFVV
S7bvB0AC063x0dJyP4cxN3ujWiGYy5yyCDG/L9DCn9Pl1qNB/qoH2AaaY5W+FIMPVzgfoKSdliW6
miG/btgVKWHmtFn+sqlFtao7KIsUIElNCM2FVzPVt4ggWxem1ic+Gg12nsblcIVPOkRpjhMog5z3
DbzAP2Z2oBzuk9QMN3J3mp7tMDPND46ROx1LLAHjBkAyWXskEDhLlC9Q9IEC0xSk2yW38tVWxBXh
sMyd000kKUAhYuqjGmV0tSfZwaHsHSjqQksC+tzBSoOFCr+IYchT62J5rjL0zV0swq4iWuA2shxn
D3/Z7Q6o/vDFIJ5yRlEddWZ9OIUFamHRFmLlQd4wvbCqNGHRgs86kiH5bi1JaTEcYE+V9Uv5GfqH
h/mEpfZa/8XwJ6aX1/pAjO4Fx+HU69IY1YeHg8S9fTHWcQBNQGLqxe+Gl2aXk/4j7CckHI9ycJ4u
8D9RpFP8Rw1fpFHD8zCVCNMv9vK5o8X+qkn8ocJoZ93AGFP0AiFqxuXFRkCGSoPMgtx6MRBZY3y+
IZWC8IR6v5sdBmKqTOt9jjOv87VL2OhpuVgx1apl3e5Md+PSl8BwvA6fURl717OwvSHP5S4S0iG2
AlyX/BqbYvh91pEeyvshoYEka+do7ialH4Y8leUFF9WWXy2mKmGXUxsRZdzsfj7HRgDKBJib+BUp
bmQfZfbChjFz69gCH2AQ3wsnRxQcZ4zkFv9KLsVKoaM+8juTE+5fg/1r2WZ+8Q5fDxyv/q7bYCEO
dMsebvC3dFFKtx4qcB0WCIEiDnZp2kaYdbTsR5OVjy8sbm0+SDetGeYA3FiEgswSSv2IwrLbTRKG
DfNRKqziu6z0BW3zqb8/DKb50rSW0IFwJvMmHWvUSGq41vtofL8ofe1j8x6UnSt1/eQ8ZqB5tMRm
WJYYdwRGJ2OXneduN3jX9PhSRw2iOgQKl4KsmvRxpvN5y6LXqHVbeySzatMvnGUs/r+0mr2wClsd
fE+IljJSIfThcSFoOiHUhQgEnKE7udhKjTVce0TjEi5vsh1XJkIdLbwgY3Tx7xdE/9a0vWpjVUCh
Kf39wAU+GgcpLH+bUgQD/Jh6GSLuHpL0sAaoG1CbbuBcOBVHE50ZZoHzqIwx2gT6P67Xl9yUXla1
oRJ+mdFHBk8gFu69EEoT0J5gcotB6YzAxHV2/d6ubNCREA7eeow8mhhHJ+E5n/pFXRjsQeegZXIs
g1DsdZ50OkWF5KpMCMNtZ39M3Rfqad0uAzxxYABLFE46Y9oZSnKu0T65scvcclFeZPdT8wgvr0rb
Q+4ue8O43yjSPzAh1Rshl6o0jDWVys94RDtv4u6MY/bN2n7+81m4PIIVf6HBXrMhVIMcWABRphIV
TRP9wfsFsGOx2CsKq8M2vvvFv/WwKa81bZIa8dDuWBoHcYFr0Uz7szzPLH26OWD/pk2PJv+liKOb
auWz2WaZmDM6ZORxISRrfGxrGkMDVJOUKyDqj33SE/ur0ktpygx41j96iaUqWnFubWBp2ch/TR3s
7Qgen9r0LESVJvAuOZysnLyDNo/pvPwsK1m+w3/3ioyEvlk5Q7T0BnBMsqK/aNEXEI8kRYpdrPWY
pwFVf9wyDzuwDds3OV9oL+iQWFz+FCCuXnojrm+Xo0qUayKIyvNQKE6V3dStJb/FoaId3W4Is1//
sUFfQuX5UW+FKkQv6tKckFts6OGnwGCCtiEYsSwc/c8gVb8WpIZvGRBf+Y3J5aP5snbRs41cpr86
vkoHLKtAXBPXdtplE9fI55p/uHq3FNrjNClwaoa2hQEtq99YECUqwKXZZ3qsFy3QnszVqYTX5MoH
P7xHRl6RNqzsu9mqsiCZXyCgFvChLc9OBJt3J8P5G6sc0ryWqd2FfluKVhYeKCuFuZ+H6GU/Z30Z
i6Yad2zTW8ccXzx2f/USmm5e7UsofPPx4vtT/MX5rtXt+k92LM6YkXmvNRQx502SmWYX4fzcfEFg
ivPlLk1ub8svfkAhEJH1TsVECcA79Ls/5CSs7QVwdWl6tHk7y6/ahRUt541jLDeNMvSjpuA8frlU
KsaU3DUK89z8or+nEaTRkbC427FGaWYXXMXvOqT7k80HGNnPq8cNWnm7l7sEob3BoarifIC9zUMY
lDm9YK9lNYmDsKCDKkWkUN5kPcXzpP0x3dsRCb/mC4CsJatL7MLJjHOgJOw5/cfgWOvI7jF3YYuK
jn7w3OerYcvm7pvaGtN1PqBPRI3getlqZ6zZ4XcMd2N34lKVV11ZgB56IhGZZk+NTepCUO4ikpby
blEXvlPwg2DWkKymWMuawdCzdKEoSGjjs2bZTFg7w3CyxNQg8BgIKqdbICNJ6fHsiNkUYIwR7d5w
FCY1qL8vL/xMiTRLVTIrr1GSgSJgG/Liftg83MnPcj1/0hCoUiwQ0ZO4wtdrRZ4XA2ZPeEgGcjYZ
EBsB4QOqfJGwibVl68xczKhcUB8jY7n4y4uYRqJLoZTydWMcZfITes5+5pIGdWXdESewV4P1rmWl
OpCe2GfBKI57GvRpLoFEDG2uIFCnx2aTe2zha3BO6L57lJJdDr4pdlf7GJrGnpaPLHV2t6MHDXnK
w71Tojwdk+KPjEydUPBasZqI0qeV/ocH0g0w6kerY2qX8KPxW1Or3Ll+cVYV+FyXfASDvNRakGVx
aezoniXIrSj0hfDSglHtXDitRdlYl/V1BAdq47/v8QeYUnUgtWLwpRVmPr6ynh/aqMwCzrsEtN07
Vy4EaQkqZebtuQaQuk+KaRCr9w+rwc1aQKq5x7P09AMkQBmKblWdqg9LaEDsa+SbNkcuXtirhET0
DS85YZHE5CWEB283NKhrzJRz9D/v0IJ7vtSbIN98nA86kScaYQdJn6zkfQXEIDiw6YPju/VmCwPY
B2zLjRO8MEnnIcOlrp0TDUYnpvEuxTBY36aKYQD0xbddYNPJpR6mZy0vo0tYJwzCBjgcS282ljTV
B/dIMuoHD0gAF3RwHKIx1zXnsW6LpKmdX4VnQa4McdhVtrL6s5GDwj/bduaXXOByoTOdsPayeAb6
MkmokEA/5TP2QV15RlneszCVetBtmybqNxgZnBh2ueA/KHZQcUJC+kjHvVGFswbsqDwjzqm4Pztw
m9UFaP3d/dTAsUT6FeSv5MExhOrmXL0+KyPZR2Pt5ekbYbY6TBS67kq6pSDjqmY914Is1F0V4tnn
zuOISIQXtX8B97TIgtrW76MQZjIkeCrXhxl9qAWknrn+iaxsV3px6qOwUewl+kYZ2VT+cR1JWupq
gBh48ZjyGxQHmUWvXBKmfssIj/Q6syqSCxu3TmXa4iiDfk9JylGKS5OvHgvKwdYnz/I7EpuloujJ
FOL7SCwi58ZYuQaWXvMssgLfbF/wzUFgR+Ds0PhrrmdtkhrHo8bca5gm2pRV+xMNB7DMXK9rYmFq
gn6Oyo4rtJdjplqSu/syw4x4nPMnsXyRnX2NoYtUUgSSoMW10NgbDN8WthoZmd6xN+wLE8GQcWzt
ttjbZ9S0ur9q/Dh42GPdwTHqlJd3Xc3zSCfVPa4bnVvM55sRr9mnCBZaQ6DFmInXOjcclLR84Pqh
prBXdDI7LdRjzbTV4QwLmJNPNvWwIGg/m0moVfKJDXXz5FpQPMLATXdLYD1alzoGZxZjXGy3T7sV
KLbvjMloAkqAVpmV0DQzRbVmmGdOhDNRktQVfgK3UlgDA9aYgiZp1DDDYq84GA3rM/CzEn686ULb
pHYfnBxQWdkzRwJridXA+1xdjtYgCbbsNbfyWwOfwv6HXYL12f0U6l6lue4SM/7a6k0ZxnzLakTT
hAfFATnrrADA1iWtTqY2pryo1gf9JjTnXOT1pzbEJniUeC3uSX6/DzCgwWY3424HfDbuYARcq/4n
5tnF4IXfIaQ9ZPR7HTGcTQVbzHn75sArKwNU1USFjfa9tNPx6ajFp5EMIHCEn5rEFbmrOsZqFZyn
AL52h9OgzPYjLHtTQgAlwvub06zN9X6m2P2GftcnK9DjeP9rm4F+U3O302109ubmD20tlmfhmO+b
MtpiRaSDac6t136a5aQafFbSd9sC87uX3Ey/P96mNpO6zbQonkgvCNSL/La9tVq3rzxOYhsBfy9G
Iyz50dYhIN/W+0RyszqbZslSuRl9knWFDAA/LuDZRECRO06EpGb1TT3cJv/MhORzbTiSZAS7oUbh
SOs8phggQ9MWukEYyOjiw2C3341EdWV1EPaMF1ZduErGLBOAyRpEuGbWvoktDjlWWhQa52jkrmo9
IqWdMQXxd4VUdgmcHwNLvLP/t/HmGqzpixkiRyiBGR+mq4Zxks4VOQlYRqaWOWWJvpC7u6CbQWrM
hLjOD3MEZHN6PWmKuMPRTiys8n/di90Kq0lc1t41FCH8FfLkNFJSV5wa7D072yj7la9KJlE1v9EP
nXSpZkRiEJDVnqjI179FQqLrTzZbh1AjyVa5UCn2PVtyrIoxkIyERE7FrHwqKz9yKd/6cDbMMlGe
+YxdQfn/HlAL0yoygDUM/uwA6K7Rm48wPZgRd66vFgujXc7HfJJMc4fJ7lOLTk5+l44btQfI32WD
e1cI5WOpWWJA06Z9TLQV1m5wdaiO7gOa3zzEQWeU1LeQuFln73z7hLmZaYGYecx+NXFS8I8EQsCP
kKmvmiel9FN8zF76eNg/Oa22xaG/DjkJlOk85jWvqXetovHxBPNYAKpo5MAfzQoR3oGipOuDgEN+
t6rKXDYUiJ3rFQkH8qMzd+GBYvXdJwGY/WoCEHRAvQ2t9EABY6M7h2zk6Q652koQPVQZNQiDrkIM
LWtBaCGaM6ONLA+DFtkLTgGf8GESKo5xjoXr/bmfzQio0NTTZ/aD+FF4UdRkWy44zGbnI0ibTxEs
YtDf9L0X4exTe9PnixgxAtrgz6bSO/VClbqn2OPG7R+UWKzP6GeWKzBrYWdciPO06qqpF/NOWPwq
lp7U5e74lYJQIDRsnstHu7FcNmyyX0jAhRcaICtV8olBucNT7wQRIjQFM+Y6+MuMCII+CWGMYUCZ
a+/pekWmYgWuVvsC3jq3r1o2CraBxox900aYI3eZmrNk8y9t83Bxr+ixaUVHnMp8JjjRXY14dZIe
LIto0z28bGFQPQC2cJaDdfN7JfBxNjBwmcEp+9IgeIvvoU/g9hluoQJ5YSQW/xkxpZQ3EVf+/0GT
RbWFxcDvh+bYcSrYIuttDFBe6ZsxjurM+ECml1skB8Y6Z1tx9ktvQztF3kFSfgI2+0KV7oVKsAH/
th+t9N2kDrX3iQJvwWJS4JZz8LRew++YLvD4pGCWFfYA2h7QifOwyJhSrL+b8Vug/kllLAs4fvbs
Vajbar5xOsuAUI6NBYV5xnAnikruvTVLiIfdMOMYa9hlto9Ne2voqsxxGtNnnpcuDijz/iBUddQz
XPChV4BfSPMXbsSVfGVTI1XO2gRu+4J6qngvBgWVZQipzBMCLPGAp6VQGtJfgjMEikb6DuGG2lMB
nZ4BEbDOidYk3BZ61C9o13fC0gwGy6d9wXuA8ku2MIrIfPDeWdq9TwIfhI8P26XglviI98bM765R
CZeW06pvCFg0tCkOQp4ag0wCcL7korqdatbYzs8EPPPVfEWDZxp/SktAhc9f5/uciqunkzHl2UFu
HvzDw4TyYSekNh7hiiTOovRz8GSG1RkFhkqb+F0Gv/ds8/z+ev/5ktUbbYJWGkrIaqA9kDlSPLl8
qzNd7oyM9Bon82Ivq5LCj9CtyVJTFZsKLC6S7fETOph+L9sS/w/n+Z/Z3I+6JpjwIJ4FS7tEfSlF
IlSKAIzpzikmr8Q+ytOGWdbXFsIr/oTFX+pgFM1IFj908M6z9XW+WUXR0xcoso+2Hh+RHdqH0otB
HI7VcayOhmAuB+k5jTUZa5NZz4Qxjc4ftxxzIPfTmTWRiyUBRD46lCZJOGdMAOm6+VvFU/sTW0Zn
EXNcyCrw1gnbZFmgDwY0aFnPPl1GpPBHHCGaVgugl5bn0aCqZt2Bkrf20//xktLsiJBxCu7VBZr0
DRmR7xxLF9NSYBqn5JMKn3STHpxsu2SwhPjGXv/15BHFlgAycBR1lb5Xooqi/D/XxII12+f/9Qis
CF6q0ujaZUOTJw6gsyItQvEgIoqrpT6y1nZkcI0YjpLCzmrqX1HKYlS5WV/08LZ+rTVdET3ZRJgx
PrMLJUag98I3n/hoSd6fNnN7uan6Jc2hwOrJncvWTZa6XOSvdMlJLziPOOD08FI20bM65SnaHqXw
KJiUNEXOPQNYBFcVoiL5HKydNBZcu0o1GLSVB1p/+tnraFlWDgt3gu1T4khvDiB17nmTITtTLNrh
9lhOVIZlzjd/ZkPY2Uc8pK8AmjTxOdutzgRuQUHsrlgl3iMPI+RCbJ9R3iUWCoWj3qqwrKL7rzcc
3TNntFweP2C4fSiQenN+dfQyjneyaLaXDGVDoOY9CoNmShSXui+ToUEpxcEfD/BuFvHD+wZ9oPwB
jyErFpozB0c0hMhWqcLVXve79puOtmfNmoF6VfXpa283iGcOKP4sdtakiEwBvkNFOe9IFSCUykFx
C86kZS1EnZu1gt8McfJSLSNW9tSQ9DV7ptDX7CFRJCiQPM3Ulfh29xAk4gFGC769wEhICkeU2VfF
79L77u1f+WMEhNC0SI6vLWih1OZrXv3bCdosQOUbzRcwEwDzWIRlCHiYLC34uECSnenye3mih9gY
Fx848NsbF91bfz3M3sU0XyYavSEZvR6bBDuj5ZGUqSMh5v7Ew+Zx5OaxfyBim1ZoYBP2VVEZSk0L
woBIb2Dn4Q3yGeRQ85zMUvLwIq1t/gf3YPCdGcgRoW+uxsqgbAb1RTfYSxq6cSrcfScVWjxy4DZ3
Ipo+Q2uaPjIK8p6oTyPHI12FvuBegVqJQkI2JR9TTSgHekGwF4mHBiLc39pcsRGtK4Uz46NZjdJi
O3lPLIfTshncRIKpazuquV9C0B8TUhG2knpUseHFFftCe5GiUGXKrUe7zf/FOoIAxtYI7oEkKxsn
xHBhfHC6UmGR77ZLZdes3uxz7QBpKzx6Lv3Z7tpm7ui1SK8cJU79ppz+ehdUvgIhv+Kmkw350KrQ
eUD5Yf3mjqdrcUkxzhM8lanm3IHHgI78HccB64oWXwVlbO7FCmptWqw3MI/21sJxXI4Zxdjemggo
WCHhB4+/Ez2bbkwmcJ8nxy/5lkrdI0YySDeLR4hbGtJgdKzTbPSEoxJYm+3iRWcW+rysakLdh0x4
CJ/SIuwc5hSYrLbyVXUTk/ABzwJvLenYr/676BNinpldvZ5V9cPcYSdixTycKUb7BWrI6cP6t2py
Cu50tQUWLi8v0hpwv1K9da+i13yIw/IuSZYPyyC5MMS0bVxnsLuUlKyTueZHBv68c9sOhC6jmHWb
rJiYJKD46lTLs/YrQSS5XNi3q7Y0HZql4K5mPRyxFm0+iWnLDJcNVGa0H6zWGQ88WbootFeNnOua
1aqzWilA0DtwSO222+PAKvudqLMvUhaA9KejBN0yGiYYiX9lprFLGWEIYMChGKVGPB50T0yOnbYO
vnyFPHWJGtWZX463JgU0/PJdg0HTnGhlKsVpNPbNGIMALXMfXL8aUEDmSQGJS88lG61SONVRp9in
uy0lBAXsGvCmTg9qOFCPQL22DboUNDFHBULnxb1YxPCe0JTk1PiQy9RhBNLSECz2o3UMHVbvnk4e
9FVdPgO5ZGI75hONUCc06CgGlQ0uHAhFqMV3EOtTbKvfD4TZUu2TB4RtMdoQx7sVkoqChfLAT9r0
M/DvafIxwC75E4pXa6ovcVeoCLc9Wg9TIekFsIJ8BrCbWVKxxQBAbD61febcEWwzyPmhNXEHqXga
Chh4SUf88SuFw3kuUS/yFowhQIxdyBMRQOpooTQavRHH8WXS1gux6pvEvHtWQjQeNrvgW7s8XcGI
zMLHtdY8qoL/2/UdblFFq0pted/BoSkVjABwlTWXhuIa4qB8G/BxBycYBp+jhGQdRzBgPSuH4JAx
yTL/3h3aLeioTUlgKgxbiWrJXeA2hq1W/x8BPj3mDzz95JIFSlhRLVwgHZAxWhosa24WPccDCLhW
mV+V753LpD5l8m3fTeV/HPpTyyg3HO4dUsW1WSH7uOxyxE+olf+nA3twMYbp6bQOUbWyzUDSpDos
o/giiwxfMtYXFfFCyYKNjvx0gztLPzKqdRSLnGKyxTeA8fKnH9eT4XoNw4+u2qm/GOcXIvSUTmle
DPVU5v7C7sw6GjH0+ss/pnsOvCW8UVb8O8Kwc9BQcaWl2AcHwrlrgUxY0IZ0bxTtLeaG2B7BkcI4
FgxN+UbJEx2tgQipdFYit046JGxE+ZPbn39TQ55Ou02xe8uYli4F2HiBunBs6g6UTIQwdh4IFVA/
EEsN0xBdPyto0EzktSvSo8lgf/D/Bm5YOQSvEFD4bBfBCbbkFrxEjpudCsSB5W7rKd9jHEOYXtYp
tIUTcGKn99bOPA9HdE+40CdAWOHQXLTqPd990X3tsFlYbLwylygFpd6VDY0yViOvC2MrAJQnpGXh
oCjEPtEVy2MYM4y9P0hNESXmTgTJrICwXFmcPkTo28q8hvoeYAFDCqRPSRujv0Wioi2VYWgQViXb
vJMgiq0RNbjlLhKlRgpEM+gzqarNon4yY8Kv4S+01XsNAvPli08DX/LHtdorxRbHS9Y3NcJ8bbL+
XkyllcVlaLQDL1X2SVjq7MwyugpMJG0uXfMw4FKMLbIRTll1RgxzU1FTwKvAHIRfr3nI1va/VplH
Q8HMx15p9Zk8BszyWI/r/z26tNXsaY+7j1880Kb7lkxqVHE9lJsNZBQ5MwAd/dUYeKWinQagsisE
gxs+EbGXsgLPyLE+x4BZEpGtVFk85ATx6AoD6yhz+Xvs/4KhNIdDfZe5SlXbO4uPBrX4xjXQKJCE
VCP3g/pl2AzzFiew+U2UMc9zetg+K2MOQuqTLtbsuFWsZBq8Cqr6bstrygPX1CJziub+7NVjs9RE
QVi2ZMqWITvDIt2EtVZpFUqDoTCD4rAFNjzM+Aj84XniTKz8ioMa20R/srOpuievgqOKWUGBKmRg
rnws3nDH2mPkLYD+ukSsp62ud9af844dn9a5CIrxsmU90pV3/rft+ep7Xd1F+eWUPVfGDULKM9Bm
PfOA2rddbSrAZ0EffC5fBLwVRhRYammN8vx4/Qxkywj/Hkwg70W0MopRBmTEHK/NV4ROetYrKDEG
GAdAoIp2crhvi/Uqzj/5J+JMOhrWEWjyjTUS3WxNArYxt2pcrr7UTuHyB8cWUhOTvUtYjSLR+SSc
jg4qrsBL7cOl6CwOGBPC3ls1j6W0jKVAm/1UBdYOiqN4JqpDeMtGKC3uSJy8O1aLoZrlr3d+s40w
Wi/dZ++cL5mSt9+PqGUFBnP7w8T8AQI7DopdruFTkqZx/kFLkJmpYYGVsuDwup2mWfDfr4QwC//r
7sdpC05AFNvJds4GOS34s3mswa03UE4l0qkQGm2pxv17pcBY4+youyhRZkiWwH83NAIZ908hLpKG
DkWq4lUhGmtqUyX0rhu9Aduc+Ce4iTNYaV2DFmGkc7SF8G0jSEp0iqte63AowMgOO0+6YnDl2geV
ojWJbRzMvxuUTn7qjzkBBrZwDAfc8s++wGDnHXTOnBzVhztmTjTUfDaqFD+mPMb8DOnOJrtnILxq
RPEP39BeRK/2B8J3xm0GRWnYYHC+RmxffyomwVg4p8fDSk45jyHXeiPzBgdEk42xjsKRFG2soIGb
Cz/E8uAioWlkZQPXiCObwjEJdsanq2y613vQ4ZeUkHbTgbhHu+2TVoD5zLiPmRL4gkTJ0H1vW+zB
TjSAN725ZfX2bKenXxWP9vTSLP7rOVec9FLzm1CvibeSuxQ8Mmy7wv7/OlsWdo6I2pUmyb5p/NbH
/YL84LHWp7aWky8e3S2Vr4aqWSYmZcW+lvqMXi+OJaiTcZA4X+Mb+rj3PcrZ98Y1TwAJoyr45t39
gvxgrq2POPmoY0ddHKLHTZwTtO5ZHySkzWoi+SABab1hVrbzw7knUbUjLY0M9eqEzEHoL4QigoZe
ZvUrLduWMD5UM/TadxEL7aGEMOcL0aEJ4T3zLMPKzJjRcSoSd5aG3Vl9sBPGK93kk6k1TPO7FbGw
8TMQ/qk1VrCh2hJ1utNJeo7iCmK0sf5yKwNw9Mjhduu3cIBd1TomY6jNPnxB/FN+BtqUsWgozElG
MX/S9Km1srseV6yFYKBdNxPNEOo/3lr0Vr+OyH5Qux6NugzYP8StMz/ToJ1VmjgkIVyD7tbqLRzV
luJQEtmLYw02bmislZqquO1Ik8HRFGr7bTkgrGwI/a8+EmwoR1W2Y3CA1cQCK+mzoMIdzDQsirwR
Pqv6JEdHW2ypQ/5Uc6JLC/009x3gUvcYSKH6/gtXdCSCr5P5yQpi4XJV5uPz7VVJObwAvzfFiKgU
xQkOc+iR7owbwiSSfyvNFFmSVruuFAFlOXiHRmbBiQqdG7qablzPfZ0PXbzsQlLuLP2zCjrsYRW4
3ltCLISmHeRWuRwMbInesx10c3wg1xQk/Q6/Ulj4Brf/HTmzqcbRo1J0AyCrxbpLFkJBjB9AVPXX
YBrmJ1yULs4iFcdmXl2GoXTatsJcGRtsUc1NYllC7nAu6UdZkIxs+AZ4G4pWvBCp0/W+XSzQUEnb
lsMW6NegN8Znec8e+w2vNBEOORYuLevrcxDRJjl6cGJgb+bDG83pUQgA9KEiBv7HxyRyGGqWfsb5
Cb2k7ktp2H0l6VqSnPnUtVkmLW5Mf0p+uU3hvPHFpg+2S49AJQhffPuh+gjPIcgVe4TR1WW9WlMq
of7xL/uaJwVsmRsn9DrjJxgyCyQ4hmIlou6BJFriAlhmWfWIn3+gCiLTg8lHuCoTOcJHohcnS7hq
K5126Jor1ZunoW4aPxVXzVMFh9aJcLeXOx/cJVPwGK6y1mWIKsqBk4X6iAQXrJ3kUlY/gJyOnhZR
OLe9uIN8ECuajrq2Xh/zFeCYoLO8cj+CYBaJKd9w0ZadV62BMCQhCpdN+hXu694pFyJfsoba2l49
dREQ8wliJzjFy+V5NByv0dqt1DJImPK0yO8rHJz4Mgo5DceXsKslfj2SwA34mii7ShRr54ESyYwF
icEdtbh1KDo8+7CW5Yk1D486Iu7uvCELP/mB8gtU9aKBx2OnLgNn6hRygxw1++dx2+AaGS7lSD3Q
2uc6t7CHC33Qchg6d1wgbONqrNiR2ydiGWXnF/EOAtt5XydW8WwxhIEXDorYUO7swKcicwQGTRKi
2BCDtKx2BOASpzoSqZOLMQDexGRzfzgGLKFJ2sVykturw8wsN/SvSfS5qN9ypHkp5r6S/EukCzQ3
hx6rlezxp66RvW+lOnvVsVjRgfOzx1G9PcGP1eyqW0ouYRYwkxqeObUa0pfFfqmCM+EIWWS+hTRk
xOIvVbOL+EpBYg6oCm7y95sIFb8YyzX3J0dNUGWdxkIjwCFex3Kf9NFh5JcbJ9rKKxHo75Z4Do/D
4bDXA5rl/cLHqIQkXPU93m/wdgqeqIu/7BV2GP8dlUZGhxPkUQiMHU239Ks+BMVbJt2pppUiVGHP
XoOif1pUZBO6KoTv1tG/eLJ5VnuV4nN7jTwJJC5+45p31mgyySGhiS1tMXgjagCLQ4YgtuFHWHHz
KnQXByKXH1/J9rM5R+3zcoJeSKAJuqkB0myu1NLIeHRiUtVzfevFOp+sOsMRrET0nDB/msGfYfWT
/2u5mtFnnOQX+psLyMzQV8wHv3JJKpisON6QoiuTB6VRQylN07iHW8XGhZpW4Jhhn8WCbpsvjSgM
E422VKWrgwL3I5JPDrxVFRLZG78CZlhtZnCarOOCViX8jCyAo81Ar8k6BKPe3m17qTeVOKU3Jlm7
WH2OU84BTi0EbPCU9V9L9pgrVcsi+QtAUn59mHXy3RtSYymZMNKms7JbMf9nyzLt/j/I2PEAiXaI
cZ5iDhqhxnth85c8MgEWplGFLK5BZ/i6Xw1ftkmmPB+6PGphDui35ycP6Hf2qjcn6fhw0agbzTen
3kBZ7/WIDk64uxIgmy3ceyfP6tj1TsZ3ftISvLUnGTGoa1oB8khBXqdnsJ6SEdGPrgyZToiO7wQM
1fuYAxSslTsjyyXfMh8PpBvVURUYOPmTExQ2iOyDDi6K7xpYxIdH7K3TWpUAsEz+2Rk6/xNMGnup
62YE554RWTyMEkr0RfJeHgvT9tyC2HNxxMCFXtUqVnjAKeM+w8bTkCaFadUO2GvtxTf69JZF83XI
iN68dI+HGKK+PhpU1a5jujPh9cbps02mnJSw2WWv8mmIOBs/7nmD4a6alCw8qqRGY9/1Nf8g0Jy6
XnSjgdaaVcmidrRYsgeJbz55WiI/vVAmotPjgVCaOTWFE+4BjHXrAfCumsLq6fRvFa/Cef2Qh9F4
7oC9hAZRTmq53pwihnqt33z5sAdhH9DKBDLNtgV75YkZwIm6IEDTToqE/3jfaiMZo4e1wX35hauj
V7SW1MOUhq1CIWh2vr/it46MeFp0hj32oGwR62mVACLbZ8AcX9Fhs0v10Ks0LrKtATCB9F7dYX9q
wY7N5dicmSjYwXPW08SJFp5N3ztE0z/mfXfntZOnA0W9ZJKnvAitIthL3ziKOp5uZHwW3VORgTjQ
N5KEhDbQ8y+/DfKAcofio7MN0mu+NVGQkbb+QgOjU9XZCejtx9l4ty1b67aUZXUEVZj+GztweN0K
KB4ghCf/4lodm1Rv24RrXIt1w2utVgvmirErtHGprNi5fot2cafDfm6NsSO1kuxcz1EIkLbqXExk
ucAblUyytqxBgwK/h0UAv3D648ZPQdM9NAlInDOGNENknNiWdnBt/hUr1v1oA0CN0L8zdviY4fnY
92nSnGNGwxOOraYhroD1jL1QeNfdxf6dC4rY90u2JAI6VtejrImq447nc0jruqguu+n4ERFAPMIa
b4iadsxWhn8JJ4s8KRhOetTx5HU0DMZAIkPkftjUV+IHUjhLu7Gn8VVo0ZNmemo/rjtFHRIbYWZC
mBtEUnpEZqfxxJJtf7ZyGaTlAiJwaig8vM4lZ+mp3cLU5Cqb0jBiMxqZxDGsOVyKCtecNhMqqBHq
KSCwYRdhN7APybQAlqMgnJZb7+HwEL+NZlfG0ZO+Wd5F4gPPjyy7PoQ3yeoRvfvjXeBzbin4tRaV
IHKWY5haQzdW1wDqbMBqCclfKf415VMYAnX9+R9MBs1MESi0vxF8qeSZqnTQQGAvvAXyn7RJX4O5
pDWb1x8paiVCa3VRz6/rLjHfAGKA6Slyo7P0PDq7Srw11EBFDfoVXSHsSTvzcIg+4qGc1khWjRi2
CzuC7KMxd7tCfhDPWGE/Uvs3jujS2g7jJQJ2PN1bMQk2BlVyOTyE2C2J3qOH5trtyRtQWEMKtine
L79BK/BjbdB4DCE/RtAeUGTC8Bjl+t+IcHauDowl4ueQHADHcX3mWux224DBDdwyhHTNQIEAvYJe
RU6HbO8ZknXCn67DnAFQBKiaystTsJNmsgcVkuLHe7YXVsZH8nWBKqKLonR5lKa8yN00b6x2Z5XZ
AeLxrePHuw9Cp/hRzGVZnCgCHgS6+huZuMi83qBKIHmIKwUzAeYBdbXjQczaYC3agcIR6Dl1Mc+v
Bf00PZrO8SihYDfbVfH6yVToFkIpW4a43azrCGswLAdEeY1CseWYJv33pu7s9A+AVm7H6t9IHEeI
WHN3yu+KrZU/dBZ0y73d9Rvw12sEVErDZvOfEQzhYEtMkWfltuYEOWqjco1NK8TjwjqIRisFgoYS
G5kI2pymPpYli+O1m7bmDLf1zDfCiPNf4hvkSlcdpGHGWPLI+RqKs1Yh526FGDl2tP24LwvJLcux
eihGgchWHpRdD66oMfhdiYZ75KLKM9P1zCJD9p+k+VFWNwtIynl9QStNHDHHB+9AboNq7cXEhD8o
YhEYV5VHCstsNxGVew94wLhhax1Xlx+usgJ2a5Ksvlufd5+IFStVB5zgjmiKQL7IWzMwcrTgzpXN
FVEHEb3vzYPXp1FeS+9oYRQgy0PIBnKw+6FT2GCb0YY/mCdOROXIUpZHrGLe5tAberTt680KVoKT
QuPvDfWCaUvf6D+wXHvYEAQVAN7czDwKA9CZGCIw/PcEXIBfr3L2dpbcUU5IPS7JxRAyIGDtE89+
5zbMnhX+ibCsacZ5fMyLAiyh+oYZdin29GeRcyeKqkg7fmjlYWBT1xk6onZHTG+prT6AGYnUPddw
46YPkolvPZme8he7H14oZDIePPtwZyua0vrbCyRzx7ZaTWaBo+zwnpjBLG2HD02V/MHSpZt7TmOH
bqDpP3Sam9m8BqgOCWDZN87Y47ebw2PWwdOYanyr2XGsZYoBkx506+fAn35HU/7vxdm1lmVwR18D
ti8unWLZD9D8yVaBCGiidaTc2Q2HbZXkukn+a6mGDkjWW3YN6FwlesyWu348kBZy9K1t+az5ZkOT
crjPJEOTAZRyjMzXxU8+iLyL6rdSuojoC4/aok9DUr+diCiw8bweWwFYd47wBi4ty8Kd5Cpajg0a
kBP1nbeE01dDZDuGc+Psv0SZurfAjqmxytFt+VSkXEASD14K9D/43EFf0gEs4vzDAhHC4ebJ1JzW
+PyIiLnBuvkEkg1zaaB08pfp/CSYu/v673iKeqqau1mH0bFOLsMfHphvwddLg2uI3N/YijUOJsJl
VeEl/ezduCaXQXNFWpSW/zIbbRBUgdqjBQT70v3Az0wL67WiUGBwFHHoRnqkZXudT46CJmcj2ia9
aCGCIsEPUXLopSdilC6ZZXHMF53WzLeFzS+7iXu9gNQDWRUgGX89GxgCvkseItMXw2LPLd5Hk1db
nJuhi5HLM4oyDPlFkfBiYix7rWYJ4LvtRGa+rv5cTZBtDDEh5sOp8EqhU++RP+8UiLGuZstjO9nk
fjVVjPS95Veqy+bfMJmPM/gkskNWTXXmqSVugAd8yFtQ6NtIEAFl5j/GTl31wldnzp6XAkcvYwRb
a4blXkWEWfdmUT+j2hv4pNsnURhiD6Hqd79CbglmgnXJf19AHE/wZF6GqfwKWA1Ljcgs27jkvhsE
wvgDZ675R0x1/aovHYna+EBm+1YWNc1CMAe1xbgD4/LvjInS+d3LX3nGbu8ALgC1i1CDUgmobDYh
lMRIudnZJeYpoLewZYqio97H12gJ4Lxh0h3Exnqmn/AN+2nDmQZ6fEtIccVJBdvS4+3+zLWk6j2D
GFG3t28quUZgGhTL1n0lQuew/KlN1eG/D64GkSfvzrVQLcts6iWgaDe7WJTKA9jRixi081LESR0m
H9YEOQUeOXwghfZ4eS9bhq33RugghLqgPh/+8g/7KL3ZORxjgtVXcR+ZQXJTP5UpCGvWXEQtzbEq
BZwQq/v9doSV4YVmrqkgyYKtzCqIJdaAPcIUXYIH/8SakhQpI+jYIPTVLFhTE+wF8MRPY9gCbkE4
go67gUyJmc4epHmgxzI4zmGEcF2QQ6YrrTsz1BVGtsPo1wl54DM8n6NBBVjlaIJhnG5fiu/iNaBS
c7Jrz8OCOBfk6DnRXIg3jGXEL0mTozgG1YkBEfP736LwOgpQDCg5whPtlmtidjFdHGOtHofoMvxX
i1/jFPFkfBAw+h8FBALAfmLz7E/hLy9BdVY+e7enOhoADG+Y2D+c6+WfLC6rlEe1zPBa9caStfjI
xqnxCKlxAh05f3qdYcJj90+YCzcNS912mMq9R7+GAbZTIN3HaNx79GClIXc3G9u7TCOdOG3qdrJE
H0udLlyXc41razMDCqJCf2ctFYiF6WVNQzWHug4Uno5nNy6D14mdJkCfORLwLDOTt5h5E9TLo2Pf
O7Ab3NaoSy7tWfQii3mceSNEonq/+ZgsGVlOfrr63g40ynw2E6VC82Hy9shp72/NgB2Kct3vskL0
nH7HUX4UYGetqWdPxL06bMaVpbQJPoRO+HpmjDcQlKtOCefbEMYKDv4MAOzCoHqRn+hsIvpVX6Tc
60kMPOC4gL9ORGFzsZZkXM3VHYACc8Kx/o1w5f3l63pkoZYI1rPy1iv1Bi56wGwoozZ+EM4UAOAR
mFrgK9ta1/FS/MN3ekGv9YGzPUt6t1lNJ+woClb4PwNejTkM42J3DPWe1P02f4grmniEVI13dYDT
f3Zc5jSFsi3ijafzfxmDPqtT2du+wsdzcU+wUU9/iWVw7uB5p07U8MmJFE3uJMIti7ZIkFB3OoxE
uyA5yKeUtfJLLzzLo+QzdFLJe4/jTUDX/i8pf26UXN6ymjIc4tEfwnZ7MfSn7FplfZ02sN86+iKN
Nq7EiCWxVKBqAaL35zmUJBedjf/NHpiJ2bzdQVfip/5bxYOa0LqkhgooKiXRW4pFql8PRKeSRMQa
hcuxLZhGfarEjt6+cYW5UD45Zkx9UOl9VcI5GD1B3M9GlKLyFNHC8dmKEBYPdqfiNR11XtN+udKc
g/1VlH80ceLGMMxA38HCiTvuwrlWx2BGEi67kUYvzp04p+RVcXM+1X0ErUzDYqwR5F/ez3FqeXbd
/qEiBCHloajctgOPZFSKiLW1Uv6FYp8fBvut9ga2V2Pz2ZNq5NDT6T8y/n9pzJ+I49SQk5omb1Cr
2k3ULtfonohtqnmrjuEbz4KxJ5d9QbwXugsZn+G8MmFjoNmvvx9iyIdrrK3KZ8zFIrDhHtFmDyfD
O6hv3NhyAH4/ckHdaIeoHBgcGdt6ZLXxXf3JMY1ZC2r/U4GT/zbz9r2qx2Ze1r2H2mNalCb3+xsu
s/STaB2ktgfYQ6GRB8OVOiVd5xPl20hKKcyUfLTzIbGAxl0YCv22QMXOotOrbKqrMi5Dshqtr8cQ
OsU1qWuGXYKRqoghdhFGLJHiFT5S0DRQsBSA5kunRnqa0TLcovVsE1KgJjxCCtdtqGjyccC++zFd
UcgBA4mT04VGPjEGZd3RxJiaMer1mEtneWCttHQGOhQCfCYSgzzTppJnwsSWVdUA67e+FXR+pSEW
Gm9y27yXUtotV9gJ3XeqROkkSeYU1Nt2XgtSWheRUX3/hZpRCxlpjH1DoNH3dkjIcFpvsAxd3F0i
KCxUrXojzOMNJTmvgISKWQxL+XhDSdUWzA+AoYD0MCTiaBFyxwDD2iGP/jEn63+CZqqs6+lVxBs3
4y2RUAItASTyB9WQeHcx5p/HRKbyoGPHA2Eu+yH6pix347myYVKurdg0t9xZqoOmanEQOcmHVawT
W6uMLTzlxxRHcWaSYNkIBfs0jtnfORhAXziFtRa5kKwIY8zoWk0x2bCReLlOHtYcoFgnkTI9G8x0
nLt7ltIr9nEvWY/laZYrUhPd7r0Z7qcQfI0pxVzcOsWUEZ93aiabPnunIXdKUguzWErErZlXPFtR
R19xrscmKnePHfkSTqFXT5etqdskh7brflogRUHQ/0JKLHw2kjfNFvPilqALXdLnf2YEk9Dmf8UQ
mbyDDfndsY566Lx3+EBOh062q1FYTl7v9uWWO54qM0MN1gJm4cknWZEpy5HMQvUZTns8ZonvNCZV
dWtHWbMO9Tc0ed23uDSllTowHgA4RBNyNbA3upk7kxLAPXEnT8Jasz7+yLGwZDWoysNsOnZgH44j
3/63xQRaSsJsxMNsMwXvBdmrv7WkH8c6PFU0LVEaMMFqwFqkEdMj+qOh3JYwUCLNRTH5y/0l66Fj
9TKcEPJn8zqO+D5+LQv6tsKq1Jus5rpz6h+V6JZMfy5fAeksDDtGc+lxCRslZLWt9ONJebpztUi0
JJ9/KSFm1/yr1axID1bKPo8UeVyMQoEV+0blvWxxg+XDvS8+KIRsRW6L1KmwZD/l/e1cAbjO7oGX
6JmLlWzHB4z/HMV8JxxjBUL7jSHr9bGa5Oe3j/VkDgCW0/zYPzbqKTX6ShH68pIlZIxNEbPwB4DA
8zKsogB0Pbb0ktlehC2domLUM2CR7fd6SoBSC8Obw0RX7fPFnCN+ZUc+ukUYltHWu9hzdsHBlKeX
mg8DHAuYA+Trff6+aQL/BDTMZcuQ8n3dMadJXpASr0sBw4mOBXgzAnhr04KwV2gms73J5MnQanQx
+p3OYhcWLxRDM//uSXtZvLy7whNULbtqtzkYNiOBMqS/pQ3O1pKTNlcNNOD69LDdaI8Qq56MtTwo
3IjHDZ5Wr/Kfvu8IL4uh+gjuZ9SzMvktsug4HbaghJAJSLvoLCEAlmViVjthGloh38OQ/4DaHe0+
a33GBGPL2xifH5sb/8FKJVWMSMwkOCEob7uEGWYU2Ylhea2Xv4Z93E56pj6sy1adu1U9DQwvB0Zt
av+kSf0y8GjBqygWEcORQfzJ8h0XgoapezUXRa7pPjC+FqknQwyRbiOYamt0DzaHwsnXmJJvMAQC
9WYBiDorH64CRYbHE/BgSYOIKDj1vLcfBYM4uDocvl/Uhrq9oHr+xnSYYW9djkmNeK2xDnYHmysd
MwQ2UuDqN8h3DjH+QtDATwCFn1sWMpLAJeqwJ6y+JVGXE6y1OZae2910aOZz2WA2Q39ULzLGtdPE
v11yenZf+/H9BHbkj0QECJiAJ2kMR0mgV6dCCFLIp1kG9sQ5XOE6FYpQvCDwYSygu+oEwqIOkEO0
GcIQ6R5zclbNY4H6Khb/VHx2lciRNPB6NKc+FaazsVSqBcFc+Wxu6WEaJ7XViZSaj1ISbn88rgoC
uALfJW/RkZlEIAxjXTbvhqGtwIB9xEnUiyLp71ftT9MvNhTmZZT3rYdZL9VrtiCZJn8SnaCXTwJD
rASQLVwIh1P5/4cSXxYl9vkIF1lmkNKm3wF3z765fSzE2Ea19jgkL8f/oesXOd0SOozo6SmnXn+O
r1DelFGUR2Mmgn2rv+lH2i82DfCxBNS8leZT+wBTy3h5OrJcOfaUsqeMCMryM/JiKcY4NDQ/wjei
xGfAN+7QsLLLBgxFeGlMs/krcwtPuk8cslLRC+mEdrukA9M0ZI+v3cnLl7BpZRLdMoyPrgWQ33ba
fMEgqsv7VMqb9TYv/o1/EndwkyPDgaTIdPIj+b1eXTLD8h3FHXkI7XriorbXa3NpbP4eZEOLov1P
9AvdHpFp+w4u9LmlNVX0VF/oZ28g+EPBgf09XDr+/OYx/mRXGBsNy0ktPtWHeNQcVZ/9WSheEODl
2VEP0EN5r7PRCPtV3dKtUIJZLOR8GYjowTnDR14xy9lLSCVj3dh/mv7k+ylWmWp268h65Mj2mkNQ
+u9f/taQQTaztEnfVadV04YIdEm74QloSG/mRgrZSUILkzSDrMuPwn2i+QehGjvuB5EVarWxPmnV
r1mYeZzSP94s2GFJ9E8mK3lQ1yjUoIRtmGffy+vWnHEtZYFZ05qhUFhRieHKesuhXaHOPBM59VME
NNZcShQS0YieDnuRvu7y9MRSkZmRyiRxPSsgrkMNUobYTAeL0QQYMf3JHU/bqsifoSzE0WzxASX7
L9g7tIwz3xZ5j1xcHC+W8lm8nk50Hvk55joaEQ0Bws/0Kp4MVKBdWRM6RunOiFsUfb6l2HMSvt7H
eo+aW2qABSolTXJNRMt7Yn/rEk3fvH/fzXdwAMQfnDDkkwySp+3/xiLJe7vFEDesshwKxZ+OOu8F
Nk8mkn6oluQMS3fnqPKmIPAoxI9T9b7adzWcWFH2LQa5AggkcSyXGyhrtXF+7rlkRAWFsV11dMY8
SKrkqNTh8E9MGGB2hTpo25j9QvEa7krO29n03kfUmfQJ6ahO34HWQiXenvhoAf/DGYWpI6HsCibW
yepojaWyjMeW22AoTYCrghhemfPxBUE6LMadZSSsUy+sF3pJaYwXfwBfEFMceBYo1Dk8bmO0VLfM
jeGWUAR+zYrP3qyxflmYBMiLyGGQZxfF9IoKhJOenLOFSRcAVszdVPjNr7PipyWqWxi/kN4Cr9TM
vYOKRDkMYLOwaSL0UfCsVqh5BLtV4b/UQLcqUOsPN4o77mN/nyLc8Kgf4zEQZUS369riFZCHhIBN
657MShcaiK6WQfP28zB/7FzS8AI9gFgYUGXtXuE0u4UboHXQxgum8fmHt8gv/7c1mrJYZ8BmApw4
DL5hr9GNt8wB5n0M6QSEl+QqDwuj39u4MouKmkFek8qycxPeTRAzFTmXNG9yG9u9JObWSp7MW3SK
V4wfNaSbFQZ4rEWaFTl+Teu9JEFbTMN1Rsyn6WL2daQFoEuJgh6/y5slE3Fm1TmJnDm3q1/LEUpq
Rd9SpqsJaYaru+NKBnXofDMW8XIUGKYMZKvgRrYWYua0i60Foox25GQ0ViFnhMGQFfNhLJ/rj7Qf
vlgmxcBLyuKrcflqxPor9hxXnPwFHXref0Agou+6PFhBfji7025Arl7lzXh4XgDGjOqzdl7PKFtX
CT54FBDzRnv99vHD+0f1Jn05X4nP3OQgeuez6GHd6SSbJBSKECEro7VTg7RfOPIB187LGOTDtWOO
zF+TDfTYdqr6jVLRa7zkWULBGL6v5LkVfpdQfgxzNxLkACaIZ4zevNnBjeNVPdL9DM3aFgsSopFt
U8DReg01BOEPp6xP02OQfGq/lFbqKJhmlhmLuDZLim2wjugk5uLHgAFCNGc8hmQhcysRzGqGmBNx
GBI/aAQaSV4nzmn2elkj0YnguKtyZerd3JXS1iJrKU7UP9z9u5FX8HSw1QvxdJcbE1m3We7LBpr2
d57P34kVkyKcR9ZPCEi8rm8mJ3UXzKp8mg5AiKkNYm9/4VwxM6nRK6x8RXgDpXxn907K/gJoaKMr
NxlaAJ08o/46Lf5YmGksONitPU8x+n5Fn6MHBPLqapCQzwahKMfLpgNwVL59SrL39GU8k4/+MMsl
VbQbzAXOUHby8/6AxEfo4nSJoRfpIi+Gzwt0VMSuQzrA49ScNMUR8MqAMrBTTTIKCPxhRNx83Smt
WMXGSmWOarhlWADc65RIbORxyStCH3eoGMQnyw94pA+3vicWESrrcz4qQxW8RUynpVfBt2qDa6ek
4N2eTmtB3++X8piuKsCJVbBaHuWm/U8ivdEX1TaxhbCF4WnWtP6UBNgjDUimmFB3TI3DU9lTV6GK
Xw3Ew0gbXVIloCy1Dp6e6oNATLqccEU0rhQDcHxb3G+NSp62dQ9L4tTspoc+kio0aJp+cESdtjxB
YzFUCGM0jbhMVpZzjaWuLribTrAdfrefPDEMcRRtj2nOSMlsHp2Woo4Y8xWA5hxX+imcgnKql7K6
LXUEVyk6u72QTe8ZnBOFEEHuRGgJXF6uieUQqpd6o0ax6DC/RsqUwgd0mRBOupZC0yO234CxgmTL
kBquZSn3if/9N9zggLhF6d3Fo6GuIukO0P3cBgXZvNMRI2BMhwMmTJc1pL/hQvbs9KCIfwZJPfIO
8SE+hVvbrqmJHug7N+dZBwZGT9aIJxws4TSSej72uyiegAERIE+EdYMP3BbwG+3rrs28PLNUptdi
Qpl5AQEF+W+ecUyCVpbpHiNpXE3iTPSpF06HrntoSdLJqANVnpJF06qvhPPJgmExFH9d2EoBB4VE
HD/XaI6AZBAk5lPZhBSITLuNfILGRSzgyYm7upoPu3rSu/Vezcaa66JRjyW2zmwTp5wN7kpmddEy
HNtUyg2oApglsFf3335zRYTCj43Inb+OyLhw2GG8H5dPOrJwBBJbSxY5idnOqeADRRo9xKcefSOh
CpPYDcWdStlaEDFXcPSbzH6OBSbEdcS7LUKEgsIjT5n1UEr0BKlnJoYbXxjX161bQoftUfkR0mdE
gGM7KSyBVXe9Pvy0gqA8suuI4heYUNbm+2CNcl+1/r/LQDut5yHqf9b+Er/DtO6XjFiUX14Ocd1J
Epgrac2cMV/rtB2vk3jfkPatysNEKT+Gm/k40CIAcx6wBiNLYI1BxCf5atWxRpdj+QkKNM6WRRru
EEE6LTCXEctt0sdlnvAgDjHTDpZmm9QwSToeYDe2bmShNZmWNqAniSt46/+hrCEv6cEaf61dPlq3
XSOMMlhDbVl9xlDimMAs5qJagHdjf3JwdU0rdNTtx+ys0abAWAaalRRjO0YrJpTamFdVCJ7rtw/R
aPUToLn6MnUUFgGBZwkUePPUqju0tao0jfmz3CHrDzobGN7jUVzjg5CABtMluWE3LmWNzKlwn+Jx
/wvbyk4m+Ndw9sw5A4SqXkGpM85WOMbK7eyh9ZCE3HR+jwdd54PbTeSJr2GapO071OMiNWFjHb/r
TbhNzfu2j8YoTx3Jh0+KEbgPh9FVzKS+3sYIEShxT189K+Hlgzprs2gOEe0zdvivF16dbfZOA6aj
U0giQWIWU4S2U57Z4mbGPP0gn/XUVZ40xpfEbQr8sTJ971TZGF/T7IO3WAwhresDpwDhHXgEDus0
ynWDiuxpJaWcAMuJLn78mbc+avoHfGePGUuYdG4YTfJ4X+fkUeO0qjgQUwjRTJ0yVKs1VXEsVFLo
syBYyJSD7nykSWpS1djxyD5GgnHL7xwjqXSsEpH7BKyt1JJy1RUVARB4snWOceEccLeyDzv6ibJz
V0+ul9HTXFwV6UqUnLEx4BnSIWdybdobAq/uqKJDHwNS1xOsGzZYiidAAgoBAgVJCzZHprEMnxWr
FOKE2zQiF2HYpujuB7B/F8pQyC0Paxn+e4/D19ioTEWEI8JIfgTYK/2GV22tS+jPCyTWyhSVFjlk
5tVzxtygYo602x0qHQgK7LppdJgqb/EX4Fvg+G6DGN9D4A9/kP70VWJbxwwkykNFBsCXLlcIxHIw
Ygg4lrEMJFNdEtnWqw5YKo1Hyf1r5I2rgIYG9ZuOTJeEMBBa1gDJEXAsW4QMEDd6xuT0/Oek8J3G
mTHjJZVO2RJm8nTnxlbhxQJMVIDiyjN4EtdKTR6SD0FrcY9GKatF3wqu91ilyvBkIMfndfQTJLgX
eU+INwcpr379N/ivAQhohwhUhJ8NZnZ/GJJ0l3O1di7o+5lLqemxKWF9oNvCkddTrdH4TSwSH/VK
XSrvoW4yQ4CyYZZeqSqXBVsac+M9Jc/yehnNn0HJtjdo4gAO6vLKwiN/7GBj2ZuX67apTEqMHhkJ
oK/lqMqLn5VCCb2fqyKjRMkLNpkKCB2DMHlDRzJGoQTm6YM4p0tEwJ0Ujt4uy7l4DE1RI3e5Uo4f
GDdABhQoD13VtrX6JA6DXnvk0hurlzPg7JVUhnLSVVhJTNfgwMn7nQlRZB6AKQeEFB2zU2b2mgXO
bYjNRXBdHsWEfU9LwCHmnFjbPtOLq1Chlb+4Mob/VNt8OEB0l9ycboB9hrwHrie1LcGVCqPPJGWO
6IoLZ0ql9C+FXY83PY8KbTj+9MlXZl9bOOjwu4/MAd5zhm8LRCIPm05WqQprvgqSPsVr2UsNj4lH
kFqnVCajrgwmr4k4rm1zfCmeQZY07oDvIaPxo5Jej4fn87827H7PBEQN8lDUOvTM4Bvea4MPu0ld
p9JlTeecR/v4f55p3hIjOQ+NPBE6bAZ63jRJzFvS/xn8JQnO+Hqz+qXR940O0TgpYsSi9jnguXbR
JvSfXiKe7umASkuogPMxSbr8rQCKAXH9oMlLDQN4AyEIZELtVTO7Wp8tbE4QgaVo3E+rM88RfVTO
2l1IzZKLYhpBuorf3ocfGC+jTBMiwkWxQjz9LilnIfDYtOrCu0LWb6cTGsnDiHE08fXXiJpF1zRU
y3J6onT4D3e5McQeIdGhb//nOmt6xB+dIdTpbGbPnqgPmoJLQNVivmRnFzcuEq8yiXJMkXJyhKYh
NJeFMFEhSjkQ7R71fqQaDxaAg9S6ry+8zlArKoodMeogiubr660BLogUj0ZIMb1hmTDlJheIt9WB
1TLKOQvhspcHnh/98+SMmCpHHxjm0AxEltFDCgmKcbqFmgUUKpKEhQuPTsCTN/QyXbne0KjguQ/i
0rRpBibwd6pZHBS/7X25Vkde2M0pPk3Lnct0MsART0+jrV2gHpJdx9dVv4ZQF1g9/CkCQ0deepHg
Um5naNm13Scp41dxfwmby24ppjBfDhDk8sury9arzTjRfafWlrKYrdemFMqmnY4BfuWXLW/tJJP3
7AOjGg2CyHrSg9Bsj0EluKJI3e4hu2eHzzlmTbk3liHE06BmXpcJHG6wrbP1wdaCMfra2poxyu4n
ypH8COubJGO0RdFgiWmsAJ7XRjWQoEU+qcFQnpe9geHZPuXsozz+p2XlNEelNtoKkq/YynXlNhpU
2GcjVEh5/bpD+km4Y47cl/pwgfHIz2jsLaRHbdgikuU86IYKKxPTAOMWcMA6eZs24ONcx0f8gaCj
vea9b+ftfvy1xI9YrmtsoSz30iu0bVFrZw82aUmpnrP7IrofjzDOX1VCdjR2RU/KEa/B4fzvjivf
Uf5Jys3oIDiYztJdEMnsRfJLquKqzgF9a9Sg/UYPvHEXv46yZhcDMiOpbTNTKb88G6Zz5PDPK9fV
6EW37U83GmPqtXyJA9vq1xbuvzhxEL7uzMlBh9/+m0UwvOx99u1hZx4Xj1AdTE0iasEih09kKAgo
leU+8jNxIKxMplGdbMFL6XahgHC+SuYVJihBkQGx+0rf7HXTA57J3prbXKI+eKQNd1k/RZcrRSTs
A+G9jrGnce4wQogX96T7kbXIbZ+A0rPTSldAJwP5+xYHdEPmMmis43aeV2Xtz9ccOHutyfB5DoKc
aCM8Iueppi1mdK0MuwZRyHiHcBn5S1U1bDSHImMtmvJKHhA1BH6NCmSP++GKLLrKD2kWoN5NfwkD
T21EM1EnRxXj47+DFCEtkpsNtAUWsG05ZM/f9F8SoETZ3UInhZORBSWJg52AJCdxx8zveJtKpCAu
RutRiQswP2PB0HYRxy9YldBoby7NhEmBWxqAzOclufIBCiJ7ilxaRBaJk9CqhYHgo/E5M3bC3w63
cegkFHTcA9YTdb2koeJgsSrJ3BThVMwU3WkecFPiQsanyt7D+PcBT6AzgNjoH89qL3BHtZ3HPy6l
aNZF83F7iCKziWK9EmIl2p3VP7vDwvFwlHYrtXxGRnEJ8KOx1gnphXrxc+OBaHKb2MN3RAt568Ln
ScLTwIpXyNBf9DbjJtt2w2FLfumbdq7S57m5y93rdmDCrrPqCWN16YLPc8IDYw7Kk7fomag/+jKq
K+fFXHjP3KHFIaXn61/Bf3kLWzwmdv0fdBMoZgwgWr5zUaY2IIQ3jmH8q4pkTokmJIScaFpnIjJN
XOAfftC/E8I9RAW9YoIWWNQkPbtSqpkEMnSZufvRazKNJlZuk9HdFkzCp3lpwwfcDRGbWMNl70eG
HT6fFlUP4aJxXhRgt5093mRoe7Km7Vy0T/2AxyDqFPNUIm5kXJ6akX5T/ZNU0SrC3DXAdXTWdNqP
a27T0/R0vEyaejWgQLbuTtWf6YGs82oO6H4qJR0GVwvLP+bgZYw5TwJ4LgcyhLJrrsmJlmiYP4BF
jgeSSCCnRHAsaBuVvR5QrRj8zmtRRwcrGENnM3vk0i45sI+Tv+btlWEsAsCDfhdoNOxXXgKY82Ed
WFH8Rk+lSPE0ETOZvG3pBDIM+0EsEbdLYNTd/kMNKwzM0QyGbAGus8N0TDCWRuXN0NCZqoB3V4Ou
0DlR8JfkvfnmP2l+5uhUsNMJLVWRpfGCq9UrAymdW+URKXCcYKarMDO05aoCnCTukxqgKy0iXWBq
5Dgu99fU6VnFmdb7IFQIiHMrjNcelmzc4ffQMb++fvzhClHu0iRLFtXl1S8Zps7CfrVq0kTFX/Xl
SyixRN++rhc5kBjuB/oxhuHrcS4YsuCfauN4FsOoz6lyqDDoL4IdhilJ/1Y6m1sgbEYuJp8JdReZ
zCuiyRQIP1ZQe3r1d67R3RN84fKW+IZ5cbTaHDF/Hi4cA/PzZcyCBb4EH6X9OTZAZkVmV6dNT0/T
bJIMheQYcnJUJeqwCctpOcXArBwy8iYmRFRjoT/8stB3vnwr/KozOQSmsrUDgxFFbBIGalAPdYaP
qOvJDplsv8tOWrlv7Q00BavOTR/gs5qFoUu6tRSgG7IRttFGGsZc8haTGR7E1M5p6964k3eqXsh5
7/n/C6xzaA4/v0m3BCTIGfuuzz/EI5J2y9yd2t9gWE1I0r3VNFHXzrs/BYdCT7N/1s+rVdwS0KvC
gEYKoBi9LExSTuTMaxJlgRjvjQRCR8DimBaJBP4twAMyDasZ0Js9utOX7W4caUbQCJ6nk33p8mjF
M9SWmRjEg336ZGQBXCmKk3edeSBlKWkvfmwuBPMRflpCTlP0P3pHho6TQhWYEbDlafUcigMWvlwJ
i2ADbqhjUneIlw13Z2JmE7XC7TWA5t3OEkNk9of2yRKDc29Pvm+og1Fsr+M9ZcA9hKpwGseZwrY+
LoOaUajWbTjhdr1yn09wDf1N+tt1Yzt6er6mMEhWizAUeGWu7tWIchIfGF/fqBrSWUhyqwrfuBTO
e0cdJ+1TV8s4qmVvwF+DBE/6GRHyACLzPkp9mjNPXepWVUaRdLvHGtywyvNS9yl5uFo0Y7nHFjbb
IqTJqCXxmce4KipN/Kwd6++WuNNnDcmo4yCQrwDJOM8RWY85CslWDu1zZzqQO6MPdy6mHWtCX4Dz
TXwucYFFkILx/tKgmMJpKQR9uDJFJhQ/CroEJl2YPHCvPrDqFK7u/RKp3l34BgFzP9h5ISfSOFei
//7mRL+3wspVgBZILrvOXnKmmTS2b5OmcGHrw2aFzX2Y7Mb9zVIHG7kFs9aQ4YMFX1FbRv0MqcIH
SqPx8R8L7aya06hHFoIlNHPqt90xnugAyp/9wELducvDykvdSrgh3941veLLObtZKmZWyGbZ2WZr
8ISyFNzjuUORGIPqiTuqwX6lpgqiS41dxQ3Tkp3ggXZwFF/ShQsaJH8ThaXhxcloD5JwiIkJg2kC
NeISXhghRR/DDB3f2HBY7N+XwqQbWDq0T9zejFdMneDM5cBILpFohGAh+Vc8mkRpfjn/4TUrti/s
NWwFi9GH0+80Oc9CSecJQRVhmRYyyrfSgRlwCtsrJpJO+X1buLAEWCtk1385GL3+vXoqVuPBwIbh
24O48zPOsv4IaGgsbgNr22907pJuMF8ROtWTvNevFBZrcLNtF2c0s+QyL7WujczyaTKgF50gmmFp
cpHvmEBhOIibcvbeLywdR7YQH+rS3DQ5J3inJyAenAROP9OUk/3Rv+p1IlYS9QzmB7rbrn6cKph7
avGGH2ALgZaI3GZLtZIUd4W6uxvD6ms0Deg5HhO+Gy/t2xJcVU6NrRDxyYkJfFGALrhpd2FrFK1x
wGA4AT6mXoHOAPOlSqvi3tvo3koXI7bOQcJ5H8hKP5Y6Q1Ccll3fxxjG7rTUZ/eJvnhppoqOI/a3
VVmkCVnxQRljOWsjsVbOCSwe+cZYcRTlT1bp0BnWNUaDTw70OvJ5HvA7P28iHJ+DxlCcSJEQj3RV
hCWAFZJ/TDCRdPHCSGICPn/jlni1WSEScPuFHcl8PfuK8OjN1fuFYR4KWSXmOvWjxM77vOqltEqn
oc22pF00wbhGI9+A3SLRYdh2FBBaOdi5VhbRGwTlSShEIyvI9suwIWYawqL1MvkeWCxbfvikd5OI
GV6kvlVGEtxisVsZoWhMj+HUR9nDejSXqTS7NSVwWHKdI/huFDRmbYervzrtTO1RgV9zvj35sVKi
e8xf9VWRIN3ZnfLr/p8xHk/OQVcF9rFoI78LaafmMR4XyOOLzYRJ43rKExqtVNQ41CfkFOlZTj8x
uhMVSKwnDa+OVcKS6VH7ALN5ooVK+suuDlgw9H9jaMwY6U95nNsmJKgs5dxXspClHel7/+00X4Rm
SvvoKwFCRK6o7pSwqwkLaGaLBOl12kWGsG/of2yLRPQTz83PSPV8fFiPqFV49ZpkoNKA68YrBDnf
staLKToeg1OHA/aKO0bfLPvQnQ0tiOZKjNRUpWMKDcV0ZaS3xkk4NqfoIw6PrqxSAoYaSGvQDuhh
WwzeU+40iDS/sraUIy4m/du7eJbYsadv9jsJjdcY2dPfqujxCDia7kfckWKvvPFRSIdu8jsC6pl7
qvimv36r8sS7B+OwpQv3/YxCzXiaTaa3zGZHr2yYd9E8PrRPn1zDHLi1xXOClW5wBvCQRUAYR/jB
6yxNDufp5VGdvo2t2agmY2eWPnaIeoMbM4UGd+4tnCBnVVn3mtf7Vm2IJLpVnNesgj35Mbs14OIa
5GPraUwtrdoROHHKDj9vE8O1gUn1wgJyou/su7o/n/7hRlKTz5/GgMRW2zb2LyJT7AHlkdhoe2GL
O8NCqNT+DWGZrmomSx+440fvia6Crxin7wtrtn0pSmX2tLnVFq+xJbNb75D8xYSATx1TqFw0P+hi
wPSgjuDzPGczDXGSBM3+awns2uDNCiCnQwsRUiBQnvcGcfMBldmjpWGk9FvzsDlfXjU5eVMy/4yz
LSK/o58lv1GmpI9qKBJ5BoLC/LbhcL9vZudNxSSbYF5SohKFoK96JPoAIMaBWm7RUyA0iuGX0g/v
4DYtfWc5qO4MfdC2kyY5PlpV3VrNr+JXEJD+AribtH3DrO+lwKK+/0axbpp0brSVkZfJJ6qOKR1/
CZJ2IJEOMUghVHLRKD2pmYLPJf+hJsZMqYjx7W1PKWtK9N/RL2cEDWmY6Sx7bqt81WeI70inlpDm
tVHrzb4P6CTb/3TNkY0T5SqDS2B8++csesyUwC3xUHphlCyJpeiJ/vb9hBBXCuwTha/5pT8ewKmD
/nSb3gPqXi/qslhWkGBu5lrb9wG75PVL69LwkNsQaBTZL16evWaOFiFGBPZHGN1KOYJZvKf1CD7C
T85CXkIhHHdw1k8mXb33tvqGKSI7Iifmf5lBAbIkvNQHjL8uh50PgrPG4H/0siJIgnqp0hEgacdO
QKtiwGAye7BblTEYTD9i54xGAkT+lLxzK7p+YyIevUe6sBBgwQL415OWqWSZkQ839Pdi3qeV4aC3
O0J/sqWd++o5r4Lzicz0KQsEHYqn8XSw6ZMlsFETYPB3dP/O9r3jTERQ5Dx4lOfMRmCNr1ShGh+z
edSXJ59ysEc5Z1+/jnbrk2mGILzh8485pSxQYdxDjDyiQCoWeQcGW9JfHH58ByXAciYRfqTSWrxm
w7NwY2F59/sK5FhOhmx66jqBGZ6pwe5BeB0LJr6k/RQg5AWtby+3pP4il1M0v4U3oOkFiJ12Sdbp
ZYZMAHIh3UyTNRF8mX6AMjuP4czqbQtqhkiEBsdb8GE8Qyabzndv4yOUTQFdqrpyH72zcb0nlNdE
HiZnDbUVTIeV748t2xekd6gp1HyYupA+8ZnF8brXRnWz8FLDQoVJuofpsHWaPKPIEM6J61d4Onm5
RGizpKCw2RNMOz27GtP7axfhtq0/qfpJ2khidB8d3g5nhvN9ZQlmk6ocZi0iHGV7gaMazSqsLRjm
scOkFrmI854FkviQ4AsrnRm2yGMOFZFry29YkrzcxA+qrWYNqxYgPbldqqbh+r/EKqR9Ntj0iVEY
EDrd/NEaJD9K4Fw/enhiNi/KonUo0zn0zw0efuN4dUDWtL45HN/LTASKakMs39JlC3js5TnQnn+T
TGxbs+RaUbhUN4moBXh6ewyqLvxCrBtmCZm4gDhVqYWkpfmhYMyburOeAXTbSgWLEyQUNrcdp5Fd
lV/9Qs3cWADbm/msNggV3BaQarUSFKefjcfjQXSMlm50Vo+yabE79EW4PftHWuFxuIZzqmzYxn5y
/t/35fXk2MnBTP7fOGY7IB9h+09mHc+TBg0FSg/j9Nu0WkiqhpM4zLDdmbX1X6D7DPRLZvkIJbhg
Ayt6DR9qgz4AsqIwrSc4jw+auLCa+6um7f0uTyJAAzAr5V3EiMnrXN9ORkZLTu0nBTxfiXVppoyO
/ejU1FuFCLaI4cpFNkrvx65BroV1XGcwe1+oAH3oKjnc8K7Rz9x2GQnx4e6HzhVAj/Qm2bHwncgF
E1UjiNvb3xtszVhc6M/AZdk80v93JWpa99iFHHHWscKA2dGeegiKNsTXhOg1XrLJ1FhREMrw2VlF
sHtmtugvwtwN0c/JUTkQFmcwCpQG/qn51EGU3vINTORnnjRcX8q1F1CVRx+aXA3QWUNf65b8t7Tt
A+/MVNL7X4RZi9BuG+dIzI9OGU3TahDaqm6g5kqrpVQ2bToIkZ/rVLOKyt4vJaYmousYVqRmZUMC
EUuaM6eH0YpNChRaYJI+4PZ4AEIrbyvaAYX9pKjEMoSXoEL/6p+j4sGssgBqlgGA3wShbwZ44zhc
2uWwgrejtlCwNgjAqxmVdtOTnjdJHsIXa5gHxKxVsBTs6RdUcUZ0O3NlJWsmy/rAt+9J6ynmc6IF
1ClOgFSygtwBkxpPdYiThv0B6pBN0O/faFw7U5bs2E6b4K93zBN0e9skdQcbK+GpCB3szx+6CUdD
WCAgBGwJKN79Xv/AhNHXEl0VNLyN40lD0UYQXl9eC2TpZrbnwW0qHoCDiHi7JQzgKqr9z4AUoW6S
LSUItF566KFZ2u/+UFKF00r38YUxvK4PQcKEjYM7g6+CObU66BCuFnmdKOZFUcWlQVPt5dx1Hfxn
1IkAERSTu8OlS4iPTSb5cFxWEFejAI3YlSRMeXuJ7BTqUCrnJRhSsAS61HoRzXAClKQseSY+6D/L
guAn5bg/bDhCXn0I67JZUecsu5xmd2YfAevJBjUnPFAohUoQL1i/Q2sx7hqwFifrPXMxe+/c8fvc
ZkWX/FcS4r1R76SnOCBS7yZBlgJ6UCWMEpqDgueraK1xoOq/9C9Ehg4V234VeUtSvIiFL6RTVpPP
YHApgEcCI9XegHy1yjwrVDXkf2ExN4HSZmB+uiS8P+xlX1LMtByglk9b/rMlBkZ3tWUTV+GxmuVj
NUl7nbVQcl1HOfnBA2uySod0Qb1XTKqPXgy52lJqWQkD8GIx1YS+7094rtS3LK81A2M3CnizLneL
LS8D30ZseGdTlP+LFVz1qJrJtDzzZ0Ksbf2ouB4d6OJxfCKHUJj80rk4kgYDRU86+rNWQ55jDzyt
Ht1h9xZmI3E51MctfzGgG7W8VpXTpSNw4m7PSRqo4uw3oJb8oOL3BQ7U7eIVv/vsM5ZlmjP64lDz
vAInpOgAg29cSdS4t2EVqKm9e+IVkJ6n+rJT+a+Txjq5yrWIJGmC6tHY7+2X6eY33Kl6FsGJmpk/
vUeyPxy7gvo74pIY+KsicCFPs2wnzeqxPsPDlA43a7nIETpZhY3I+0Kv5q9L8StugKbac/gpAiYL
WHdnhz5t6CLLRfzckO/akz3pRFRol427K1STCHWjfyZZpfK2UxAzWfXCUs00T1T5VjCh3fJt9GUS
ANjbYfEbB7SfeZyGaIrAom8GzlY1HdrsEzk5H6KtjUS5YyN4x8Uix8cRSqoF404wl8YFwtoSNGKN
qws3ISQHqTCSegGcyUSwhP84bAt8Gu42YGYB8F9NN4ezepRaOyo5g6DffXjFfHDRufCUY6/iBO0J
g94jOtPC1mkfE9Ml+LQcIwqqNpdnwCm0ChwwANG7EB3yYAOE04TxgUmCgJqijH/0NIdv+kVjISVe
fKPTsThWg7lGOqFdXKvW4E7BZ+lAgedLzcDUv/MTLQAjePgEC9RV1V1I8B2BBB6zZn6IWfOgeV2a
LyZfcvd1eZnPoEV5N1Uz3MBgpcxsazi8JZmoW1iVRYpGenCqG9fX9dA0lN+5O1O5LvsJOa48ZGhU
4uuFl6VtParkyVetbFgjfSlPa5PGab4nQCYI2UEYzQM3xnFCRphufuj/Ov0/ehO5OPvQvFsEbEBB
PqmWWxCB4lrKsg2iG4Qeu5pcwyNEtKW1ccm39AadHKgUIy6qVE4rvl9RGkCGVD8k4n431fujoRDD
sciK9kHbUlNw0vu0acbR2Iyy6XxDt5kHNnoaTYacIfsQyFINh7fDoRF3ZNlVAtQG3jkyz09ePGxK
ILUEe+5o36O7/hBvyTw4ZHtKXDVsZGjfcCuBpLlCvK1fbjN/gzVXdyl6/zpaa+KamvjxLJUGN9qO
1aK0Hn9SGgCHuJeUqDG2/h8183nt3uZUu3I4OJYbB5k2XSc6sxKGa82ehUY0KCkUf03EIGEtqKmt
YVg5BWXWhFzysJI/YvoUX41iD0Mj5Dy88fE6uSk/vngmWiD/SiFjmS88ZLyo6eUm2uBaV9uCVR41
m8eDbwD8VGgBN2Tg/E1LYRyxAIDAc1Kb8G8zD+JcSnP7ZLP8RI/eXhSx8UU9v9dDi77ijch42fTC
P2XrBEJcaq4QHcu9JD1OQVdmCl+MY7WSPqjytRfs3zfzDkWybuKrhf7OY7jlcSsC/AqffUP/YOt/
9DEEN4EYrPmWpXZ/PDZpNoLvoveOmHTvpCDX0HGH7oN1OyyQBUesRhAPG4TYIMs3N/ZlgINdZ/45
gLSOHklQEalB3VO5zCBqvhsafcRUQuleoceianP9z2v+WqFD/mSZCAQaGOlHv+jfPCv2nmVyCF79
cNS660V4S5je7LTonZ8rvJIq+aD4cXGyeJqBguPjgbGRP7mDCK7BzFkuwvxR0K2OItF1j0rwQF2c
ESulisx9SdL+o7PjPTnkuyLp4bdeN73xsDIrv/vjm1SWOdSKEDpVSAZGB1kYIFSMd4OxaJ5wEPbg
dSr2l1IJYFcDOY4QbkMMevBWK6EXjdvqxb3aqEklW3J1DyjtYUDFXjbx6O6HFBNPBwAdZkfrEAu7
xvBnKOIPxqNAgfD22e7DQV26aRoFwUhHnyF99gZGgtFNVDQwjajA8juwfGRjkDI+REGFhapxjZ1w
q80VD7s02Fyl8ZkfSmTuAcKbryoGGV0njR4SjrSeW38SoOBVJN7mbv0bO3BcQCzTeoCC1Dr71Xx6
b+j5wa3mblGtW4VZlRQVAibkH1oXowPCnFrKDIx/qfLWAcyu4HEHswycLghHWEu8ZcFsvaQB7UMU
H8YymeZSI9MnPkDm+BYmisjbPioCwtxtGeNjRDeGYh5oDoZOGMkc/F1FHBFUb860sN0KNgNKblZQ
Z3Eulu0u0f4YWvpyqFz5RdyuhH0ENI1DB6IwJsQGq++HN3wQsZe5rq0pf1auiG7bDcuWtt57v2RQ
1G13NrWhaFvvUZkUH6xlT6YBQv/IR8FqDJUmznigGbULkkZT2X8J86J37kqAeQFxtT5tXH2GWI5q
JjC3B9+qnoTE1gGgMIeixRjYIewdYbNeniHgWACVrPhzD4ZbSvOJ0h3bjhmCK7Kw2m8DMJ3tuLT3
VSU0LOHXgmyeMNz3vD7BeTsZ8xsbfETckFpkMyq2QcLcnRb+N6hURCiO81qZeNPYVTKz9Qz+K9iD
pYnVjsoD69ipSkSKmGyqO4eMiOO0ntCuZ6keXFfwmCqynDjsVA3etYQOseYBKGS+5VtsNx8qqjbp
GzcyKIXAV04FmIJOBJTl2+daytvNPzewn2FBE1/3tYqWotL+qXYQ6Oiv/OmTl03AhktHAwVOS+ay
QYc5b0i0xdvrw4c1/3iWaEppKcA/nEo4Hfm9OCgsG3SadJvXtx32UuCN+3nHURVeaVqJNDaDIvHE
r8GnelL2Ie/8j05GuQsCl1afOhJHL6nqbG1DeHZtGnvCRnmQlZqn3ZtB0cq+HZ0oWPTZjmz1ZIN8
1eG6bhMgkr2vpwyM3rCQp7CtNWpLMi9F8cihPbFmJHyK74lp7Br7+QT7dScwO7VGvM2NX8divgm4
ujRK9scveElHn0AnFs08az9UK+43HQOsdefWT52GrxUwcgLPk1X8lvELo5eXX4TZDhsT9aRSs1T/
+M8RRqSfjAxWHVWVZBeNvfi2GR8fpgaVB/66Jzvi5RAVbA4RHZSjSIYihiuc56q5zYNjWXtYAEPA
KGELGGd1lAEkJ42/1tiWeazmoBAb6IePJeJTMa8IhIbAgMaGNRfC/T6FlZ3dla4wT6zNSAeJloq6
G13O30jOIM3bRGF9yOX1tlN3yNQ8Y2FTJe2JmF/oj5R5F8pKYTcm9uCbq5/Qg7Xq+wgy1SuyxvN1
W6u5yftb4y7bQoH6Q8iSDsG0IjgYc8pZiG8+Gne6y7ek3riPmKWuZJbi2JnCBC+Yaw8rLfGhtRBg
dJSrI5vYccn6B/mKOhctJ4joRBRx/AagumXccGhOOzaAu1+XeiBUjWifhlZCsHD8BUgxZBAucvRp
ae72DvWDjBruentrt2W2q7M9xnRTdN9KjX7OVNRHWpsMwZE9HRG03GZvBFyaANJlj2uF9v23Owx3
BmndgmCXyCHprIvOElnVLuCvaI9yN4iBazLIyh1McMr/o+YT5fS0iXSuno89ukYmHcuAsgUDl+BB
9SPIYHhKbqCHvQqHiTR6WFAra6JCD4yh7SWtRO74t+pFPo/wCUM0Jnq/vBptcdlNuNXAtlYyfdk5
T+d19Br+RFCZ+BNaocQtOArNjGJ8StbnO6IaLhpdUikZ5atKDtFyXdmOSmm6ltqp3c0ytzPkwX7e
2KPa9+Swr5p/nO72Wx2tsd5xRX44nZILPJ95e6agby4O6/crFDcQmramDxNrX63UWYYc/sfVjhxa
Bi0Q0CXDL+Xz+n3C0afTvTLx4bgelBSN1NGF0OUz5OCWl+kzcHeK+lQjK0x+hq+Suhaep4Gkplpq
CUjuGnhzKcQaCjcUWBa9Xaeon1BWhbJBtXHY18RRCscH+FLF8TWJCnUrJg91+UgEefOddmZ3Tjis
kerO3UVMM8spAGTtRXYchY7btiObQq5gIrhpXK4bEJkgih7C/asI6/n049Ss3BpgGT0+hOFzQUCb
glllQr/UXMEzt6Z7EyyfKVx1EkpU5QQjt287jmWiMAORfLzFb+I9qOQFr2FBsGkLVySgIUcTLPzN
vkkRjsWb7w8ftEstjaSyY0gjEnUgXu2bdkH4PJldX9NRqhY/7Ye+vfRxjS8aZ5AQ37371M1XhO7n
6+0DAgKt9fEWEDz2T7Y0frXELsvgH6XOb7UPP5tB8+lsCCP4fHec76gmlLfixzVeGQ5vaxDJf7ef
Et5mfHdUIT70d+b+avJ3UPtUkrHIchDmBZmrXgAxRzkLMjV3yYPziTB8/fhQr4IYKlJU4MxL/6N9
TAh2uEcijaYR0d1R9vvcRnhSf0bIJTKqzPqU0Ua2KN/AUXXglk9xpoSpoCiavBgfHV4SEzHaVW2f
u+TpQH7VZGrNrARaUyf8WavqWl3z7mFsouipOmsnZX20Vfks+C9PC7AkPIGUjZejvf/8mxs6mObj
gyKkoOm3hExfm8hFgBWSnI8Dex/COqxxn81U+ZDNuubGphVHW4EnSZ54g4QJV0i9FwDqUrmhfUQw
8GnGp/5uUD8Cs2982IEPyBkv3fZCuYaSrYn4hcGa7Qz2215bKrR+egoI5ze8beqPTa5MbRB61b5M
nFSSdZENN6WpBKx3hVx3QACFJIwoEuk5y42ljr0wVnJexXm0zCNEQfWuyFU0T4LlJZ7ibB3lelKL
6UL/VXCtiZEtCeSMYHqXd8RXDdsIrglPDpI9nC9/WBTrbtjnTam6TsMpX610qftPmpy6hAGmTGrK
rzgaGPK/URqAdJhrCMGnU0SR7/C3j79WyIz8zlENMe1WCwvpHQoWRUvDwOD8jv4mqfvJjiLS6At+
kbrAh85y4yzBCCXJRBUEhEcYDlOuvrXnZcCM3CsHOVeViYoP7osTlswH+0aDnf7gQjTqFSZvo4CN
6dIX7QTcv9X0vTK2sleVUSQALFLVnuFPGxVGeaTaQ3880FWHBJyNaoUa/j98C5lLrFja6uJP194S
usNc6RbB4PJUq8M28byOb+c4DMLh/T06MJunNdvl/SQJZIi0yqONplmxSF58OfAGYtEuCMuLPvjF
2rNyDdFpwAgejY61pCaDc4hzXv1DyBP9si0WPNT8msj3vWS9jDPHIOANnE6Cvw+HVpRV4onB1W0u
xWqcu+GA8Yj4FgNN0pYcpnding9gJmEI6S2wkNr331sEw1tv00Grj51oYwvGrvhBbs5dvt4CsK0u
iESou5yO2hkGfDpq7voNrBKgEnAEhCyG1KM2lFIqsL26KFXB0nO/JafurQJFqY4iIiKbZN9dWNpm
MBM5rTLCOXxY13AudGjTaPlWf9Rxdkwwv7vYI8Eur9UT6QUvbdrboRAAgyy9qO7agucQkpo7Oko2
9F0LgSMzl3WGtoFgEekmEvdTWi38a4xgWlOeDhsck9n9HHHTgLaaoKIVY5hH1kmkqaWhZJ6Szghq
hOrkm6JJAV5K3cZUAiqKwbFp0HRmRCgzMhAQoI7iChAdQ82tJuIxgq7R4796ztCGEuboQzDErHdm
F3QTKiPQnvhJ4cj8AJyDVMc+k5vUfGeIyKqw/x0grCndBotE6gTKNmNuZJPDDsbC38suxP4PVTX8
G73Gtjkwb3iBtpBxSMX8w0ng2E9do/FXaH6q2opTeI0gWEPfo5Fl2WgoOJMmDDCAjlwog+Z3Tnm4
LUFR//1Dl1AHWk7p5vk8S9pep12PHldZFdK1Ifv/IxezeFVXdfMoNkHyY2Ic4kqSO3gcOHKRR/d3
Z07bQZ/7UhPPxbkGweQKB7eePJEZTjCKtu18+73tFzy1lLofRcG7y38rHBAK0M4yD8wPlMODf5ps
NWPSRUDn1N7EbmysDEGNYCDAtLULf1G1qFzKwJsbsnxiBjIKqBWVHOj26+4cdSr8MVpTpxmGgSk+
vj2Qyj6hTXz5Ffad0aNVwiK/wpnJJy3HHQRpTf9//a5u4Vij4KXCmmSRutTEeLdbNpu9Vah3WFPk
xQbtK/NcbyNvvQSt3l2bHA1fXIykhYmoWdaKG2krEjLkkfESomkKh5E3UE3agibwz+GuuCGTKtct
ANd/v1qeVQP7SLCMN5qNumk5ibiVp8dFvqEtNndUeXdsW4I/Kn1stGG9HZc7IdQ/8aiPHRBDxNdh
kyjdHKMumyMwO3qsC68R0qPK4pK35T6lpSFmM69KaEB6RoGE1foTg7ZWy6fHSHh5jyIl0KXrJphW
jOMxSPQ7ZjkbeLqqcXTRGP5TB3IzUeSpUExQ2v2tUsQv372lUwXev9nmB8C0VMjbnv7R727GkT5x
/pVNS4cQLv8AL5x+aC7OQPZd23oaVaNg5/+DvFBgJoI1yUNZ4N/Xug/rgTJAkZvfskjDBZcIOGLB
9Bl/7tMCsHrN8wG1GizG8bkH/ddUXwDEKkWGvti7BbSjdkbNItWIUkXCF8YUPxK8rYoOQjxxG9w7
XzNpHgJweOCY/DgQ9KWWixMzxdzIZVooI7MAkyNFsNdJk6EJiezs0j2Mt8Y2mTCgNphbdIWFc/Yd
Hp1Odh/+lh/S7uUaFWji7sbAShG/uZxHkLt2ofwShn2ZFtmtPShH/oHYMRv3LycI631OM27gBaHk
8DFiS3AEho/SDn3OuBy6fq9TytVvBsyQ7DoJeITPEhhn0+cMNUBEilKquyf/OgWU213yXDAsKK9y
QxKJfaU5IJQgXjOKpceTEcn0X/fvxYov3YOlzz1HYfXZWSDdjkL6rDRAcFMj1L65hO4qFaZ7UqKt
FK2vdJNn0O82XeSqN8COqPQLFuksL8APutZgG6fqujSo6XbOYu8FAEWlDfibGGdj8wZH3rHsL8Kd
C0pXKAMsLJc2j9CKQYG7sXXvUzmYhm8Tl3SUqUr5Lf1MVb/1tN6prlmB8zgtysuK/wRVmyo+R49p
LmkVcSh0/tRpensl5P8ZLU0wlkEb7l8N2keukCxgYAXmcG+MV7oOjB635F4EXNYpziZg9YlBk3EL
HOKW/pzfd1ronp7V1srNqddPxka4LD7B0LA6lDuEqZx0B/nXNcxkEiz7PAx9sKGsvYtQ9/FHDS1X
Te9uL4VU0lqcbfNQ5MW9Lyurv+Xdkm1cDnimaVyjeMuJdrDakh8Nnz2DmMxUEoRsVqRm5pYbq2C6
M//bWbfjRsYW1+pASPQqlhkDrvxWI54nYks4NclMvMnd/diyi2HgURdNhQVUnygsGNq8o+IKBH/x
2zNxuTOGFdT+ciCTgv+HXeHKeeQeyXeoi0ieEBWL+WR9rcGoSrx1TQl/kOCPaAHmvwtaFjAmW6MJ
cQ9eU+5LYu3gUxlIqAwysKWm4QYBKskm6bqnqKI3Dk1zwSZMqDYA9Gjt3p6UuXhnCCbacIR7jp4Y
J+yQm1Q8BwadobYZDTdC9wbYuhTYqLA5mALPct1XCw7WvAh49yKKhLktpzb7AIN/b5be7UJ1qUto
l5QVG0fwAI9aZmf7dwH9vrPO2KLVglZm86D83QQw67iQl2Bk3B9UHhgCFzSCw3RwyuE8kHWgaIZf
UEbaxPrdItuFJuo4jpntlJdjNmjdVkvrkjmClLs6nQpLOWc4livQvLkyu1zT6W7uWXebMFN1tedN
mJOoD4YzCvVq97MokpQPFrYywYENUCM49gIio8nL+CCeyiPKxS5BYSkYrbqe4K6sMxPHywY4nN1f
Q6Z1lsgahUuQ1wLlDC72mOieZcg8CMAT9AzZuDIKTcS3tJ3XGX5bUKG/Eg9fTxnSAsJN9Z2MMDcc
aDN4xrxfDQ6hZ2ljHPVdaBE6fkLE4m85UboO/odDNYn++UdAVfAOdlOD6LNOtmq/6eez7kEHb/FH
epYvNmEuLkn73eP5/wGYarfT5S+ldx1ZxvvUpFCW5eJ5mpW2zlixGPCLGXuL/kYTsGVxO1vomBxi
IhIwbqRllXAGQq/H1nijXgAuY1PilUlflo6Ped6IfO8hfgmli/7rsB2U1W6jDHZASC+zEIQIlPIh
dVUwnnh8TVFD4NSF30grQjwHZOXKSbmSzR2gWtmP6gTs8VqwvDkbTUpeEquQ85MHaxBIp5ymMYaC
TDkh+wBLYnMSzfCL9NB+ZMEJmTE0GF7KMYZgmqR95VRjpquG2JXxyaQrjwuFCkc4+eOryTs32Xwq
8/DvMZh+YOOyxzj/900A2fiHtTUE+puoYr0ygx1aguCSYP/lp6C1RhMZ2hoGlxNcpebu8zBYRlsF
amygRaowpLnjX9/LBa1JGbw/Ia7qQB8dgFfitsUZ5H+lwC4TvXO80dL0tOKSbGJC2pUx5ydOTy92
bs+NKwt6SHgeagQd/gZVi1tTIfHIjfBDfXMThLdl0Agf1MmjwYhqIVuDe//LITYZfxQnnwFl2EB0
X2Y0bXxENUmCQGd2iA8/PJZlYjbr8v5I4nQzWNVzNV4a5g17Q+urUuD8zhMd6EyyOkplsmKvDr0j
3WJvryvn1kQvWDocfE5Ge8XejPl0MzEwIZYwcYvodav1RhDaLO8Xo/Ck1qrOM506DeXJFDqercr9
hoLEZmcQE96FI0zPxwfegaAj9V/YO+hmm/YimOhYPlpvM4L3CsyHhFpRIwGeY7a0qFjjlBOr1nL6
ZKAFRlPLn4WvLvHGMGmfOi504hrw/izraZgjNKKStBHBB91udo5sNyJ2XbUQ2y18Aax9WiOuFouX
CdFp/oICykPNa9WQdM5eqvfAcIwXXgLrGyqcytR1YvdY0OZP8vgBsbgzcA27E1PGWyHW0dasWw5N
osrZwKISQHzFNeA7ZMA+93UGz2TSOBQCdCqMBI2jzB/FnN5MbvvnMVvJ68hLnfNZ4R1yMRgCM6cr
7nSOcqd6sp3bUvbLltgSgizC1nvZfgsFlfC6csfSUbEXu/Vc4SbOeLLASZuQ5y3PFdd5SEN1s87M
D3OgPLNYs6zR1jPJofchmfzmV3KrEoCdtPWJLji4UpUWSNmS4EkADbmeLTkZBlVoTLMYY0d3Jm6Z
r9kGx4yPOhrsFqcf5zmEVO+ONod8kda8TBVVN69DU4uOBW/dgs+5pYujjwJ3BkDsKmVpvRh0KEsd
t+yrRt4SVcVX5ccdgoEwlLn6MW2D+kn3e5EAq+lMnQwnV8SLZykHcD1/l80S2kIy1/KfGS+YJKsr
pPWSCxfaXUD9AHJonB99WlA2SPpmKBeTB+Z0ot8HT9S7SVNSRhCouMu/HH4a6z+WTxcCWJYH8Qwb
aipMkvbFz/eek2IdyL8rqIVmlV+Tvftbeddi63rFiuGMdOzCNA9WYThJE9wdD3AXLfC9vJCYD6a+
HlFOsmj9b/gN7vefmILLDxwpzscQxvUfwj/C7tAgJ/ZZIDdNf481Ws8VCSN0+k9Isvi7kPaF1YdZ
6S6OFBhkYAAA8KeTV3TMX3OMJd8QoDkP7gY3PmuXHEnpJnm77Yk2Vemll4rYflxRmbtY5vxxCcqQ
P7+ewra/YZk1xIUbwN7X/g/yJS9x5euUcAHx0HuAdlhudivsP0m1KraBtphUVCaHd9UXnGPjHC/n
qUIjw/VumV2UN8wSvqqniKIAXzAA+hMCk1jpU3ijk3WrUlfRvB1aoCYPV2tGDpN6iaodjnEJ0tYX
rKHq2STMzuIQ4TAESWncE8E+eJ0KUShOfZ2fsSo1HSXsjzUhUIp8T1Lu1Uze9zmlU1CU876YTnj+
xJkqrRbP/PH9OGRZ0rUu2XUNvsEsFJk+xYtV+2RuVeOamEtvdlR7FMJvpT4fI/MvwRT9wMJ7Yp6b
7LtlOn9VRacW9KFfqRGg233CiJRunCaFesFFJGmLOjFI+6jUY2cnxNsuexdacAdwckHt5ggOOnSE
maIB56sru8q3CoKOD/pgK8wZiG1jc6qB/aHVgIUDFLsKpHLJDWf6JSshw1s4QyNiN5vQcVYvRQxf
BL2T0f2qaVd5v+1eaTnEez80OwdTgTgcSx/XhcOKRaDNj3NAlqBWS3BCaU6yNyA9gcZCGvTM4fD8
HdQLXJLpXatLWwCoEgfld2NcblaAY+WQiJStn7tbpawvZsd+9Oz8f4ASZDCEvg1Y132iZf5Vfmv7
dHH5eCC0zyiHOCEO9gMMsV2CPAGYUx9dzLaN3bedKH+TPVdYYIUSUp68w+0hqWdSotcM1pQ4i4tl
P+JpdcV4hk/mjZNa/62yR4yt72eXR2oeAg0UtYDZ7hLfZrStVCU2A66isX10alxHP52TX5/AFMnz
8CNZJ7YGhknfoGvc/D09Ok6mX8zdWGWgG3lFPoVA4AIS3lg8DxQNosUp5SocKodo8bkjR5tfk922
LS27TCBKIRekmT+nTnUca3/7QZnDYYVuZ5D7mN2aExPu2OaV44nZ5InEjG9zLlaaFIVAC7bBwk9I
HmmfCDSkQK88t+xKB6G22HN1vUYFFsRhVTvA6ofQWI15TA1/0QdIUhDDdxV+yleVt4md7+shPrLt
t9Rps41eZ7txMt33ZtWSkZBxnSUWNuEBSfRK5qGqbj7XkDMuOgYMejtmCvSjiSJcp7BiqFM1xlYk
fHAt/5uqk9ZSDfWenoZW6zV+1p2wTqlxlCWyRrjM4WKFJzbeV+qW600Zmdksl2hwmbOud/ZSXa6B
zus30a7jXv1eWiiaEJFNmJNioeQ04Ihc+U4kOJVrBRZZRq6MF3fTjaRm3HZjp++jbDapBgDJkqkq
5sa2vkg0j+mZdRdahaRUxvzBD9o+2ywYZ+OBM13OFpNYWaj0ZbrR/msHFOUIWt/O+uDsHePdLk1B
Dia1z75MByJNtOfM553tk9TqvLgRuUt1EPMW6vW15HvRIjtyA0Ggejc546ULlL5m5iemrOCpAZz9
FJLOowhK4x6oGZyhX3VWOn5Z0Kkw/zhB2CW3+PYbktcDUhcaTzFPobXi1rN0wd5I8OwmpIjBG/XT
yxfV7ARwHiuCN6nW/j9tnMKutmrsa9B8ZuuuHty+RIVWz8rDl+964md9E7S2fvpaRf/gwIMAM0qu
oaMvLz2+0kGU9L72P6WN5d1L+IGhURNliCnPUpk3uIhPgcIS+CfHPrKAR7QbIFHY9XIcdaYRrAB4
AXAedkPyzLRT+JSdBjsMoeGfQpK1R66ZXbkMNXJB6pbigjtrVuBLV6uiCBsY1SOyksxHuILI7DMF
F+7seSMGioRH/f1hcUHmMFWVzYOcDfOe39DF5ZNMpa7MYyS5/vTKpgxqZU5CXx5vioLiI7Qs8Psq
An/c8NnmjJ92ajzv4Y2jM42Ci0eAg5tKndZH3aOPx4rFcEVeuckv0nW/k6WTNr7fzUGbASsAz1kx
2mlelBpxSGna31VBp5oAI8w5XnwkA8F0tFzAs6IQFHVyceJgls8M36Jt5LFS/0khjBwBZLR9llnp
7Xqx8WeQcugqDYck3Y1gX0dx/ogeDXjhYi4V3yIAsApdL892Ud5br1sCjQgfyJkXnoqER4m2DPRo
VrTymylqL5BktHR4GORAC/zJIi36sCaWapefyd63s8ZuuVgYBesbjwKHEzfubyfhYkACb41roLxO
oAC5l56S8ik0wvjA1Ouuc5xWT/nsV2JQJ5OLDDpXVXC3reQ5yMB/8epKjBdlgDD6qv4NibQam9Zi
jm4avdwQ7wfgTzskOWwSp3xhI7pP/CpAhbtmeh048+zPl5IrEzwX5mT4s3WWU/l6PbqaFNbU8IlP
mmGKCifer4D+gYoYhD2vzuu6JFfeyhKC0RUU9Gt+YWiseCLv430mEB9ospG1zWWtBiMJZZD52c6B
30sbecLiR7XOUwUIVF4C/iHWJq8aqNkDtDtoCB0yuxqqAcefhN7stdOCncPUlAkOloo9qGrvgUC3
fPUhEeeHMIgd14Yktaev7rIfmjJmaFrSfUtCLuVYtzSJo2YpdE11j15CGpSFalTOdbF4+rJrKSdy
9GrPwzfMdGeMeEXXUHrbhVKMvlIJDeFJfns/pnrG9s2FaTX8qyBgMpOqIsCnle3WlZRJofJNS5e0
j0UmYPbH2tlvXkRrbfBlX216ca72bQP/CmqL47YjLjJmYPF1HVpr0LlRlsqkM2kjRjm1/dwEe1Ic
gAPj0iqTl42JV2O/7ak19pTxI6wlOfF8F1rIr5iX5E1h89ZMgCAzNhwo8CrRv0+pKAsXEzfyHKgN
jjBSpvx7KoiyUnAvA94W/ZABqMEM/y2/QloPl+nKNgeoD5NSJVCedQwP/5W8FAsgYita0IkkUrU5
8URDElyqEWew40JYx4HWsUyWeWzOcUnmDERF6pJYOjR0lx6tISqjzOeC846ehd4MJzz2uBz6/JJe
0Aketoccwv2pL4kfS/lSohmVwqKctQ1HrAwOH6TRORg1fIgXFP3VtBaayesmh9LTAGdFHhmtnwIp
G99GktSfYt33xao06scS7RgPS/VvBfO0xxZJnmZVHq0D6s4Guuk9z6Y8/SxLtcX5CScRgm3iNLCO
rjXqtlyv3vl0iKZL96gQyrQGcHfMkowpA1YRWB+QwUvfRq/+3gbNKlc/YWmsFOHfX1duHd0EmHFH
uCGGYBIZAfHjk5GiTrPnahqpuLDV37NA+bWdtvDOJryDWfpGH/DrB34iRA9CwVtYPMr+5RjdDIyT
JUoixMQB9sP6uQ8EwfsWllA7BeniULxO4u7tJJZULLcy04/+Yu1eaDkA+al2/O44zdOWIxjWFvPb
G+V8ql5beytCTNz+sD7fz3EWG/JMNktn7/1Qjo0D+J/47CUzFjWw59Jyy8jcsIkLD/0TvtLfmEXi
ehLrJHFAsaZdaHymQkBmSnw6ICDOKXNE8f3lVMBQFC49DiCObmoTX05PAzpeWMGnI8mz2Vnjlmuc
N99TlT9eYVEvld+d5KXJk7Tpj7jVvt+ey0eLn1luV8YUgyhosTuPuj5L5YW7wpFCYR5uXDJkDr7x
D1EKhPLvy3SCnZGR4vmcKxSQ/ttyWb4BKK6b1RxS7mlKRLcxZLoE3n6xnzzclW329dutREPw5eN6
Ow7OnDZkKEFQzmEWISXmudtIWsxX1CVcD0gBQe+lZ6KvMk1pzhfGj6OxAb4jvwTg+PRd0v11pkSa
TyWhdktFB1TBp4o7eCOwjTfGjE7HuHBbj2MHWk+8c2h2XGFIxBSan9zcRWaoUb4b/3hK/vXGe0W1
29THTc7fuY7Uh9MmqQrpRiWAAw4SI6PcQiuR0lAo56YGAm+SFFCnfYFIEV2DveLDQnVj8dqVhKNz
DKH5jdUN31/ODFj/D/WPVaCxxkkAtWe2o0ZZg9HBqDGTGZu2/8E55aguWhuhhbfrqxPbXzguilk2
7nUwkDc5LODM4uG+BJgGOyxGr+n/3aIAb5Ym1kT5YfyeDznnTacdmWWcgGc+TYiIfVTxTT/Ao3CJ
s6n9xPaS3An6AVCblMJWwA5dvq+qhR1UJZ58iXATYnzHni2er6Ap5rIBSPzW94774XzkObUS2ZBI
YMHbH6eutTxLr6q1k9iMUq3ZXIiujdWBxA1hd9dB2nmMbZznJ11ViDIfDxl178NyJmw+jcsH9AAl
aJxhO9fq58Gwv5zHwam+oKug9Cs8ivbN6ITqCNE/gTzBCeUCRTEkOvhEl/uL7j9Yw5oMpta3T/QO
YanJro9hba0YHIdUaDfKT3Tn1YRT0w9KWhMOYyPsePzpOChLxXSMTw2ESsRT7vCvN4Qi4N4nUA1O
jDMjFFBZHROWrCv42Ti3qmotf3DFGdEXqf7T1EjDMTor+b9XeDaZlbEt7ACLo/559Sszaa39WAC0
SrN28SIWsBFviZQn0Na2gn1MyXs3Uw29X6qsjViERaSvtQESV378I7sTM7ttU0ZWfpzG7JziBRp+
DqRzMDYwzAtq6yiM0bAhre44FaVrj0jCJKJ9Lk5TEM1HglzjWgBO3H4+93Tbp3aJ25VI2+gqcKZU
/hRIFNnynbx/dlaP2P3yg5DkMIsl4UVRBAAcDUfd39QyXprCJ7d4seTcGc82CXArK0ysfmIxDI5a
2KEvNxrqjZT/NpL/WgBKM3p30/3t6kYVlrb4xiSDVm8NPxtZYQhZ5W1rb/ZpCCOnQKFelfut/IIA
M2xXq6kjb0nuVlX5+UK9xITwdjnZnsi5fldnyPMTrgDR/ZcAyMuvOgO57O4hqhTK9lkAQD3iFMgR
1/bqXYmKERQkZfho7IpCB3KrQjO6l3CHZjY10K500ZEvYNe9UsXTutqc+4MG9uXpfbDGJqsTOCIe
F0ON7K5r5anoHdUrfjJEpP1stMZ23/H/ZNw6nLnDLvHQqp2oZBDorDLVV9h+mmHQNzuWT2EiyOa8
HcEAKT7rEPas1Ngmu4e0CiUWfn4akU1LQfqd+7x/XzfvgBMwQyNFqgOn/Z4pFDJ0a5+xKxDUdazt
rTdcqaq32RRh8hAPtennSKQ1moNVAljQ6J45k1jBmSaskRqq3oy7PvvB+6Pzrf7AFzeCBHecGRet
JkgusOhp8TFsRSIimePJUhfKlax4jxZcXRVwvbk2cFHuR5VU5Zob5gQAKSA47EaFwUI+utRgBS/h
VAeWqpCk3TWnb0xC1dtfykG9s5H6DgsCmNbT1TI9RhlRpW8iGfJQ1IJEOpvoyjxUjcOytS4zJWFP
sFQvNq8CRU3htidVSjVG1Y8RVb3AB2xIbKup2ejj0a7ktUL73yBxViJGay41xWQBbxjllKU0WJmZ
sMoin/gyyo9gC4hS84GmVg4keRp/FJZkMsaTmhzMzM6R/74v9iIu9jRX9i1k2LFJ5ohiVf2jJhDz
aAhCJwJg6uTPUoyaFy7JJpD8x1RPPB6tcl3gJLHDiqD91Nhn1F12IaWJFl8qWdjJQg88jhYwhUsQ
Z2DNHvOuH6cJrnCgj256DYM+fd3jYbA9R+UNzJNnxwnDCaI0zKLsWC7CUtfawMKSln/jrsrko43T
9YRHbmMLHBLrN7gh17HW4l9ENjpxbQKGmlCCIX9mBHkI9VPCWIjiFiOrVCnqd3nzrwauDUAVYPA3
XH696DdXzy/YJqMy5am6l78JW8flGgRcfeGkm4W+ISLHnBPNE80c+UPNyh8MRF7EezlAqSsNJZE3
uiqgC2monfK+W9iehMREJqusXr8Ri35RNnsXPsMYKO9K51VnHhtDPuetVxIdxlpEVfBlk7CdLM6Y
euLPdXA15lE38tU+iHARxoUgJnhU3fWd5r35T4ds9D9l32MS1TTiVbgimi5rnI6d9/Tn4QGdygvj
qUUBKH55W/acTT9rbYr2uDIXYOdTi/y+ulBspPlxcOhxIz8Y7ca0yJxiMKOOSEBkjSu4Zjpb34Nl
A307vCHj/hj7rGrYsR/OY6wTGmCqsH4dKjqk341MeZKsoCFpvDpEJAtbSKiSB4SkWOcEwTFWzy9x
TgGYgLkcrKnhR7HsMRHqq9mnStG7enq0rfQ3G6qDUpo6VI3wNZnV4WRy7oepLmBr/2P7TOGxhv/7
KZ2QouqjvVQvveRYsusg50mmuThdCEh/MUvaafjPPoH6Ee1HGv9qql7263JP9aUwr96RcU0el6Ve
weMrwC314bxAPRDP0DjXNUg6nzd8ghSoMlTNKIA46zZQ16UfutYiOVd8W7w+ym1dQG+3sNLatDmr
Nz1GzrG3yI1371yxE3bDqOaziF2az95VdqfZDZlQeZpuEh4Y+slvSVqpNteExtSKb2wmQe1O+kq+
zQyDb4bS+40H8FSmg4TrXLw3BI1DxL0amHwpG6asoNUJZlm1z+HqiytHycsKmb4S5Qifn772AC4n
4ZczvodNyn9GY5FmiTU3X/zHmng/2+XK5dwhia9Z7jnsog7N959v9v8UyXR5wEGVnsi3MX9JJLR+
9rVOjErrBk5Bxr5K/ILtk3vUd2UUcwRavMWP17Ui489Dy20sBgCZTQ2Fvapp9riImKQUI2sXGJ4A
4xvnncuywGi3RcLbQ3K7u+0d+hQR7uAqw6YzgI2zoSHXNWJ/69EiEG/CvlWAffPTO9ZslXoL3Ykj
Bh5wKgMb/B9cDvFvCch8na245HOWV2WIYeGZugQtTMKdSpOoZVUdAamQjhJNPZSZ+xY2PYt74E6z
bqVDUKy1dAx08dKqX8HCGgz+jw4tHObs2G5BVd6v1V7xzr3tbRc+bhGusot1BDtdQ8z9SKRf/ngz
skYE1+zgNwPORYLITkIkX4lfwDa2gvhM38sCW7AjaZP9odQiQdTPf4Y9GXONt/6j6rLb0OIPc3vs
5QGBC7bl75suGDgxbrRlXV2nFAqHI0hI36s/DTp8Lis6vXkiKYJM95jxO03CHIGHZ8AaTJwK/liG
Y8cbVUqvpd4UdzgwS2H2NW8C6JkDHkZb5ZhPDmkp8PEd2pe8XiB614UbD/U5NG/hEHvQx63I+Ko4
DntSUdA9iNjE8+vYYEf1vQJSX1T3Ma5TWyhtJ1A0FGUnpgyzb9E1ond2Q1pQmggUCPZresphTcsa
H88e/S5A45UE4s3nnxTyidKEH8m8/Y87sdV0HXgUBh6cL0pz8UZNnWlw+7VMSAKb9jNDMgtluJeQ
kiqeNqHF6XjmeE6vscYiR1hl+3zUSGIPsaRsHaI0sHJ57kbL11i2cxxP0NybE4Wgv6z/ghX4IgWY
Z846iQRx8s4YJDbWXzs3vH76AquXm+swLcLNcQrMy1jktFujWk53L7wYeb0+OqwuiuEI2oBA7ldO
HsyQsdGBxV8DiJ6MmgkhE8IX3nJDlUilovmcl4appAiNzVC8kV4GbOFcVteSp1hHPCQtxmRbGkUr
9KkRRs1+vzceAqoWXLjzvZEwbYQM7+1HiJxCNw2OXnwo3OJfctvcpW4/VFuLSRRkFAjw6SPVJPLw
HQFr8elECszrXRxLQ4ghYNBYwp7w5M/NHr9QKcwFl+f9QPmkAKffs2cc5nm/Bt1oOSVu0DGTaxVD
3tJBiH9RhBNWO9jny3nSe+VrrVh9bEAcwBcbFoseoBajPnfrgR5/Tiy7S17SV0neg3xleH7lWpKV
G+yaL60SNbfUFrqk0r511H2DhHx7R+yPZt30xEsvtu1hxB7PTC3030KpyOWm8OIUAmKrJDu46Ael
ohLzS6Ps6NihkqJvPpbeI5YjnXIekQBIkZgCH0dojGylDckC6S8Bm6WW9WTvVDXsVD5MWc8ed/tc
hYsvV7fANak5WtyGrouTBrFJuXzTpVu0LWHQBLaKRfcw9hSraHtZsSq1IgMZ/8SG74wMd4kzvEWw
aaPCYvhDG6gUz1998kOmMWMHRPi1iLrP3nJMUp46xVOzgafp80q0FZfolDPiwivuKECN0ZDIvexN
B3BTJQQBb6zP65KrQPVS4lYBnFhNi9Tk9o/H9kSMxvEZ8x4EFiIJTLmQ/XSNMdh58pBRDMGLhSZZ
dOXl6jMXksME/Mf4j8/Ry7a3R8Sx8DJNCbCn3NZRIMFCy4n/kPBbLqb8GOiSjcJA7qRLyYBprCG5
pDERa6V/boXV27xCLMH2ml+5/eC+HscjrcH6eCANwQ+AOBvaMKY29tJNmYa7iIC1maoXvH1qnvU3
dGROXJ4jtuSVJMBJ+nX+KdGKxrgF4K4dLWjCrOS3+NnYb2vf8o+K2tfuIhnYxzcwob2uYvMhH/wy
FWTFeND5mAM7WR5WdZI5vJGe+71jVa5lTt7ZeJsF0cdMtxsyFNi16FzGj0fqXdZNTKDpNSKMFDC0
uPIGkEocyXqtLuzMplCKzUtswzP0AId/u8W5nNI8s3jLtCJ/4MCWRtooJpP9yy77I9K1o3T/SFoP
igUvOkQLMyvgaxJRQamgTVL4Vb94WB+qUJBmRABfs9rF+x42ajEWhVYOcWVptmX+SguhXug/IDFH
jH/kc9nNQjvXLII9nDOMUJufWuX5+Zeh09EqdDX3kuWc9Uv79KjyZl0f6t8xskCeRK/INnb1o8YK
jKSnU9xYH53nFnw0T0Y9312sofyzIGqcCtOWFC4qoqkQ3BNWt3BXu++ty1w4YtMAgximd2itBjlU
1JdoTYB5anfALJ4PeqjfxMDdDox7M3dOoU463bFkwvUCChIBFjRouAIZlwIdj2S3I5s0FG7X/5QM
cYR5/kwa2zUS1zclUWrL5AG0YC+e/IDk5AjJIGQJ25/6SnzO9Bw49VQ9op3ryYOhLSE0OcHBE/sH
PyxG+MYVinBnjZaX7VujDCjuEqD9bzfp91bHmIfkYTzn+W96sGGFBHGs3rxlzzgVTbNCiQeyUlZY
ExxB+Bo5a4stZ55vO0dG8yW2M7326OdebNhlg9acr50sTRgtM7gg3KFTwZe+DF8A0Go2KbU8y+Z3
t54Qy4yn1YkycUb+A+JQO4msIsXcJsOJ616TT/snc4rbre2PsYkoU9ScKqjEvN5ZYxK+6KEjWpRQ
WPUSG+Ov0cQuLWWt7nzYspI3HCHQgMbyeZt3j+jMq56YmmrXRzfbRrztfGFrJLFQ/qlZjapSWhCF
LqP4EonMNcy5VxNcoarAmey1q8/q+kH8cXmxlZNOxDeo1lMo3p/MUwgPcHDAW53aqvetMlHCl3Om
R2B57bQSKUSX5PrxTKhDx999zCXadK1MmORxbxe9W8uXSnJlQQ3D9eqxT7voYleO1rjJ8nPwuXHy
DiYGkwHOfS4fI4ZPdSMh1Hl7xXq3ZIWsHVJS6Vbzjv1VW8NnwprvuIh6ivFfOTdSU0oAcMhx7fHd
m3Ib8XM3eXIgEcuUxt6fkpvkvpp82dQaVl84Q0OuxWP3KJoKBjW4TS09QBHokG55IOnpWm4BrZYf
edcFN+QZaeLgIbL7k9BTeVw+HFHKjjYIyxe2TpRTOoMTULLuUJcxMTY43WZy1FPeZyI8x02QEoyP
VCBJgBuLlyxUxNYGr5gHrTFJaEpd6mHU2G2+ZtceAOOIwldiFFFP2fr8YwXCTXakWOXU1aX8Zhz5
MvbjReNuDQB+/ZCvSwWd8v1F3mesljY+qX39Qp2yNbngFdOoYBQUzhQ8CAfHpKxPExiu8p3nIKhA
daSd8NPlWwHSO7aJQ9DXizzoBn0w2YvSg5hmkVaPLg/PE6mQFXnVwlbWS9sfBObi8YWeEQG1ozV3
YzQNdl640WFQ48tvszO0l+N0wO63/6Df0CGnibNwn1qysXsdTASxuZILbcu0vtKjFlodsqoZUaX5
OfRS5fFEzCYzH4DqoFt+qEMEDRMFDLPDeiD90Tr1Ec18CLpqKnQv0pGVmRt3+uasOQX5GBNDotId
tzSOTlaSIr+4CQ+9YYnmAibBhr1WpuHgTjHO1eKwpRBsmyjyklfBTJbWFuV6BfBEVWYXbYBqHtf7
w8tJEuqt61YchnPB6dLgrrxjNtKexP8SHBbhZmgodS1fZE4Kc9JPOWBsOo6P6w8CeRR4G26WKbPw
ZDRB6j7Xsro9p4YL3wvX45l+IQ9FLqb0oRtC2gElvbm4PO0C7+6m2wTBaiQsWZpHIWTCyS2uU8zp
asjvWdl7ctoum1F+/nGrsLmPZM6uQhUR54SERHeBK39uk9KPzXSDwBH2S+EFyfRk8qsuBL4Yk6T+
O3PJBFa5LpAjGgFBlzWF1pNzVIXkbeGGiXbHUKMrVEnSxeZ2wGckQnVFzUPvQd8fBQj6Hi9/YODn
nmKJ/CHVWGcEHu09hnzzYNovjh63WQrG5LVjaz4ZvdmTphaVKTHDjHSRry6SHxEH1MICAhP3kvWN
RtTHnuvotTkBgUrjyjQQLth0q1xCfxUc21HSgoD84CEyDw2vKVTbqdnjtBnkVnN+62H+L1KQuWCi
ZwVltKGJRvb0pAGE+O4tAva+puSxypWrbZ3BZ7UZ5v8b9Ii/C8SWkm46lOTr5ykRx2Nj8u4zIL+V
EMMiXS4edWv+8dXUYW5fSaqr3f9HNw+ElgOQT2eufmVK+jktw8xfnKeLOnhYP8zCvFyMXZtRqSRA
cV3fWrX/eOZjS/aOBo6IrdeXatsJSc4jDQ49oIyQRbSf9XthoAGJIiOnvNjTwq5Wppd5SG2sT6LY
48KoQ/ZmgFHkIqDLECcsgccXagzcnt8cX2AJK8wcJYFpY1+q5gouWcGMo/90neNPSZ/lC2/gCBwJ
vp3zCk4lOyP4xEE7LtjCO9WhmssZXsYxKVvVSURQDj6shnli2LGoUWA81GSJMqM+7Yg7Y3WdFqDH
bOBvKcNfLjTWUgrKsByHO1+zTgTyshoLxMru8DJyusWlXqFPqR6EeExeBzF1L9D4I/wXK1qo8GV7
qhf3jBzCPDY8c0whi3biF9dYHzCA3zOpO276Un4+w0P0ITZg/ag6e5fj1ptmH/PPQOurW+epqx/9
x7tRO0W9D6f578fcpQ5isdDpBDsR7HYgSPwQkJ8G1Dzr3IuIx7R3Gn9AW77YfZmxfabLZL39R4/b
pTWpRup7jBDfb2xL1xNECBXLT9N8nJ+JUUPVoirK3MkOzsSXzeEsOrPiTbYTbajemvAan09eelaU
oVcnioMw6CeYBXoHPJQlOyH+z8PgOSg9YtH67+xXlE4xzLfpcotwk7opP7jS+gbHyO18kEobFa5j
D/iH1g8OBnfw9RfIBIpjH8t1X+MsxzSZiY/jCzTBCjytX7mIXCzT+3jrt1XDsNIjHVWv1WzILoJa
W2W3Uf6uHc8bxFc7qr3JF5Xn5GybiqSY4iCI4L2hci08FGav6LEglmUejdIZ0LMVaBIiOhGLdcjW
Ew2g4MS6h490hcx/oZys05cPelp3A+3e8AZUmth7UN4CMeE/xanFjtWku8hl5Wc/9xXHDfSKSqvw
2Kh9d2e8InkYEDVjvpIf7Frk78O9E3DfSGGqnlwotm3VHEbbjP9MNebIOFqWTHTr8OcBRi0jZ5Mc
hVmhcXr/L7Ss6NzbF/j2FMjggz1K/2KEjw5eEq+lZbfZSjPwxspzfuPTS3GDtovlu1Ivu6liAouY
iOpYS5Ys0/JeZwsq432pX0Cdbj+/s8uQLnxIionND+KwHLUbEmAyu2AYhgzgKxgeUSxWEbG672+i
kKI8kB43SXftEUOPfjC/JardLQH0qmJNpby/822uv9/C1LMx7n1jWIzw2NQceYI6UVLqO6wiN3dM
pvKzoDApilSoH/PIPTm+Mt3Be6agHLBKxS2rx3BBwYYAFXYrhf4gGlw1P93jdgIGq9TyFnrizDry
2wG7/L+4FTvjvJXH9cJO3L/wc+FN73OeEtv3QjM8e5TniI525BW2qbmSmLfjwD22NVy8wbc1DBhz
MDjBCnFH2Al697WxGh9XYksJAPdJ7drLAvh0n5ERdKVeRMYnUXLrLA985VW0NhKwSawAILAmND+f
m0IsjUIB1jBgdDzUvRfFUnV2m+jclYY4reQk5vibn0qmxDkN/rzMa0Sqa7hsxMt/TY6dpExgEkt9
kENNEzsQDYs6zYRVr1fyah+XjDBW6Xo/jHtPAsIhkZWo45onKojkPEBuJ+EbmhI3w19iB1xr2atH
qP66HBmlWCWSuylSD8uYJjaNK5NgkFzXYR8GvCxkok0LM+Ni8xYUfq8DgrIqSePurw3/2SaHuOx8
WW61nIS1wb4ZYpcfuy2mgek72+4tEpej+JTQWMtMFpRv1sz1tdwlQyhnVWSOJYC5VboG6LSj088s
opyJfw3xTJnTaHpumFKwzY0MpDpgzWoo7iHP7up0ji2bQn2UthmBNbyrZSue+d/nJzaIkQyYHtAz
g8KdKBvkbH6pEcy76YpfDlY/c+anfrGClkCoghW9Lu7Kh6iV8p9nZGqDrNg5T5VF4Q0EDOCEMeZr
UDW9ASNTPscjHSyBLqmZWPzM00IXzWnSmJ90UUfcbw0+VMCxvWfL3u8fejKadY7OPzazeVulIgw/
tJN7CWkuRh1KbvvOf5A6SruGNIUUHvyW1EVdr04AdWsAMa/ugJlhFTpVg68bu8NJGOtr05dbhI3m
iJk/VJqlGyE76OrlxQ45j19RTGcONIZf21p79twxHdztI99LSb0srCMw1LIgL9zYxVx8Cjxbr3nx
LaCTPTsITeptlnVZNHzbkJOTx2ZAWikZWQP61Gps/yCksID5y/szAbRTIm4WNkTKP/VhkizZ+jiX
PFog6XtrYs1nEtFBKvyFLlP1/PolPfiA+hYXnu5Lk6Ftkx0viTFP6qTE6PQrCGA9ZPBchWgJWZA4
zXLAhtsFXgw8NocSW5bPAx5PKIdd6+IhweZSl8qpXUZI2fHSXtCyAQgut2viY2rs7n4kUYXvNkor
TaKM3TMio6mcYOmm/5rOlqayVr4l3zt1w220BhyT94tW14HarEKcxOA/p6FFoZ5fu/KI/GvCFEMt
orQaA5iOYCfBJbYIBvKhaqa6AXPg+wXr4+RJ1gHyGR54K2SaxUPrUlaBtQKs2wg3VRMDF+JikNDM
n9+k/DIc/ye1CHl16lELsBBkJE/YqVid7ETEFFn6YN2nRexcOZcqdUC4COBUfWiLEVoFlzgKJRXj
5RfpSxN+zC2304XdLQ2cBq0TGbQGVuV3NSlvyEfacdQ2f2dQP8OWWrV1WaSu87kXM5OnLS/tpxSG
XP2hcH8byzBn3B5XMR2VLJS0YkDan1OsJyCkafo/nWUXSKhoQoznqUqrMtSXAb/W7Kkduw9fcFvB
9iLEQ3DbYU7R3rPLg3JCbEgsmSDcrz7iSf3DYFqxzFzzE0pPfuB0aF42LOo5E//uUR5M8lVToKaY
wEIyA0D1uRzKAzdM7ZgOqgmQdfiMLpVyVFtuOFziSZkGnLEP0o4Njp48CyJFm4KcvbLD9CSlg2bJ
HPPmUnOB3UwCdCd5a7seeV1rChbB/gQNqq4e2nmutws7eo5aSRJtssL58QXDPYnqD7udkYkMf/UH
0I8b9UKMH4fT8qdGkbHL2SWVKz+egEWlz0qefh6n7QdR0C4nv2c4a+Esh1COPxyudHy/deLE9GGL
459SNJStVbWdPeZavbaTnI6jIyPUjGVz7wISK3HWRI3b8e2Eo7Szeo8tvL5wlnFfc+8dOQpTDfat
0Y33hq6FNAwPR2+vqT2+5zwr2zQ23bv3VkJVo+A8n88eYyXvIsO5IyGT63BdhqnLjoCVWX71gl/k
71ygz0z8+dkQnyd2HWhD1DiMLW6Gu5tnYGGZzNDjdM7gqq0ylREAM46sYOroNDHSJY/VbGuBVNjI
oATh9nGATMHI4Gz35ozxoiySXRtKGoPcsXH107IccWegiy53ETCJL9whXgAVlAoDulTn3nhrerXc
qwqF1xiYkT4zHcJTH3XJnBL4Yl7wBzDEH/6pQJbW/9g+GI0N9644v3jcEW8zcMUhl/iJMLyKG3a5
OL5DEfAlXnvsCTzcK6C4EFdyhZc81DssukTvnzGx+0li4C8AAih5C/fw7BwHyfiMxO6GnKlmr7Od
AYuyJaXvTTjGPh93q0+hesaA5sSPiYqGC1elpYRjuMvh/HK+FnZ88JqSD2hg/JnPaFvNJU5WEGxS
OBwbAC0hE9U9CVqTYvBidO+rigi35TlCByLCeroiIQDTvUEqf47Yw1PfxjqFJUx5XJGfhqdd8Nso
A77oOX59Qr6l6ieIdG4T5ZHiEnAKJZwM2reuvXVGQLq4ezuwTOAu2teSflcWhkhRUYCRzS92R599
7OfqjeulrkhQsHRV5jrAas2XwPyhOPCc77wR1tDHYdoS1IJoslGnRkGweskjIRqnX1JjYkAMOps7
Kcfz15ROw/18fuE1MiVxZ+Xb8bAH3tvLsXfqKVWsUM2tjtAyb+vCNtpWzQ28QSPKZfNK+bXL+tC9
v6HFYkP7VXwUuouqGbjkf4mRIUmbeQuRtQHKUJDaUdNZobV1Z+PiwrWnSHMf2szTMVLaR+8Qi+DC
S+ht7QW97qe6/9rzjynPWRv2qhGwjJtJi6df7/55cBS48GupgPbjatN6CiN3VgEb/47jXVgHfV1O
wMK+hr/JgvEV+C7BOOXKSInatlnWNMuX7WRdT6MmP6W+fC+LtGZgwgjvlCPmobgIvgJWFtoN4PN+
7dsQP0LepZRzd5kPPLBQyw+jEyHyIJbdIbiDTVFlkb3OUQlkiF3RJO4RCM3nbGEWG45t9OhY+LpU
Jf8jbYmAEB9eKjqLURk5IiRLc9ox39ewP9cLU5fVPU4ho+pLiNjprY0ZHo4J8+zby9ij75FBLhWT
t3UPx7zkdIv33fdnm9/W0f3of7nbrssM4ss7Ysupec+AQtqB7bbOGI/sEhv4zf/W5bYhHFqEpRvM
CWeR+uEtQS988tBe/iLyKBaixO5LJiB5OHAm10DpcKqgn4zgvz+4johJSqpKrwtQ7MNbPlQ7+wN7
BdiI7n0i5DEmRSNZXOgkmGkxReCNUc4oo16HssXM8dCh58uhi+y0BSRsvPrl3Sv6AKp4k1ZjGI+l
rP9s74xiItAa0h/CkagP/pA0uj9OeKavihhA9BPCkNcwNKxs6EnZTAhugbdtCgsXmCKkC1yuvN7r
x9ox42wKd+0BB+cH9iR8NMOXzykfhJp+hsh1G+dxxwAGTGPj/hHiKGgA/pNWiyvAiB9z67dpmDUY
oGhllBuw2EzXoA+1SNQxgO9VhaRNfF4MO0Iwkd0vla/ILEFjJRAw5rAWeOPznWCt9SpDlJ72F4Bg
Op3qqPADqS18rmb5Fs6lNc5wVcX3jicMSbT2SBbus3QqLcPEoLyR54Cq0cfhIT+p2iGFmJe/B2aK
7LcvyLBaRtH/+ISXKd9uRDHFWn6Z4fNoqIR91dbhI1+q/U6WAxUV1bU5HUYhxgY+Z4YdBdG0wfHa
4zGYf5neh3TFnSr0Iwk87QxXHH2hald1ZxTOhUcgvGd2bQm4+i2FTLySeRdqw9ZwHWK8WTAzolrQ
sb52iVcKCWLpdLGhPcqH0PWAwpjcCnkAvOli3Gxhsi4VK3epFx0V4mEqhLsiL6XI4QVizFkvLHLo
OX89RTzDUcWKlUghtq9ka7kdWx+jkSzHZCW9TpDA7ip7UFS/yHRFPc55sqWhAMzvhiq5RwLfcWUy
JpwUkae//OJQ1IMWPIeOTKOttJGgxzKSYHroLVrnzBK22fpb2gE1fuPIIIKkmRM5uXjD+ckY25zW
YlBQfM9rJsyw/wPv+gzs9fhG5l9D+BIc1JIHOqZEjLCAyb6mPpB35WXOK4VjgFEWgsKJyl2tvLwq
NiRE6hSwRSfYKReBD8bgmEAajdkj2JaRbY+B7TvYG0o8R9Uyh1uL6ABgFhlcp6iuWUw8iGkQ8XzW
WtCyUxWKboKeM0cl5Y6Ny5lFrXG9GTUoc8tO8ra4NBoJ40BwelgFBllCdeC0ykfTI860w+5PToha
E/r6729t23eMid8X1N8+m0ns1RY1k+0nSnbIY0PtOS1NGAugAPsE5H9ltRjTmvyNVqXYVsMwyv71
m2wyIpND5AQHoKmMh6hqYe8hlbus/bo3cY3xXAB7njh3agbLLF4eOXw+eQmiVVFfh/cU96TQlnDo
AKbctmbgXeTfY2/cfvkboFHsNvcOCor8B1w3SUTLMU0lLPg3Mz1C8Ntl+cUKC/r4WlrMeUclnq/J
iEVHp8ubmYXiVrRZwo+II6/SBkuC2bfAIqQaT5GT+v9AqH7yhcdDpbt/e+68bGY53ocYiwANnQxA
6a8TteQtJnxFYkhU47Ng6hf9sqR8BRHYERm271HjaI/4KaJFpZX5ZB4/t3Fzjo+qj1DTxccQ+9xZ
Wy4IlD2dNxj4optkQmOzxx1Ct48ZAEzAE9obboc9aBmeryJ0dZ79vI4xw0kn2RIZV4/lZVHeKin7
f/CUcv98DN0Mjn1VPv7Mpj4R0mPEk4O+J5YlAUB8qiFhTRtAQ8ofNX4TLt0yGXJSK1AOtddnsxIX
im9rHgZ78FuqiGr3uKIgITzJoei4Xx+5XAa9KgfgVKGTOZ58K+4effL8hlkNyNvDHDTAEx1lmoIC
yMdUlTM2KPtDNIQ7RU+c77iWeUHsq7twwTKjYSKO/JqAaFYq0MV0NYzaEea+XzVrBD2Hz8sDFoSE
61DAphmdOfWHuuVriN5z4BEFOXRJ+4gLVkbo2TVhg/JvH44ycrOm56Fj8yx3sfjaG/eINFfk7Pq3
oWvSWsC5hEEf5LPMFAfdgSuBev6Y+vZ0YKGh3jCKslns9Ps3w1PUjY5iIH46T1w3WUITAzFJvW6R
rQlI0bednuPf9cw0Q0cQInob8/8iw2q6B0oWTHSJApZiDlhLI/25G/XrhD506hmLrx7RK/tfzYao
wA7s59Qq5wSGjv0Y3/OdyVKGIXTY/zECvNd7+Gpzyh3NeihwjUyiTiN8970UmzfCMMewpePWmGLy
ouBhMJpJgmYjE6i17XFOCnN+GyATmZPiJZsJMiOJickcZ0tFOuuBl4llHrNJTllQLehknJYAxg36
ixaKCt6u4IclUhSLJL2z+RCKmVXHdfeyPTxpJFeAPijPHDqyNWZ5CtqEprWz0/vJuLPrW2FeIz0F
63MLvG/sqexbfPqHUWiIYXIy8LGL3UPPEQdiA29stWdZg6hVYUhmbL/xZA0jhKRzj969uzvk4rGp
PPr1STi5Dt73zW6iK+St41Agly1aS8lLtIL6sXXXYa/LPomcTC9KVNEkjUi3XezwzuvfKbxDiEOC
P0VBd7iP6yQryAffBkRfHSRfMHOJVcq8l9mzbxu8NZtL/RzYgFChQ9p8/9039T5x16Xw1oyEb8db
JXKn0UbZX98k+MBo6znS1IDDwgZ0r2Ub8yoJXG8FuLeWbSSmpZOkZd7nj4mBHImTwjQEalRbMAsc
HN1nCJjuTPkhrtuv3p622MFI3/iDsfjZrJ8hVG23xWKFB5R1q+zoVUSq6HfNukFP3WoT8Cg4AlCv
CKwYkLstlPb24Wc9bau76vNU2yNwQsM7DCS72qwzHDVSvbjDnyJO7r5XQob2dqetBSs+e8tzISOz
UyZ7DNdUUXO2jABVUvT2DsECbX6myG32IG624Htu7qp6Hlay2olVW5CwC9q7hS00mhxBR8K9Gs5Z
XbLDoXa2dUwh2AZMVum+YDO/k24+D8oxOOW1wI/fEcv2BecuArckwlvODd8w/ekJ86tAknJabl2c
9soY1IuiHQ5o0Xhs/YAAcvYWnDZSD1qeqeITpjiQOGI1rgs9lB3pgsb9Z4FvL453CIIEyi/lM1fa
rvqSiAolJFDZVJlppq7rPMlp03Ox4/ATWBXunJSMNQokUdsQPMCstBKYChR4yNMD3lkjq7Y7MGTr
dXQ7LFlXOBE4kbq/8pEQtzNLT31VeG6HRdzOZYW8PihOL0XKg1fTOmeHREaEGCzURqggHzvbM0NP
rMkW7fqowrixiSmrtVtyuseAO+4ETSGUeAoMiBCZvmWXv+HN1eVjbod0sm9uQzPaXMiQsXWJKz0P
kBzf0N9FO4cQ/coI4m0eFX3uZOOWZdXHf1DOzcsRAb7GV0g1prMD0CXDrysw/eLzT/WegPrJU33B
WE2GmBx32sPoQe1T2JpCSm+Qb6sKzFKhQXlpQuVjVKupL0nU/YJcO/xllej5t9TfrLzrXt+IT9lf
rstd/ZK7vsQz6uImi/S3g+xdtfBzxua2jEr+Vzy1fbnPA4vEcFTD5OvXmyNkzEFr2yvwfsLc0ypi
7to4EFvrOhjodMsnplPY9hq3wGNhoD2KVGi6SqbTPatnMpY/S9BTR5PMEyZajMg+ZWRb+DYPSoMK
xXL4ILxFWMoiS3P2JvkvUH46D8FrgutO0+TdH9US635wKEOuBZfeM2OcJGv8UCawnnYCdC67NmNk
8VDgdbdUU0mTpcYgHv3uRs02MmZS6itSm/MWz0EdXcqu3a5HVlOlvv/vF6p9i4MEC8xUcEQP8xfz
juUTfRMZIOKIyxs9QTaiJOq6B8QJrheGXJjrVfB8jPKGfhcXgQW1CTGy1Ew0djR54JQqV1v23x2a
GMLmfpZn04FhdStzk4TfSw9d0FlTL0KAtESsCQIlmXCEaxyymg/mubuRfIwzWly4bM4Y7rxpzzBF
DISmapeXyQpNh5RmA+wvpbPkxesS6+lV1aXn9vD+2gR59nJoaY0UATc+pZKWfbzp4BHTZMMrhSXg
nFmF4P90lSbY4KTX09cutLewclvet5/VUGfucCZsSdaPDpZDdeoKnAaL+73K2jVpAI6EVRt/lP6D
yNKtbAFH1nWowZ0EH9y+GvKBbae7d38T6ImM6jcJWjiZTtTBBBKFjZX/Y6QgTxz2OSWcx0MihUL7
x04ORQNzi9w90K4necMJdAhU2kggMA5OlhNCiPpJZzBKB7CY7jjfP48uVNR8IKZpDjwSYQdIexsn
Swl8aiTwZa/aeD317EPHW9GfwOyP8Dz17f0BU2OyzHnzNVyxnAthzZqIy1kYMSaVWaYzPB8ENkCv
SPMLbFFTz2ijYGvACOCCz2M0L8GomnkE7RQcgwUrOgqhipD4c8V+Ih9/5aviL2f5qkgFyAGM1WMC
NTJMKwEv5JAFWyQdvcDLvsSYqTy7Y01QoPeC0sO0wxM0EeYT3y69M3ATtp22YB5yMP+PH12jwq/A
/m8SsK9HbVEaI1TQqtUJBQAI3pH3GbNz0XSbcp2m4H/uzI5Wx5uzK3z88z5yhPHR2Vc2RjOPWao5
NhJylsOTZMQxwRDK10LNrbVu9HpYqMCCtmMC+w8Rs6Y7Fv5Rje3/I1EHTkcpLYEXKF1SxzvgqGWF
d7t3qoBM+yhlJosJ4rmxCY0sBJnPa6cyBpxQPsZFKQZ0Ts2BAryulseSyLV+Dv5uVD+4FsGohBf7
ptKyVIzy5/PWZGpOWGHtWYdaV287XHXuOGRwq4yWo+AKvKNsw9qmR2LYVzzc9Y+FALl82szidNMj
Yz1qsgz2YHnXLMXE7M9k9iSKFJ2JY5J/zZqBpBQNMLVVFebfXvDBOUyFu/bHj3OKKVlsHjvKdoQO
RUveSFCCv7e4ZksJbOKP8JLn9dP9F3FFI77qGuj1WOxsZQ16z9bTPRlpEMKq7K2ZvcJV/V7eBvyS
GGgL5C8xTs3610yBUimEB+sLAVkYJIDeqVuodXMV/Kc0Lxv+oBzYLz2rHiztsWclcmF6XHbWYIrx
M2iSTv4wqw7ublP5l+xXs6uzzB03MR7QUXvtdKFsJIRtcXetCgGY4qf5qr1q41p1qQHoFxoazNVh
7YPxnZGWG9WuW5UG6YQmi++h37HBY9Y480cqlfpvEE/A1GEKVIDM5GGQN8kfFAkvn3dVHm0QNuqs
IWFwfiXBGR1In6d6OzDxZ7erejkZTYgf567VevGzIwcRSDMewJheWsMrkhY0KEHjJEVkwxS4eBwm
dplvE4Y3mEYHbiLUxdJVZuz6kjWHEpYEXQefM5KnRii7zOW+NhO2PmbdbCQ3jYt9vwgGWqwwELQr
UCowsNNCoDo0yZbPfA31/X8/t1+qWzp4icgr+qClbOrYQbxq+cinng0Va59KjRxW8JUUN1D+u1dS
/OqGhK+sBAbIwU2PWlPpXev/tIuTB32HTe4iagqh95qYShfuqOAa23vZVdeywxN/yNbRGw+JPXm4
+NYsDpjDcfGFRmVYwy6JTu93RF2iMSFRnseymHqiW///h/FJQQk6ycipKSkKjwaGhKd0qiQ4PrDh
dKTZenMXlrqtDRWT4EJvrbGgy/G1h9khELLeFDC3c+t4FvFDkbLMKfH0E/MS12IDAWOkkSqymV9l
7MuydnvqP5Mq3CsSEP3hgtNPy+UoGFbLg/CDoxh2wyIIuXUu3UO6a2fIp4MaAggS/kAJsa4sZRvw
0DIno2Joaw40Yt7eRf1UcQvMURkJLNh2sXIYQ3RLK90Qs9VaNTSJgNHQ726tIzVHCRZUFoGKedrB
etjVSAtFlUm/UzwpL4A0HRqVJAfquQN85kLbXEeV8ss8vZjfrLH0AW9Lr//d3OEothP7zcHKTm1T
7x6G5mNgs+4K0Ahrxxbe7xJ8FGFlHg4TWPBfWVjSGh1ElPe1z78rsSXpPNsjxGJ/Ejhx5FeNnpEK
gPMFn1PAEt4boUbWn4fDBz1iD8BmozCuFFswa/4rrnxyaZKrLb7k618wxUCpz8qlaKC+zsDkYvc+
3/PHyWRQp+VDpw33CxCbWy0l91fr/ZjN9QaywcFuJEAL+i8hzrQde9usf0YpSryCdIhJ6tOmTsT6
EP8W8HlBQG6O4GkU20vao8p4RY5HC2LGWuhL0IAkwqdgHS0fFVJGQN0XTjB2vEYbG7RutiGiOZrS
2PLHmmlhGz7di7NmCW5H6yZ1LqTgO6WwdPUGQOWsGSR98uSAZsS4ZZdRjnNzKby5gCXVr33YgOBn
zbX+A6AiryZVSLkmj5MhuKiBZex6HGY/4nT0nJqC+baXX9v7hbhDaj0AoeDzZ1KaK5F6sZ3a+huU
HqdpnSb12x5yFvZ3V4YQpEkH30wRFECMFhl8xqVD9wJzPrs/QABdaGFyCWl/6VHNrA3RfecSNpH1
EgBp3oQ6yodFtJtOILJNA+3QquxYrsjIsXxsmsnAnlIgpV8SmjY7XPUhYkfCmbVVruqNUTLSAz21
rQ7UUq57gcGubrH9Nr6eF22fA08PvH/vXUGfSczy3tU/p4guDf4fd1Ja7hV05qmSnqUbqizuYZPb
zi6cLHUxFJnKv4iuCwvwQWVgilYvSX2hnhhwrtamxvhzJfIKb4qav64sbZwpgF7+SOZvFQC6McY7
SnM15B3IMcK1FqHeE8S7KzvzQgP4RVDYS7w+fUV9RRx7ieQaoWetYST/+iSEVHMy8wXK2V7m1wiy
3zYsoIL1eMBDMFUh/GxE9nbwoZsqypLFPAgVWQ0ul5lXzUo2yc/W2OX37MBmoND78QAaROXejLwT
p/ST99aba1zWZmORsp6OYqhS88bEYt+eLz4MX0kDGa11aMz8RdvQyiP7jvz8Cu+IcTjRhpGuCX0U
l6174//1xxbpJQSnKmXfo2npfF8hQSRY1vSij55XzPo3xd093toiN51f+bBBByINBD7vn3j2aQVb
BzU4uX50UtenS9UiGvaoBLYKLpR9EXAHQw5R61gBbNBkKMjblgoZILVDpZ8ruLyxqj5X7O1V663+
6oZ5ztFS+R9wvN60tMAojhICwvz5TFtKdrNNY7uMnEofRIHAwpnG9bo5TZpu9gEw+Ab5bBrKXSrj
nlr2GOLuveBrhb3ZGwiccLexkHGAr4bZusMPEMsuRlJI3uZAZyrgYcGQ7Pl/G4EBdluNjFIC6IOt
izBve0apySO1Knu9wKzTdkGAywC9JcfdFFgT+uygNGKqajLkB1EY7c9rasNuTr/sqVcbXbCNBgux
q74MTz+11ACTtK7aiEmPDGap8yF4EGwJmb++8Tzih6d+mK0TBH16H20AFgOMBQ/yqGKGJnQeeYGl
1iwE652+KgUp9rHyXSNE1WbUVcEuRBuNpuTK7XPAFy4IaevPXylmyr0OrIAicnTumOUP3nVPEoca
GqrNliT1CIJ6uDEhijOuf9vKeIN2LhecdHeWydjIiqoRN0ZJsjBjsk4ndBj3KYdJ/+6AF/DycZRm
tsMSHt1F/aIA2HbcL2ngf3+eLJbbTEn6R4wTwAvkBQaibeS/ulXNkwcOoXNG3NuVceWL2QNejnsw
W/3ww3AKKwVpPlmPhny9+PObIZUOuAXGCT9sW1NQGhRMIZ9BD0g1NUavFTrw0AvgXXTwMBQBqLZY
feIA27iiEbVKcxqSkfMBKXIp5xgLQxBE7T6YaoLAQmAIC0qG88iyeKeB9gOxGlPComHZgtDKfIBn
teXwFBUzz9wTsa2hX82yVL4nsHqrMD5aqqfd3FmYiiRQZi4AerQPgasGSgJ5vKBZhmQfzChhuZr1
x3gLHWpCj6NNt29TY7wzr4zSnm49qfok4DOJbr9PDXGh7gkqQyxIRkKBUurFRRUqjY00MlkFxMJd
oMUQclcqxhEfV+5vVPrc6FguB53VLZM5dsk1HfUuNbK9gPXtWSoDva9UPtfEN7rysLJUdSgjrUAO
N/wlEe2N2ahzo0uM5iPSVOPFIQFP/K0Rql/CnRqfsDKijHUD3WvjrcfAnYKqK0jhQCKOsVyDqSd4
gPvyoEJxnSfwlmoHrnXK2UBiMShy0+7vr/TXQEfqmO7993tjtvCcdHjVcp5AjfjRUF06Oii7jVSn
MNNcJQPgyXzAFD9LpSsD62zTKqEuXQmEAIe6nIlbskLIczbE1Wf0gPucX+2MIDKXJJPSWpdx9Cnp
smyFx84B0S/CN/rfy63AujBC2VcvIaKmAjuR0C8Z9LzjRgrc8Itl0fu3PQ4ZiEzdQ9uvxQZLnEWR
O8WYQzB290jvxW5K82V8UOqp92ddGT1etXuP6TQ67C8KDgn/VifGf+m/D+eLulk1ALDxxqg06eHY
LIveVoVTK8zrp6hNCDe77ROneiVo2xjQraFd1m2oRwvnU++I8mJkX7pVcnDutbh7klM9UKOItTL1
NqYe0qwNsn9wrgBpOnSqVrI1qssj5nen/WZ4VS7w+RCFyM9CiYnP8n4cqfXEud8t3gaCUbfvbXCF
MEd+TNJOCh6KAbvoJ4m/GvH7w/gpHJItG8dj/sjgMYyXmNebVnIGM/i1dB4vUE7O/Q6tHizK0R57
B/ggnk4O/FTA3eDnoUzJ+v8R787ofj8jtkVjOOqJr7gLv3jzm88Nys5HnEJEgbl9lS96kx6uiZaO
d9wYnbH5BfIBHvTb2fk+svdTmW5JBJYKbJ1kti9qpu0ESuT7N3Neag49UL/1IwrqBYwrhTzrn53o
7ZPQjxiDgnCX9N/G+4EbEf8JDCvEaP3dew12yxUQ29dYrUXFdxeDI730VqUk+lnJ6i0QITnBtDzE
xNnhTEuB0XEi6N3jOwmA5m0nbV5mlrT1HV2IEWjY+vblOe//AlCamKK/u0DSBFYrmEgANxzfreoh
N/nzYo8vAme5yJ5kLz8kDdoxP7s7fr/zf9NH0Y9rTh9CFUX8RCphzLlFs9SWjsuK20di80uyzM5P
7NDbqLWYiAoNpvRazF9LOuX2fsBAaYYXb89D5zjldx+QDqD0FwPhkcoB3VJHOhBtqKMYkO0jdBxN
2+jwx0bFumUz7lQjOGlH2VdfR6uJLKi3wWGrwW0OAvzKRUFb2Qb4Rgfh0NEa5Y7B4nXxGWJoMoIf
fhMlawBInt4gSFBCAE36V3ih6MZc+2blEIx0unmHvyQpOBiXoAHm2uNlBS9VGQjHXRnz2AuWkcZK
CYuTudVMKB2fUAgHGYm8nEXQZ5ZNjuk5aKeIwF49cMKs8+fZ1U/qxAfZKAgoVrGbWaLP34MA52cP
bxXktrhEDHGoFS2UjQmxmuRb109ASw3Nu4LKAogK8f1NWeY5KwfAgUWrVVKVlxTFBk4jo1uVw+tu
1pUwMwE/FH1zaTZLh9PIz2gWLXIbRTU4FtgBQ0TeCg8MYjUWWVetYIlz5z1wxUJH+nRxSgVMKZa8
PeoDtXFXlwerm+RlemmJNyOse/Sqh3ILkM+M1CXGyoEFHtm6DEHqmILUB+Cs/yteXvdBa41ZInrk
AlS2ClfquqBRFplF+TA6E7RTnzAqeIxkDCoJN2Wb40TDHm2s0cS4ziMyF9Q/ESUVT411NdYgbnwM
I8VV4Ipml6J551lHEzrDiBRYa54kEcKsalES+Wn0JQfMoQIkaVXw0+m5nMEIu1oGqEkri0T345XP
oxwZZhHBD1MO/0t/nNuyPct4575gRVtOl5GbsOUkjFPryOFR9oLRyPOv8Y70wnkaQELwu4KnFmnl
2vwUCwaIbf0UVPvKIGZ9Zfs5RvZEeO1LglS7rwRGyAk4rZxZ0KTr1/LP2bV8g4IlAqrhtW+M1f5a
JVnqleGYk84cXqsjh8Lgn+6wDLwnrPJTjkvKpSBQ0dBTQ3g4BnUzGBb1LA6k9SROXv2dSt+kWakm
vVrsZ55zQbBQ+U8R2RXEHhuV5XSj1iPkokFNebAI+2136R2ltneyMvKvET+7KZSRiWfEhHoNX6CR
XfZSKg4p2gcozueoDRMSKhc05R3LwSXl55BPI81uvJfuwyukXW2U7SQy08AfBFR7CTCUVmXd3GaE
MgNhkpv2LrAjgfzGSbPoOBGVys96U3TqeyFkxSBVBz8xo7h7HDOEf760jIKKvdHhCt7gNZC+c9m4
VUVXdOq9xfXLEm6QOv5rJliT5puGDj4bySDjxXGPdh0ascqRiFzznb8itwyrfgztgmKk/OxlItEn
FNgt9FEW9do084ikeMBA+cyhGAaX+83fQGtspcvmAh6UmGtF9e9ZFbKBzi23ytuTrO/17tPXd9k5
SBFE/Wu19e0x8DWFbuCjuagBZk97r1gJv6A6VOUu9VcTTQyRyB0SBxYYUsfwacVp4wbkaXxOb/fz
U57jdVCLCGVtU0XHMpjuabBfVehjFpXkHhuJbVnv/xUU5ff7BILazK8+CG4V9OGodevNZdKocbmZ
TX+/kiaO7V46/Ag4lwXRWBDd7uh3cFChf9A05sJuZbE3ygU7xFHeBWB/DSFMjfedKc4545On0CJ9
PPbZ8leYiJGUBmsuuoc2AFKSyFSxhorS4Em/Izn7jkP2YDgAIYQSb1INlvy0FWEvUCmdPxdJvW4p
iXox+K6x1ZOAoJ9UcX9TfbymhUn6XzZTms1Xgdz6qkeCYVqxPyEOTeIyw+m1B0XVyr6gayXZfPPz
fTsvYi8ZFlRG2Lm+KrsaOBg/VRppRKlqQ8aE5AUQWpDgDC5KDFHx5Md6oNmunwyykQY3VG3NQZXf
cHKupVrmtyXGPAUvUKVt+nrbvwT2f/OnMLDQwwBmvqyJcz4oLaaj9aqs5KwrYSzFWqQjGiZgNhZh
cF2Tf/ZIQtX4doo84Oww82waBxVjettx6kN9HKkPTWhSVYdXs38fZEYoTgvOWDymyjCFxFiUnvuZ
jS7EalowfwWXH8GWTba5rjXTAprBuMG01knUFDJjhra6oL3CeRcBh+psF1pZMXFQTCQg3H/BvU1T
OWHb8vD2wq+lbm3E/N/9RIjmZ2FKzHqjPuud48ayVVXuGumEX0O1IbtFnsaLGR9qV86jzK67mnOB
tcRIIrQVdbk9BcLejz78RNQF+frx2kD8w+SwNhsMon8OrB3uj1kYtoX8UZpJYPN7Bx+Oh/z2hzX2
ZBWkbvT/lWOqEz/NWnQHFgSCHcS3fL66zhzZ2TjR5NeoDnj9x9cY3pH9iJLxp+RYeYnTpArriTSt
uuhVZhzTUReDTOhleHwDaZsbwRHHKnSb3z0IJn0Eg2dB6y7SBoUmkgwznx0r9ybiYH/6LlM9uE0P
HqLY38gp6htRrt8JABvG0DWCZEsqeockii1Nzq5HbJavQG06sG04kr5NyY5g83MXC8cJ4+eh9nji
VYj4EdWC1nTF5RRAhbfdAQbAQoeFAmM0S905I8HaEEQh+/l8+NjVe/+2PH2xxXcbrZ9Xjsf1U5yU
k3xgoZ3BHQ/F5EZvoqjcFUBBbZzcfkMMkp1OQvlEMYAh6F30vg7R72G1vD/QKpLpZUXcWQ2qIMuv
0YDJFLFOHUMmum72bNDy25W0pci3axfIDy2tuVvuCKIqs8zWOcsL5dNC7UY27Loc6Qkp+MN5xalI
8Vr523ZExL7bLk/lWlYIrHJZwyE6gATqBqXy6wwuYjod1ivkex7DW5Ed9ycIW45TE2wkZsLKXxiB
QjnIdh+JpQCYzJc3kSWbQtluO0tqzf7FwCV+0GJib6obzpjejF5n+DskcO4veSbmZJt33vtgGSUm
dlAo4j6rqH2aCo1cdW7lFmwwsVF8lBUMt6gJCMbX/4zQ6S6pMKc2gc15CuBgKf8g5uuiythHl87+
x7E8W7MIErUqOJPNUBtCHQyWbJJ9n57PUUzVAmHFZfcBEc6ISyQKeFnCs2JAEX3TbhHKXk5EUrvQ
PcxBCgr6aH6JXfnQ3hdn2vuJs5o/tkREuXq8KylsWNejPcLk5+oMIJm3f4aMiQxZE3nSU4QNsXiq
WAItgE+rXKb6hBym/SQvVgEra2wBRxtgYzUkCTlL89JsF72SPoTL2mbX5Zs1a1dWIOOzgq5qD1fv
6tS/WVszsQkQhte/JZ2cDgi7zyMqpqJo44NwQnqGkvHo7UCzrcXnB4arRZSMP9f2jqJ5IlyARvRV
/C7vgzv+MQ2ZBKAkRY3q6CeLwZTe1bZA9YAUmdChhTijoQvv6x8cD+YXjbtEFLNdAwsL5m0qFua/
BUV23NP/Rdc/r+oAuseIal33xcIr8Do3QmX34jTiZNg+wN/y5PmOAn1uIoFZG5sdU+qr+BP4Sh3z
OzVkZYGNwXqb99Fgoc76TIcdUu1VLnsJPUx3e1UZcdVURs18MwhUvchA6uSePih5X0wBn/IlpE4a
MVIYekXWo9ZG+ksoo0nFzZ6iKB+N7pKJx6MPwA9WaVMQti4iaH5xJOtaHHkxhT3ml0wR7cqPxsh5
tZnDlRHXvJBC8zlk4PytzH9hqPhk+XVpx587oyR3LlspKTfyIOG5MarA36v5AHEk7v8OiVp3Q3XU
LJm4TaMfVYFY0HeMt9Ic0Vg23rb9BBJ0TJo/eLA3X+oVMHI2uYQBm//hFmODaGhslU17Pw+BIC5J
Yxgrs8wbLJIxwOSXfVZCVS50v1ijoGIwhkokXMDc26Rw6KJEuC36nCp4v2gM1LPK8F/pJ8WU5qCf
m8pQ0qdU/YT3yNM1raKTVdoPmCgrVIJR2FU2z/b2D1aDlprtcYA+giBOdKujY7lXOU5FPEw8FQYW
NjcbGfXwt1nc28NN6YSz+Qc5D3qgJ0r9majkicxKNgzGgn4D6n5sf0apAZWkt/rwpDgm69/41Wj1
yeceJ19tiOoYXWlYU2odDPuEf3VIhxG++X5vPJFcFDjmDSIvSe6HAJgVtGU8C/6lVuK1iyKFHqkc
HFusqdraPuBmpNSb7ofdxqd8GtO/qiPUGb//k1Y9tKQk6Sk2D8n/5sOythbYWwmnauj4e2CdAu2e
K/u09mAvWAq3A3JAu6n8QiKqC9H68YMt3ehDqlFYEVtZomz3ZblZifwQa2tIBhCKYHgy1ZSKHHY6
3D6sZ0zdUbHT9OeJJ0wyCxGfCYTuxRQPwcDLWq9ud3BxglI52PQu82qusuEduTRBE2ugaSqk3/04
fdBZ80ikTsxZgoeHFDNwbx20eorXX70d7a1iPKogwEfs5opkoi5tFXzCRhjvg8lcPSx5FbHZPM0x
WE8K4WvFgIWknLjfCZa6u7+p2e+I2Esb3IZbIM2GIcwPNpXhwlY3TknpjtvcLBcYB+rSin8ndbkD
E5hWVb1vWJLVSkDPQ/k8UsZRhXuolJGJJMrhslpprYOWiM4XNmM7JFmsoJek6ca3vUr/od1weCav
Bsyd9AqQjqBBHBB8F7mlAh9mrA0iDZX6tQasKHsJvK8JOiNAR25fnI9lAUNpeYvCJ3yKlDTArxyQ
3et9z+zx8Do/SpTJSt4czh/FCZHrFKm6j1fZR262w6HySLqCzDMUt/69k/ZgyGOozO0KuyafN0k3
3h403OmVVkRKIy7PwzgMqOg0+ZXTLGuL82F87Q8GpFl6YqMr6QcomJo6QRpKwyxihU5Z0v4lFbRj
CYr4L9rFLJWkkIdtQdlYSURU1I5Ar2u7ckzSGiEwEeWD9y3fSbxrhYo+W6m/ZF3WAD9nfACs4aLZ
4n72/42ti6FUgHWaoGYRY+fF8+/OQMLG0kVvVDkVfC03XPsFKkxk9LOk/zaiCmA9WC2dqf/FqnKa
bOX87JtTZS8XRghkQ2J4Jf5GsF6sAbo7sJLvn7a8vAhbkunsY8RAO3OyBDEebTirWH5TB0yomf82
oJt3JM1E8TtAuvLREIJOkgGbLZVud3BUa4/p5GiGa/7H9h2SGRrlmBSJL7bmbTOWFRs/mAaP3wGr
alUXmSWKJKhnyhA73Mxj7R1QWxQtCfiDOeeYAmyEfXwv9cn8AWkO6SvuTbEa4G60w3puvHmsfDj0
cT6cTn0ulhgVRBkgxd0oMqQqak2Z7FzSW32IfkULLT0IECYFV6zWXqcDMcPOwlF7gzgUqn0vik0V
VSRp+bQKwtoxPERl01rOlX0BWIXc646L9T2olMVrWvX3UEU+DQNfiCgl323j8nS0ziDxXnEfX/Ay
59woxsmOTqqIy3PcbL7nkaXbquidmWU7rrkm/4XY9uQsOjqltephakhT6VSGsaOUnqjLkTEUXcSf
+KDkRwPnxdDvF5ji2UzTY+ZgTeOK9RkW4SoLxknPU6J8bVqrImfj2Q9ELqHhPQeIPzz6Yoq950K2
HJxmWQB0Vr9wK1LhULM7pOt1w4BMe4W2czhMYurEK9nR6BMYhJ33hDlD+lamyUcBATkXNMZZGItN
uIis9LTeeDTTnNUb8UQEapgtADtPBaImLf94X+QVHbAcpeJop4SyeKUGk7lIqkEXRKxDz2zJEA0M
0klJ2Vb+rbGTr5Ih/Ep55DqRon8K71331Yc3HInzcYbg7yq5dP0b9A8GgmqDrDjJjtyXfA++dKET
1rK7sWaedVBl2lx4jD4NbKAZXksK1zcmGc3Mzae51KN7ZFjY84O5G4ayhkGyJav3c9k0I8LWppQH
+iiIULqVQ2sNNg+ZVoeatuEK1kAIou7p1LxVLVtZHuEPz/xWNVjD2gDwy+MF6AAMifrdwYnzAQRK
Rap0aRNL9Qw8YFOlAPTyE/bJss+zG6GeEvy8sgbAi6SwYueMLKR/we/Brr8dEud5mxceFFWS0Lsr
3DwTU1Vp3YgRz0zoFO2ktam8272Et9QRU26eN7aAmLuiJQfzJ4aIqVG0MustY+yg4HwtrSt/5PN3
YYbpiWNLbn1oD5RfW+QBmuIZJjdE/kizB0tn3b0DvkgvQOqa63jTyc6YF/qIVI5v1grTT2ousQI9
Jd3T3Z2NycpBdedCHGOxVYv+Qnmy0XDkfdL2GS0o9vFyYDeX8LLuZav9TYfRRcq7Y2T1cHU5hJM7
kkn+bQzFsCG0DcoUGA6ZBdR8OlLoFJ95fWZnEix6jagi3J5KS+2O8KpwMfVIogbaUZIvJ/YgDN3Q
2MzOyeuq/SuP1Miua48DHQFdoA3ZdY4tL/QeOjDsUGdV4Vr1Y1mSmFEfBg3xP/3U7IEO4gIKzyNK
ZMpo4uj7IY8iSxTS564XRtsz4/F2wfujLcmU8AKoenFK6c7RKwS3pECkJzr5AuenX8lnY/uwG2eT
v9hA7yOT6Z9OmdXE1HaAThibIgzBSd/oSne5BJbsfqTFDz012p/9D35hK02IxAPIPrrYX1OI5JnA
3bfujelMoVRIkC62b/+T2y4JuVpkArAI6CfNXPFZJ+/5uVqNmKd8l1Dhpjsvvgom3xmRccCvzhAM
vfLDghbmPDH4iFneMMk6Be0BrgrTEl9xV2CDHOK1SnHT1XlhY0h5trD62SetZhNY8THqVXN9HCDM
LSwNsAuOG6F+imZ6ZnGEY/SUeemr8md/jIGn+k9Ip1GJ36GNcTaseu+aB5VLKp1uZqRMhSBjDk8Y
Mq5kxILEdTPnct/iQSYlSg2Gef15Q6+KBu3P75sjpr+RHKcsd4xyyGV7yzHh/H6qemmx82pe0EKF
GjEgv772xbHkwOHLHv6KvohNh2VvwBXpBYDokMsXpzfuNu5XQs0a1tjPZFRyTrVAH+6rI4qmml+k
sea4kOAP8b7v72dZkMb5MD+IacisRxLVhit/iwklfqFp15oR4CB9zM1+hfrGw9KWKFiBg1hP7WlD
BhSUMmd/4TjjaRlxbs5wSE+1ynJKGP2tFIlGEvc7ITrY1L/00TsLLLvmbNl0GAIRAi9O+xB3jSPa
z5Qh2TDBi8WAYRsXNheHXvgjG3kL/35UxrqcgQzvweblDBT+opGiPPW5FT9fe67wH2xaQJQWZgM6
ojahChX3UTWBjpLXCwb+qP0aJ1ZrhcXdVyGEVgs3eJwJYwc4LPVhz/R+5i/I931ap7HnxyC5DAk5
B2geqgw2otWE6HDDHm971HiTGoKIdp/+if1dlpjbpmtIsMegvGU0O3d2OD4nS6pHlZYN+EZNjKoC
20V+wdOjyzdxo1l5XFaUYJ25ad1wyXjSPEdRuOEaqCt1ufsk56VFJCjHKp8CYItlSTfnaXtOlxDe
3xRs4A4rzRIB8z2n73vuQqEJqi9/uNmuhHgRoLoEtiYL90i+BxD0GOUPijld36xoYmjzug9g+YVS
I35dI3Rtr9KyG5rxjXRLCBNYCq7d/4jfQCDvzdE3OWp93XNtewyVZ/CM4twEThwV9DLlNBDfCKqf
7M5Iafv39Dq6Hvcp4mZMBNvyJNCa06dcqgLdkhJ4YHwX3o7Ne+UsNr3jxSZwV7P3Ss68kbd9/x9c
2Ik/+QG0XoTIb5V9PjsxvMEV4A1Wnbvdi38T7aGQEVePPQD8MDbt6kC4Q7IBvnnm1DawL6dQF65I
XN/e6lMY0IW+xK9HJtu3Q84i2/Q5Tk9RGCXip0CK/24s4xAryT/yiqkdAJoVXuZ4KWbcZviKvFHb
u0sGgDGNEtmux8aUMkFAGAfVWBIfU1ZM/K76sJXgWaPtzHfa6ES5Y41sU93Cq/ooM37t02ysJr3k
BsWEjjQ903nrI1IIkvMfUaPNfDwoAeS6E5OLWZdsWRCLnPJZcaO74GO2z9uIa2XZ4QeoOBvbVnHS
trMt43wC/m0LNu5HVKifU0mYRrPK0JurPNihSYztdJ4MnNDS5d4ratKeaqp/Nsar+pr85OFcAeV4
qp+yTNk1hhiysF9FfjALaerHit1ol6ZkxhNUblrf3P1LiwlHE5jaEUlASnKG+WxVt8UoOiPchFFs
6kvI/cEytzUFBk5EsAx8gjZgc0/5kiSId0TE2g+KWjTlBWOyd+bogjYXvyDjlS/t//BrZvN3Esjk
eCSKl2s7/xsPKteErkIgDqZru5JhvL9RaAB8NS4pYiVqjZBesj5xJH3m5XQ8PUvW8HDcpFZSVAkj
jMWzoEqy7sk9NopMJB6pznANFRZgXjTbf79leLB2OSYbGMHCeh89cuZzdQcfoSBcBsQZjxk7tQGG
rvl35cJ4TrQzv5GaQRXPwu2IwvXlYbxC5MWEps0jAQDf1bgG/vIe2BNJxWACHxxtocrn0vCtCG1o
V4RxEgo/4LkWkifG9eV7C9vlcCZHeWpQhfsQNfmFJGWkyJ2kT8IeM0SvFjw0eea7QM2fANvDWcjl
Evp2JsUmo5p7VN7QaDX6xsU+rFZwNzOn4/ObHY4Idjqeh+2ka9DDrujE8W/fnFM/2VjRYwxloMAn
ab2OzXQL0spjHs690GlYrsFW9M52/HHpAa+POXOW4uaXxOLEnIH9FplBWZVqj+iVot6BusUgsghk
Wh5ios78kokUQUscbRGQsWeo2+GpW7Oa9tOvkag59/nelN0H5Kt89XRiSxe3UavdqB8Bzuxukynr
7gnjjm2DQeLPfwEvTaZDoQTc4Kv0UZFIhrxrSlxR7ibCqG59mV/voqZofAtN2J+wA8fXseDb8sUL
PiK7D37QCioMjOUmV5njpRDz8/bHwFSW+aGwmbGsL3NQIOpD1y4Psmlj9lj6Bbel6ddBmwAT0qKS
4UMqwfCIO7kWZEp2cMhbo2UYJ7E/AnMAklxMFa9kT+pzqkf9wpF5c+0oeTuHmrIwfxi0sgiSEWxo
mB6Op0j7O/reDf3mD8egqXrTS4UnAvxgeeYRWWY+/u4NFbgs0Hh9OSjB2KT9/6ppI1wu5wMnSCxe
t7zXV+tmbBr+hs3WEo4Efrz0GxpRlpKrygEXjAKeT5rhlhaQKb268QOFj+q7NYrTV4ZPyq8FCPZR
4ez53h1uHZqu1PYQEJOsegnJaCekwa+xvtlNXJEtMrDX0Nv2ETvfwJOk7fvyv22Wy9QyNLPyFxKy
t8aIfhOPKCLXQsLkWsvRGE950LwpR83y+/PIJP2CKLelQ32C3bzsvKUgPnHwcJZZ/qFj5ZfEhF2B
IvkVPotzeLLO5K/JWGaJGGeYMLteXFIG/Gg18J7cZvrSBoMmy+vyG8cL7xM5RkRUCvjnu+FLvcEw
kRpJdKzKRPgQ42v1n9fWEp64kA1MfF+v2o+A80hlssViaq8G70sWHrDvgWKNXzF/lILHNRgBmiF8
o8gCv+cx2HlPL8BhPxrhw0HFudQ8FSlbguY1Wj0NoEC1QTLTd85jqj9OIsl152wmxrmcS29l0eyx
xKXcXi9Mp/7t6wSt588XJJdRwtl/MdgIppOAU3wSlhO2GSQnl5PeIo0Os6lkg9b1taYDMwvFXeY4
F304HJ3OopYsEFG3UEE2tM6NrjftmLmaAziT8xq9RRZbDMKzzh3sDqYRHZNG79c+JKQGeBQIfn4v
YOONhPCa2p6yvhOPJRNYEO29CSScAPPu0RNAh9G6lrEK7eMxAr0Pcc+KZz84k8Jzv0cIwAXRl28/
mRkppaxajMkE+T4c+rgnfsv8EiDJeGYdFDq6D9sK83ZLheM6m7clFgCwJHPAHzJd5o0rW27x5g7Y
UGfmQF8REOibryg0T5r9whOunf7jFR7CAIljNj5LvMXGQEMIQ+XbcgidGgLG4mMN3rQnfN3q+0DT
cJx1FudkSL5bzv5L2CL+MoOZpWtWQnT3Kvgm5vt+VI9n9FTiy3bNUbxjIAOGGT3zlYEJipWUeY7M
M/3ZbWW25YkbPUk/1iWICyuEK/xdg2CP6JPmTbKGaDMc1gabIDeeHAKDg4OfNzX0u/fwcp+9MFk3
uyS8knCoABsGUqqogAMW3wnIxB/I5X73MUddcjx7EmRV6iRTYV9Q00SLFhMlcSiNzERvxj+tUXhn
+ckVD5JSYBelwpMmLeRCtSi3RXR9ioamJRbD6ZQqy+FoUFKCJMGiziSKb6nIqdLSvpGNlcXuvob2
PoRd9QQVC+oPuZhrE6XwMkntSIAQrNRaiIDTWHF4Rdsu8n8oQyr2PBjnTioBQ7Q13QdFmdMqFmXI
GRJD2G3pJhcoB6XneYtzQ/83MOZlXxQMph73zl2WevFJShRZJP2l0bFL+gdO9/WPli9tNBkYqGxX
iP8Y8RSIrZELqaf+Eg+AhqcAUtOT0fXrNfS6zISUjsvrDpQkWPryuXHWu3Yi5frX1w8+8k6MT/nl
FTudJmzFPoBEJJ/6AF/ynjR8VtT3XYcE9YR04w0fmtfST3+dt6zN4MVkoaYQ8D+xjLcZFxmQ4ydB
cgNJ+hRrjmLTyRJkC/SrycB7v+nvLdSCztrbjEzDL6QCdmSqHYcSRZrbZs4QqTzzahCl02s7JHz5
ePYcc4M1TMJ3QLTCLJ2WzOqnUbCjrBitlZtdSA/1uKuW1Q5eFFMOeJMfhOvaIMD0tAzD7UwAIueU
hbHzKwpD1nqZvSqW//MXoPwC+mQ+1mnrKQCCDRvlos7hbIw4u/O/+UAKoaOvZ+f4SQOLQ4d8rd62
GCVfbb8gwks/wh1X/gwnW9BBnaPBuMdZqsHaklZ8SS55UBo3GGNaW4swk+6zTNYHtJjG2+zwE80t
p/9l66z04vuMkQtKXWDPm48Sp+ki4px0Bi3VPnuipT8XBRgeRYycKps/ieHi4SsjBtTvVSRErDJa
7vk9jIEIPOnHDNKtUcJnMxm2CkUZr3tOGL9wioUjLcbNgTHpk6u0G8n5u9BZqwrtV92zDZVWgxs/
/G5RsKafDmOJAylI3tB/ZGDF0xyyEtajmNgtZLVbP766nflnw1xPQPSUey0ODcBxbYA3I8ec3bxw
OJHg6FnW52zFr9bUmKNWIzQJ52LjqtV9lhIOscduuuKyr0vdqLGDtvZ0cIURl3meANsY5g4C1Ed6
59hoHhpZW7sKjw2uGtymMbcANMkKyJun1ovsw0aV1u0RLWb6CYNk26Hg/jN+I58R/Z8Hxp5P8Qvt
ZqKxb6pVRgxYq8AGTuO2SgAcGfEKnVb92Ax0pS1/ZTpkB+aD7hcnT9kzb0RtndTH4UIpO3j7bfdW
8rM+m/UBLXB4yf2mz21oYV/t81KfMxGk0Q9Rm3epdYyp9yH8M+rgrxNJL3xyDDNlla63wNjE9y4Q
2hpcDIjE598KE+5JLBvUYK4NO7uhxzeboFX0Bg3VIw5Supvb2CbLlFBcyouWY5xhX2feVLkGjQZE
oHScBBp4rXllHNUg5uJd8BpVSk+Orx2JnnMnpO/+DUogFjJwQAYaniWdvv4yBHZgJ2YBGgYRR6+m
jYlRV+T3750rAj3Q+lSD3s2IOKBClqBeRzLT5X7T1kpUhBoXz+7LUjgAmfeAhcV386wdCq78EDGh
eXI1gTD60QarLFKgWA6TTJ0zSczy2bPdPQtmhQLBozbepQuYZBGDwi0qGRv0OxW1Cuu9OgnWV/Hg
uZGOwTfkq5FD+Prpe0ZmVKAr/Fw8pLK68MCqC7o/lJWP1iwmZSnUFK8RtfA1J8Bu2FjE3zbw1PCC
skRUFbOds+gCTgO7LmC1O37oZUBUGkUH13IYjXpX6VuKH1W0hm0SAkpj2GdVCKLvqX4ai8aaKRg7
HngHjkAdJirpblpFpAUH3euyL2Y3aUTEKbK8F0o5yeiYPNpPtXlp/oNMdQaX+NyndQ5og09QCpLS
S1nRnO8HZ7hRy8n3gZa/42qD8HSFmml9fzdWAnNvdy980OYFY9HCof60wHhHR7P4qxsQ8DA8D6P9
b4kDxvSw4zgBHSQrXEn6onO2yysgsqkujxMERTJlpJH8c0WpSnWQP8KzNx7IOmi8LumLtjaAG2Dt
+FtpU2d5Vs5GqLz0OyFnDpk1AdkJnAT73rgF1537O6d+s1FwBJo0G/hRVQj6Pu2mE9MdSCxF5fVt
UB9a64Z/7EiB4OSfhU7w/59Vsr+karhXAdanlfD6tlpObw0l9GLKZOpkVutr9wPlixmRYiL2Pouh
Oh7mqYgX6Ts0CFNz2fgkR/m1wSLtnIjNgEjcNv5wQGZs1chLigDnEb8fb0xeEFA3Bilm4xVLsXSO
Ulvx9e8Nz8MISOfDInFTLLUIgtfPqPdKorFtM6P4hvhHgbabOVdsMv0P+UZ8uop2jRRAmKJZVlYn
wQeK6oJlF2+eEJpJwnjWZjINUqEaKuynF12blnHcpDkKcizCgsLdACO6nXI8fqo6/7sqcMgSdBQQ
4Sm/FHEmSzhYAITTkpucr04ZAEWy9USGDfyywr3SI12D+iTevvs00foV20lvJ6sqGdXDNe+03Cho
jLOiu/AIUtk43FBIU6o6iXmxeItrJtDWKtZ/mbvN1EeARBUxJiky8zJeQqkJNvYQxdy6BsW/216a
qSt3Obz87MKyNMxbW5nXPgGw127E3ZRcvp2GOgVMlw0elPGyTAC2qaXN4VCKO7xd7KZB1BB+xLNg
xDeyzS6gNB2FvUy7db18yeR/rWQ9ELHvXRMOy3Cq3cg1GL8yrZFHtroERh9paEAOJF7grZbZ6wTu
/LtSPi7lZC8LMwpqFDf8rWUwBJlFZrde/k9hA4oORDEIs58/SCzxGbJEn4nqpLGtNQd+4mjiDewC
WyQ1xsg2ilFGT9sgyxPhBXblEpzf6a3eOrH4P8G0F2t4P5Kmqlh/EzyKRTUMus4TmIyP1pv+JsV3
kFPMwLp9o4WLP5C5Cduf6GL+9YZ/tkBEBK1gOVomBusgoKBrVWHrt2azupKyqO31GQrPRe7iAbQr
IvxPWtmtIRfFGZLnd/hiW3UszT/e2Z/S8ISqqNH5hdWXEP4kMqQLzdk3kOwUtMF/UZASa9mS+iXM
h94DqZBH2uzDRxrAT2I6kWEawr23KH8aF6MnblkND3PoAdYysfrcyptkwUD4DsAym5ZgfrtbmTTi
s5ZhPdAS6B9V83U/FIFFH2f1whdMRohyeZmtYirAeIPBEgNykS5jqJi4OhCRm1gj51WcCZxjVB8X
l6NBjZMgx+M3GSdgi6w7zh+lLGWpcwP6e6tYQ9ay23rATLgbwX0Wmg/6X8WmduBjdaFqbGo4xce4
q+xPMshUxbKJcOBKnYs/s+aSXO2uY9pWxE2zZGEGVMU+K0tOeEAxMhi2tv0v+Uu8jYzlcTpU1JyT
lHMvByU8e2N3ncd0iaLHHweJe2nr7Kn9prVTUlxGf68VKTlkVHjZx7jem39Psv4viOLvnoMNHeYR
2OBhXLDexfvp20RJgkWNXXahncIp6GI4VJFjZt9KjBFoeGEcrQRYkjgVucqHDRt1DNWV5A+qvskl
mS4zhCDUzMiPj3k+iMXqxnpfInHtMVQoLft029GHNfqasVLAPSS1fJiLChW46Gjn1LgcCyCA80aL
5cqGedk55VzEKr9vuiG2Nd5p+Ha668dE+3M/srgVr7MWvZcA4xMpBP4XfeKE6LExRLJHjzG50oyl
rGrQ04B6FAWPanLJOD9fNQ8FCrLNPUfd9OaJD3gd2/QEVZsQTH1BaSuQZQ8wSMOLb6gCasmDs/vC
lQs2yktxrWd0pWz/ZjcyzQ+AUASG017r8MyKjhVFgh1Dm9TUpOrd1e8tEbuuO59mBxc8EZZAjB9M
+ymDP6g52bMOmtVrZPMda9cYnagiAKEQv1y3slx4JR2pvIKcXeC+JfRx8uRNeRIy1VEqMZS3UEoi
Yar2hOq1yO8lROyz+uouYdqK6flhdx0f14kG4F0r2hU08776L47xxaqzcx8onbdnplT+qPPIBJF+
K/3Un+d7rmjEpntDS7tbnfHNkkHmqw67vxWlRqVXbaNuZ1I7c3xCqkU3OhqCoJKa2pTBwz7uvdsr
24NImbs7PnkXIIwCvBym
`protect end_protected

