

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
CvmaYyJzAT4gGJRlCkE1yXt5Lv9gJbr2gC0wBzixkhI3TupXRLTg9s4Z9WVWp43QDkUuM3VRZjAj
RVnqESt3JA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
hHyS2uxRkJ6sHR79RwG8dxYfMwySDoNzo0ZpVSoiAp/93R212I5J1LxM+7EujDw/cO/x9djlyxbz
erzC6/tIqQ2nS2hUZANmmER9YkiA1RlXlIqDOWo8pOFHNj1c4jf7Zdq7OJMDPvKF+fLgmk5Lu9Y0
15oIyfQw7L+gXpW1qEU=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Cfhh7YIOGyVJiZpd5j8xa2ugbHZdDDpkNcw6vvVCCgnGCfzlen3wlGk0omzzJqyVapnfg0aPFCVf
eH/noQVGu1bQkowx0JKcNE5x1v5DKH//UNI+lq09SNF0WKlMcTAGlNSUzO8kgVv9uNbKUHDXodcD
5iGh6bHMhVPSu1QKpTfJlIMd2CMz0JfDQiVbfTaAGKvrQhaqVte7pYpnqiXM7povPwt/ntWHBH4s
XSF4J4eDVLMuQmQNy3vrqFdEUqmQFtLWgNRpG2fwo19Y2lRzT3ux5SiA0Iv55uR6x7AG21x8BZlD
JC102ufirdrREfWUzlClY8zmr+TUHpTF/SgPMw==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
UWceDgHVHZAg17Yudaw03bncVn75AJ6y0RYlYeqdZU3kMG9E1W6q5REaQAI7sMZSrC2g0zavsx4w
utskoq80P2avoebtdvBfjr/nBCQqUN3AvM3GSk85froboZgk4fCQ8UtEj2Qk7ob+ox/md7d9P9dw
2YULi+eG04dUc1g45wwF0ZoZdARk7Ml+fXMnm7zxmvqVieAEsVq6ETZN/P0pwvIpAakLTayKriGC
qcrb1S28bOuV+Na/FX9rxN6hM5aK7vSdFqja5GGs32r9UVRIkX6i7uqS9pWQDR0Qa31W3z6wrRrT
+2wzEwNMDKYuWVIM1FQo/Tp0NKa1Y+kyjahSGA==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
tLsJPLnIUk5FSxPTGLkNhAFldHrP7oFH8h39nfqyEmnC/AmGzR3fePfCEcee3I4TYySABpWhyXIf
m1jGiCuHfIpFkF2EJqjWmBev0bD33cbw1av2xtJRFa5gaQjxChO9URfjedFvCQWWwjlxejc9nD0N
O0V2XUDQxd573YmSBuByzshlxt3bujEd6Xeeb8N8NI8c2ZsfY4693LGdb3k6gtY9ZEoo4XuYVt6n
S2tNFVJTfQjyBEXbuCPqpwGf6bPdy2SKvTE/s4rSIVTO08J6bXDaEOBUGg13XVoJJqrayiJRVuQL
LhoiPzgOqS6ude1uUaMHE/SN9X/vt/6uOsOl2w==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jgk19ieS+ZYiySHKvgAHMus0OAx0HPJ59p64LMaYK8CyW0wSM8LIn++sFz9tsOBdLj2gb8IKpSVr
SOX9XXXM2pQFSME7x8q0m+EPg9m1+ghIpW4bU/w4zVq4NBjYydZCI0Hpy+X3op0a3+eENVEw5SoK
4R/zOL7aV/2nZ//wkaw=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
L/BPRr/PHH5da1O06dKRr5ST8eskM6lzR1UPuTvZQ6RCsFEjTD1HgyqjW7/ypnIq7V5TYDC553+Y
rJnEENzDc6RSpzenrYxw7NrURpUedIWlCc/PEf5Zq9gu1ESkpND7t98rc+uiAz7zsn/pHD/K50NR
q9l/gcWkOCgArmADo1Lw9usrfZ8ECIPKY2kLxeTYbh4fsrCpPQsQUk4NxX3N1Q0h3RRUCdHSFc0O
lvGip/vd24OK8zXDMaQv4fPmgToFQMUvLrJXErEUeRlkpxkcX6g6Zu4RMWwwmkNIfZHpc5K8Q3RL
MMc5rARUSXbNbpf28H3iyAMZ0y+EgI0CrKwooA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 967856)
`protect data_block
unvYCsvaDdPdbHKQym2cLOTVZD7oI7PVY7ko2LSc07Bd9gnnVqLv7OebVVnb2bOYZnRS9V6hPcbh
ksG/iNrBHeFWlJb+qQPTOydRsef7xeaC2S49dA3i1rJ8RivVHcDoWyZ1Au6hmPse/W45qkkH+Hx2
03bL7ciuBxSs3iXLm88FPDuQQJb/gOyfJ2KnIpdRiyUqBiOgBgNsvJdBRvgWXg4xVs6p/QolSmD1
18osMnhEgGb7amr4m5ZLCxhlPQ4C8r2u/hALHW7xatCG+Cf3VklkQ0T9AZbWKs5wWDUo8EnLUhEU
VpG/5c3uSdU2GZvKzEhrBHcNUSojsZCkiJyZZCbBCqA67HZPRmB4eqfkwqzDeYVQn1olAmlmY4R4
69ruGDiDA2Kz4M122xE04uVbmDkWeI/Lpw0JZQg5jZI5S0BqKUVi6NEDuqJ2lUEEBkli0LUnzRvP
LHttuMXf1+pewozQyTyKS8UOVajfCu4MMrg4fvuGPTaHQxvj8QNJAFsS7pTTl1feUwKSOqSz11a7
kM4mMC4hLcME0PEmzsLwQbf9IzaCNylRS40NosD7nsKBeD6D8PcWVZF1Z78e2UXY2j1jqjfyCxD3
C/mmDsRX8Zwfrekr5fDDPFdVIfv5rtzoXE79YHPoTjpv2326I/ahS1wFNISpKtNV36doa3VdtzbC
Q0M67OpEFvyQWEzM84s3BIDI5f+xSs8Ns0GghyIqhUQWLo5KIDY3A+Oao2ABZjQIpN4iYBx9wfPN
LP90vwhvwjsZMNZjuioPeGWyyTP8f1HTNGm0Ka9nIWxxhFdDumPSqCMjrj9Ni6SMuGwClXDcrziN
AImp3P2S0+raC3FLeTPcXKYRjP5wMelQWG7xwu/TOuqZ7kLld+UPfnfGrrIofggiQSVAU8MjRMoq
0HNGsl5Fk6J/9/8R2AvK65yHhPpaFAyUx1Roe7w0eCsJMyrflhLJDwctsxT940hD9lfiCuBGqcdE
/o9GtUyojJAOMb0v45wdxI/vp9S98TTZS+OqoQN286VYjKh1+C9ISPVEGEc0sn0Oh5zo8QUiF1E8
e5fuMqgemrGtReDNfEurs7NrR6slNulphwZNrdRfM2jkXKF7GPNebbU9hQtN+GgtGD7jdKSIGUKg
rTNXJ8XcAxLTTkNS70dvjdwFILi4G82qqfy7VTelpexwTtnTca9GViBF76eaKjCeMKduQ9oaivip
JRUmZonOSg1oPpngsPjeiTKqjTN3V0QHPdsBWzt1GwVpO9R/miQ7YToonayKrMBzJ7o1PrpR30FY
qb7z+spR76Hh9uLzGFvnOtP59SQMDkzX4M+/TnpmwPe34aOfEXh/AnAwxECkIt/kCEUWL5MSqinP
UhUBvC3Pr5VZtbSIVRNeV/59aZJY2/nwf1LOU8i4ZFBCY7aT/dEdCrtejPc6yucgA50bbpFEJYqk
GLF5St7gZ5dk8aPPjx6Qqm02QybDKYHnluTieh5IN2nH4A9IaGWOOpwIh/lDCMAJeaD6YdPopm90
bPwjwGTog8lT+AMBAcIAiuI1bun9t+OLAjelchmhTWKvapa6n3nsfwuAjLGhvtvK5iChxjo4up+n
6VrK/HfJxtLLQ7yjjVvZk+Cjz8ybC+n3ZLm0gKV4XirgydwvN+ynnH+Bu0RodlW44+BHCVdApHNH
U3XJl6Dux01t8guUdbFu7erUo3WZyy8XYMTn+16UiIi90V4JqUZW6Do+V+ChbAmzgQkRwlRLjBFB
ARsyVGUbuPuBXmgizaf+ZuLFpt3oEeKyTVAf8ci8/rTEufAr4VCWzGvZT0jSavVtBZW/oo75XM40
jy+T8ZZ2eF23U/1dhZgW+XQZppvsfQyV5KKdsZI2JyEX4VxWTD0JQXmJIPRI5n08JZe2k9NpRf4t
jjKG4Cl88xXq/tiTawh6eYH/Hzk3SMkQfiNj/ngdfujhFThOJ3cVIZ6Ldboh2T1XX1pIcmj6VY2B
Krg3g3ZjWTMXA344QoxX0tfoOubblOSslnhakZRzUQBmWJWTmp02V4yZFhIp1P4jw/uvWIy0mPcW
Du/IUL8CC312Y1kIQWdmITH8NNAX5cF5dXmwvOPYf9aBiOcYQjFtdOnXPgrwmpTpLA1FI9Bxfth9
MgfHWGQFjsiauQEggTaONA61wwkbiJdEanEQCdDWnBDVyLjgK+m0vwE3GrXtS11zu/lBxhRH49yk
a5leWfgPeJFiSne2yupHYnXLnYWC+leXRZefctzJkQHtyCjSDOvu4tD8mdi5klsNR5r8A2o8Jvpv
x2g6R46U6s5su3hRCESrKvVbeanw3Du7D0Gd9byhatCBfbMzDarPRoUL1h8HUff43FCjUGRDDYWK
1l7PSIi4Dol9DCORSG2YeCXu7DoSbafQclIL7/eHfwinuMb6ZPm9RzQQgTIEDsNMUItoDKG10Ro1
85X1LDDORVQPmoVWQwh4J6mKsTlPZWSDEOzAN2Ml77A0q0M/FnqhQhr0nT3R0wGQfIinIaRoF1h6
Nf2mgqyvYevLJd3mLulUaZY7FLuOy6ILtYDaEilzj8hog88L6DY3JuCcKgLoiUbf/wNbLR3DJ08A
DFvmzTcUvCzMm/RZzSZQw9uBwU8468vvXT9Nf3qvrO8vJir3CJfkKotF24gieMMuhEEyb1VehM5H
LZ4kcmZZjj7nGco84ZkTP6LEfAMQyLmg70d4Y4NcVyrOow5cakWND+DYWizjKrkVim+BbeCqvFNG
WAEh7igLUhAeKhbz+EjsfSqwlBQHHCBXNNUpn2Xw+rHtWeszOwOOyyo3rIWp/9OnJF2de6HB+44q
pt0SNqenxWapKMuwVWMDH2hnq91slaRK78HZmkLEdwmlA4AOWkRo6etmtxzryBxOjFSNMA8ACPro
6ZJ40nWsG7TQf8eGxgGDSKhnWIW15eBFlU37U6rOTQJhhcfcgoC8XAoB7c4oXl6yYtbs40//gry9
QHgYX/pv936UENHSOSEx/WkklbCOR3mUynpzXX6P52P3WfPjAh4YI2oZ1cAHJJ1StaNBc3Pslj0D
8aJD6RfDT3OmHLT12EyXd47wAaDce8PFLkjBtjPIb714GPu7ymuExfhJY88+6VV/nFpa42B5pisR
e95naGZB000xxobGpHavfVelOQKv65FEF8vP6OyWdrnuECymI2fkuek89PC+EicqqAap0ecVp9uV
1L2/o8PhQK6IW8FdlOUCRoC45+GzcGmm4PtWcZdXFzqRUlGLQGZwhzkF4Jl/v0MZrwpwHPvLxhgX
91Ucz8jmqKd6Qi/hjOOpmbGPqhjBczFU5y2gfXrRrGvPcl/7T/+2v8WAa+aGBdodmrTvg233xavM
kY9J6QMV6ybQHq5sSA4D9GOP1leYj66IZiLW9CUuLlbu4C9y8mMGcSQAG8pXupAueXQVpDccHf/l
R9D18XbjMQD9QU79KcSvIJXnnVv9zAwm4VdokjbTvQQPy44IfjftXFKasXm+lT+TY+kiGH0QZ02g
lbWxV6NT9/iY4UNMSc5os9W6uiED1aIvzaz1G8jBWb0IkTV39tAf6cYXeMWBFpp0VXqe7qJp2zZr
vZhaYRRH/yqTvSae7IIJFPjFGgg+HXdwCkZiJaUU1rno/7JVmQSYJBbwNgqenQu6MVEf8vsVZXqa
WXOfRfTXV8McHuPFEmom34suPmwEDj4AK6lIETilHC//9yBI3SRXA8LWZpAMzxs12t9sukgUJZ3e
Yl3vjbwwUZ2KHkS13fxGoFAOZk8BG6sSXXoaTlzRQ2bsFqD2HKf6WtXMRR+8KtyZW56UKUAXtB3+
clWVlzU5bJgRGp0HULUH6ab3xCtgDXH5U2FgNYY6ImQwDktVzcI9bQqTHHFnEY5NsXPKpzJLZ2Nk
6LvgAfR9vTkyOmcf1u1fSw3f5aVyaZT3edZh/OZQon4g2349J6yAcMm+YBZ25h+4IGYwgQehrC2K
T1dv/cAtcD6H1ID1H6cyYuYmJgr0IEo16YpkB6k/r9xO0wHSt+BLDOcnMPaOSaVztIeDOmnMHvRy
U788AgzvwrWsDffJ3rbHkkUcPNcRPnl9/0+9HsOlyWEC8dn5a2qLUs2bcfgKD9Hj/7y6eI2W+YDT
C3hsDlPeg1q9aBKC1OUNyFdOVURm62mHCxkBAiahoLgNFq+B0k4UIwr39KOdm8qrzkf8JhbEEnh4
4YJCiwFIhfDbPHUC+bYKuLeZgOj/2KWZkrH1Idy6CjKp0WWbQyi/DMAozAI5z+RUDGwaFa6QqK7b
WbfshyYuo1lXqOXQJvIp/+qNN9ibRD3Cbhq/1E7xjfJ9V86I1d3OsxRmhh70l+FTOCVNdGrpH8d3
4zOR9TUfV5SpHhRg0VnAxUVtYxsk/x1sYUnCwPMfABkkV/6K/wQN316bcel7u9yQ4XCoS6EL5tk2
I/XRYdyL467b1ZI9S+fT8jlXLu1RLaWFx1vPoi0O8DSIPNZUe3Zd+6KXjUl958WwmWrlj2AWZ9Vn
02SKWuGkvyPRf9nPjyltUksiHyZ1iGLiJIF4QCNP26qlVNCORwAxZI2BPKsLPK+x0Mz67i96hyIo
IZ/Rb2ABHCcmA/Qq+JCs/AT/hq7HHux6zqPmzsVqkkvVIXGqyr5zksrU5idA8Xd5+J2UNRpuTLsM
fY0j1ygTRlPwbM1fY28sapBBUAT6Cohbd1ZUTy0ZGyk+NcZQGp/lHff1WZ5NA3UhH4h8wofYwYZO
CVUyHRjKH1sYgeBp7Cbz+Y0WcmHTDIA0JCB7kUWTLwyGTh+JRjh0pp5zCfcdqICAqMkfXL7tGqbZ
2YQ6EnV/RXxJYZ0KV/hsLgK65DoAf1uF4G0Acna2LaBbdxfVm1dKUda6K6VPm7R1wpMlOTm8rSRb
xx/zRZ2b1CZwAsPTzfBJHujqysndDcs0bXATpMvRpO6oQyPs53GP1ocTNkfwIHaTAc5aMKIDcfa7
g04HxlJ2yK/VsZ5SYXv3ROkNoyADSf3JZgJP1hfQAWo8LckJGgdkjIsFEp/Msf9De2dlJ4YvpwmK
ltCP9Dz2q5WDxPWA7Aft+XRZaUMlo+8eb9c5jAI4ZcBGZwM94Kwj/3qx9XygcsEV47m9LvgbNWDC
0Jmj1fJbV7y4P2Q0qZjQQgzDPjRJEGVjEUDAJl0N5Ob2edyrS2OjS/8S6OHpih0udi/B9Ii0hI7c
0ae7AsJvpuKAoCZJGGPeH0QNGkt/G0op+zO+KbULWc+X+RInf2G95alpAAdzrAGK03BAO+DVfW59
iJhBrDraFeJUyQ9RcKrfot0i2sy9U7W5fIsg0WqPvS+NAaCbgRpOI+/EM8R+kOtaa4kjVakKeirj
F3iY5NXqLlWuwi2IbtH7OZmd2UpeQdyPEK7CK+Nm9tBYUuvXKZJ32a6ZaylwE6Zh2J4WrLegKZzN
WkpimETiMxJ70e9zN2A/C6OiTO7pi1sWsBx5ME28L4pRhVYmE1BA9J+UvJr7em8EIyRV2Z3uSdGT
gkvEzZkKrkz77UJaQR1g5dsgdCG9wxNqSjV07AtZoXnduOQ3MxqCIufK4DQCzVgaS/6s9JktlTbx
nIU4fs3SYiuXxKJF+Yv7Ke0fvU/E9bHhjbyLPDNLljQl4wAUxCAIUqdptiW4qk0KErACtVtjoCSq
g1sJQsJWMQ1lZ7Dp+T1fPq0mw9VGqVbeit00g6Kn9b0STGe7UiWD3/4kQlwvKomYx+BGvORa9lup
+sA4iaFcSkN4gldd2/imhX84UOgG+DwIQhTOFawJqeUt7BGGQpuEg0SsLLpioCil5vcw5+K2OYUd
19ZY1xo4qGp4vNLjWmvyBHA/NT7BCOK8P87sOv7FPiPSEMN283LH3R3Llaj089le6g7yXgoH6s+2
OaGS773kQI4coHsFi8+b189pIZEtze/UWyyCPOPNjaAqVSUimmi9briOZBhaAD7MpFiGppCRTJOq
34HG3P72MMcUottXJUakBTQym7Q2A7et17fIlWEj92q3JosrgWyiLVlwS6feNygBqsdF7dy7ZesD
PPYRnJSvV3qO9J0S3mex4TKUe7piqfeflnGSRJ3JJqn6c29z/JNYDsSssaE/yfWy1O5vdgkM6xE2
6D+rOBmHPAZ+1Xm+d7Y1IBUvGYUhkfRXKHahZJ/j9e5owOxxqsSvj2L2PqX8SojiJnZjQVdWqi5B
757qb4ZTWBdQ+lgNJT1pqPwkfKWBYctTqQnua19tSBelJ7mKw14jLK5wgSiJzwkSm6MHMd2hdfsK
umHMCrFQ1KZh60CcC0pFUSG+aB6JABSdvCi018DeM0UjwqgXpM7QQYSyy2TWQ0g0eBzhpOfwZRBi
uIUxp08nIgV9Xd5JR5MeiJyKLcVcRJiAllqPERjr8Rlw53zrSMb01LHSv5yFlmi0wtQlJInqETI2
iEu0SibXW+YUvYoumZG+3zBkQPM8RZV4SMe8x0OLEi9v0FFHxq0wM5VvAIPmQVzy0DHaG7fQjhkn
GTpCrWhh8X1raw40mJq9nb5oxnxp7iV7C/inpvMXMhzfHM2RJEg9qd2hx6shTJBBXqW4OtyTpou/
zBI0cKsrXjs2w7Nm+wAqSlAwHvyRqzPTiJM0mQb5+GV+pRFGhenzUD8efgmK5E8VsjVN1aDfBdDT
Y4aVfwjZOjNmC46hFC1ewscjmz13GLBEGyduXd/cVOnbjwJg7oHm+xcYZM/fj/+YTEy45VPJUL9r
pYVOzcciJSvOWowp8tJNSbtdSqwIMrTyKCGVHTEPMr77zWf1CLuOMHKvPdfe0rHBLIVeP8tEJO7O
7caBmeyRgNvq94zz3Am9prtxWZp+gDw/9Rm2lY+r5vju/+DEObCYzS1KfLIn62Qcj4AGyZK6auLr
iPZHgfoguNtXnXO7MAkRy7fWT2o0f5e1npyOUyc0YeUH/+OJ9QqVEFVRrkbrXVFMSQn2VTUnLpaS
kQ4PLjRNiGNlZ4PWpD8qPE+zF+nEMvqrlc1DmU0tZG8UVtdiL+zLDgu4H2lnr35LSNX5a23frAkA
t4wojP/LYz7M6mHwcBnAA7V7zWDuPS8UUv6MP8+yFZQuWSPLXaKQUo+uYJS5G4/1c91TVVlg4Scm
H2bt6nrl//qA3S0ptqkd3zKjqYQvQRp4kq+39IzoYBghL8E6Snv20zKc6vJD7lkvL/zgTJz8n36o
6e0w93cfCLfUmXUw04HmJQ3Pdq0+12pOk0iHwERRZRAdcgzFio1XEOtx22PbR2g6wVFF/oXW3KLH
Nd9+37fxwiKAi882jcA2bTpm4MToK3ZpSvNKV8uhw4LqHHrW7aD2BIQBNXDzxwBHFqp6HRc9Pbi3
VEGZO7iKmTm4drUsa3lp2hsvJZtD/goScYZ6u2WA48bmm94tNGhYpPVEjggWg2srqbcTflCLysFj
gIQ60z57TLYr+u7kv4fktGoehOJ2CzGm3SEOOvcUJwBzV0LIQG6+md4ZzVOHSN5pgQyMq2xllmzc
baCYAQM3BkkoCekHmfGcli9sfWsvPilldF4Kv2r4xtdgXPl8+XDs7Nh6/W8ePuqQLoSC4ruMh9bZ
XQgzngiEZJkgzBNQazalKloF+kXDdYW4g57KVveutMAQIhGR8wTnbmrhHUaqEN8WncmT0QonlsOB
xn0R/xZEMz7TczIfX3/og6lZzOL6EAl2UGGSDgXyjK4y6XojUydxP/1oKc0qd+6AA6vCFU+FSnRQ
ATKqgoBwfgtE9Ya4E9NLWMUiaWe63Czv2JmurtvJRI3I3uLdUOY3b01xjHveCeIBf/OSbnGoK6bk
O2RLePW8Kp7TXOTD8Xgq2BzWYPhDfRkeMdb98rYpuKg31pZyHPf/+S4tWRZGpBMeG3Ddnchz5vwg
tGNELh2XxipD1nCHpkzuZZ6MCCyt88PXda/y64sihwU8VWHG7IzZAZ9BzGncWwfqPYtOJmykFWy1
KdieAYlHx2JbA02uQ/PtwRu7gNmAH8qpPHafx8198h1SykE02sQHyWCS2ynT789gRdbBKc1/bmrE
xp2a1Au0NIiuvxk2g59tyVNgY/C2ZgH73gtKteMyozdgT+PDGBhNjvLh9AnJltmO2Cq+XSLAnNVe
4VuC2zQzyWsicmViD/HtgCgj2cQFkyhAbDNvHUergkF0u/qfFQyKop86bzAoh1CBmvOK5T+tCEkg
CTMbN6ZPxB9oZEIJEqlD5qlY6ry+RjkMW9ZCSUmgD0aIMG0l8+Oe1wSX4wY4cuEfHhpj1kNllChf
SHATMOrAeQw78JUjIChsCtHOY3ir9mtRS9tdKNk4COCdYjccayF0+SpI6EbgERwmev9qB/owxq79
AqXZ0K7IMx6rk4et47xgrqyZv3O2dDst/h542qbJu73zitDMynEKHCKF9+BdBYNkkRFqPwNFrkHM
+k6ZWFKjz/4BZsf8dnxykSYy8l3u5Na3I6bSc0c7k0vLRSSfPK0NoXxbdp8I90Qd8qIw3GXP++F0
RoYIqggYr5oZVkaYKN8lngATXe2DHmOQ7tb/pKTCW2f2ZHTaURlhv/lwfHgS7aSVPYq+rwImBGZH
5BrO9o0BfQJ+FXHIPGt3W5CmceuWrgVNILg/Wtwu8gXv5SjvK4SGcXlzqD+i93r7SPYEI7O10PAq
i9vKCC3p9W3nr+mHAwJhIfDmobuLjEnLygz81YlTFAsbz7lRCQHaO6NTuY9zE5wbUZBVr0/fo/Q4
Mr39Qy6V4hyoQCj2XFdqw+O8yQ16YNClh1KkL3W6zU9KYc2athw3879z+dOMMqsF/1Pf3mIWFzSi
j0DibwAsyfUrm1DvHuEyGp30vF0wAgHpJtS1Rnwoj2OQpx+LT/s1NNEMFLX2D3ov32PjfFWG6C3q
1abinMFFzJqFwS0olZdYJYZTnm8bhYSTDHSLXHlauhSUP3pBPWdOJw60wXJaa9LoePUyDuL5HY1S
uFe88jBXmD0UUtLQzCL2rFoDJSlWqDlCOdmzXH60Fe4ep02+V4Rpb0NBJzRVr2jDU/dJkQpYF0TZ
ew2Lhp0usRpI2XM1z0Grx0p1XRNkOt46VaSOAj4g6k3NjfHkygO3juDQpFnexz++YiSM3CT5Lhcr
rKpB2bADxXbmYSsUEBi9NIeUEtDTOQ7YLktR0S9y9lOsOlax/sWTDZdf4C0filytiPO5wA9zdltX
syd7FyY0c/iENVIhz4BxQhItZQTPV4Z0+8aqb3fmZ+XZZKVkw66YkSVWXmCNWKjC3SprTvlknh/I
GDvkM2wLEhw+kOKEhlXNbaqCOO8JQa6frVVpzBPzsSUBX3yej4S3pYzUnPI+8TTdByG5/ZwEIy0z
vNY42r9EoPgakC6CvUx/weOfrh/vAz5qBkOcSge7nONRs3s1cSjoN5nGk1z3q0+xwA6W3PRynbQ6
Z9AKdkSvxaQT+3tWnHGj1Y/YjYosaUMKnT5KPWhgJkeMku5RXYrULJWe0ATzRjD5RyY/amBIVtxf
yWPsF7ZRslCYyVAxxQWtG/8p9gLvrJQ1wJFPYSEMHrDKVvBtu8N5U3UufF6X0dl/AXxA2mqoStnk
3M5JQ98GBxd79GHPx8yVZX/d60lzbg5siivr3U6Hkbk8ioJQ5aKZrg7G9HKefFFv1dKfuf3UcTam
oMhAFqCpeRVPWef3C3pEy3FdYWaUyuoWAvGJUZ6zf34qUtjLFaqJgq+RTjxjKhxnVvYS5rO6Y4l2
A8iLtkPy3+HxY0ithqDD6fs69/enQVgpn8LZwnNJ5cwda49urZKefxSLMvpZOOM3TQdLQaf8dpaX
yh4rBGIp6/oUEqUpQxeCpglaJ6v6JDBqsmcNTb0yhpYBlfkqA962XVpYGCbMI4ba73SubTy6qO8+
WXPN3IgAVVd0etec8ityMj7DP9wA6S1neU+A2MUFTgJanYDwJ4S0wtlDMtiFIla1VT5uPkJAss16
H0QzTZdxGXOvdXKx4rLeaLtB9WtAc8v3fBZ4xminagL7wXDP3NyfYO0QSl9KqVWw9az81YxZ1ipw
9aB7X/VQWk1/5+8008J6Ks8R9bPqoFR6p2WJSyO7qu1xowIJZEmibIKEKQ/tmMnZ1o0lY9UQtFIJ
LiUxJRU/QCLkXBJfkPPtAXk5+M1q0Bj3ewp9e/edLgnWFIHZStgbBazj5IodtoLSNoxmIkJmIaGH
FO7eGwIWK+4LtYeI2MF4ugp1WquP9NjbJbL8gPnDh5hYroATXCaLQpVL3trS5D8AE1fcngdn5uyI
sJNZtkGg8cKRTlN6TS7jsxw4uVgbEi78/P++/AdOlWakXZ+StW0jY6aJnIRWhLevlHP//xdXBKIK
ewCRXngB2YL4tzcUnDkPetS5CALCBnDK7FNbjyP/7+pTGMsTI/DrMZnvFHmPJnyoSUJax6kdptep
/wgEQPq3HBFy+2RTRG70aZuwgNEJVAlZRBVRgi5m4MtEVE6Ja6jVulskq0oFe5EkbAN3CwnKkdAy
eg3XlD8S1xkR1FnG0/rthXVv9yVP4C78/GaCsGCXHLkt3NymG2p1lwKJtP1PC5EdT9TjL5zPritB
UYrEGNvw4h8kJDMz8xx3QCdjO+XpVHwfoXGRdb5kaPqGDFCDg+wPUmFDhen6OQq/FmPSfV33HFU4
xLIfH7pplKLpwxMbGVRtvPgfHAwOcOT2JYAe1XgT4pVQ5GsnXmLwa75VQH0O8PllLf8z2gzoamMA
liu4GUkAdXdVZ6XArOKUT3/DbdfHfem8vEyU1LZZDqjxdpH7hYkwUBK0aRJTcuwPEzDHtePtphXj
B7YVPCrHOqZrgW7JeLiulLMYFA8iHctNbCmaEoNPDKWgO2ApI/KBjCgtzvHu6T5hpkQdTx5gBwgT
on8b7KZTaAHoXKfU0uiBGM7XpPaRcsLJjoYDwCM/veuSaioQpFRYykw9f8SnBik3qKx2RW4EJgoG
yuD97THOQ3esxjnmWvuZI+558+Oizy+pjHDTkVLWpQvYsXp6eAllTWdAqJE7WxP0LmeBfHYIu79M
vmLQEoZBbfIcluwT0e3DdWl8BsTnlDVJfN5SQ5kt1Sz3CDXkh3qkqKSsBIvX/0FUMndpDBMQ/Nlh
xZZ7IdOxUfbfyoBBzYNncFUEmVzU9MwiUvuG1lCKAAOG6gHS9k0W4EgAzuprC+NszjeuuIsbNOik
rt1OcEzNCwkcleIniPuwUZmn2HQGbzjPhyMtc8YwhiIxSU8RBlpFRQgRvo267ZrkjtLKBg+7X1cX
ZKqIevJONAWyYVkkfPFxVKMQzqLDhGpCrJHQgcEagSnJHYc7L0boFKdqi4hFSOdqLmslbguSl/+H
WEKv93pag48iZz8GfEzelKg+AYEPkBxV7plbw1hy5YaxLfkFP126Ps09zDriJAd1G9KG3dt1VTKS
ORDunr3DL7dkgQphsdNjQAZT700Y2ye0DC9madkYpGOG4F8n7zo+7ZxOg9wUDKfzc1NKiC0/0M8I
5/ow6jQk1LLNWjUE2qyTlEQVfdh4YDYlWMo7/phmqCi7POecH1/VPv8YR7GT9e5d8r+1Wm6XPPzN
xYAiNfBhvkwveSPHf2WxJ5p9MMhV5WDf6vg26nO0OV5YsWg2xDwE2j1cxSVrVLyWto5Zg9XnxG1l
wxhgM+qXWyalFAPB0YrWw1TLdKcSWlCyVZBLKk2EsY/cChkkOHvOarq74Ik6bsW0Kd02yGi4Rqv8
AZWuhKqa/bVbICQiSZ3BZbxjTOjV22IveqtgGlX7YSlV6HJB38z5sgGoyI4MmfGe8RpiJuQ97pwQ
DAeX9KQC/oymZj01cATAaxUI+Y6tiorcxh3Wh4BwKpa8NAQDaAuyPeSeSAQd3dEssVtRzD6Vu53t
uiDsfiwlrKm0oCweMceFEBlneDnUrUF/XvI+4g5P+AZnXC307MRHxqJ/cw9W9/86XiLbQXnhRHhT
zOSJxDaHuafdOdsyo5fEdLUMXZh/xNl7zIWsc0Y8iWPXx84D3fxWmQlgz569nH92E9eEc+osNI0s
omX3qEks8eJ7g/bGGMWgD4fncTTwGKpcXN5RTNKN4pHbeiXsVBnx9ToHdAhjotnZy+0kOIpPFhvK
D0j3tVjgbMUkB8ekXpApGrS4PajecIJeE/0k/BqpBQIEuHirdRh85XX6iHIemoYLheWcDhgsI6ka
CJrYOz1Ez438XJTD2WCX5wxUmzpx4Y/YxmLMJbwLRj82sFHj3BJJvUFP7xfrdJ/1MQM4g0Atm9ji
eYLYQGXy53M1Vw8DGXtiRpaqZJ2ZZC0VsXLVqxLi9irmSnCIyCA8R1ISPR75C7nC40H2Z/h1xmIO
wTT29GQU3fJkRcJzeHDd4rSz8E2N1kNe0ALaqLl8q9FU7rI6X/5vOr3diNv15pcuh905R92ndwvM
P2ycM5b4HfdH2Qsi8YgxATzTHa9mKBlTizpisVrHGnfa6z638lhCKZhWG487CTAOx6+WJaV3gvLT
7O9TaCWxV3cfFJ4VVKhu2zhmD6G99a18inGFrwEWnXnQa32BIPPMOq7kmbREhKrHuJnb4cBBfEYi
tEutbBKcQaMcTCvt404Chg9Pk5+yhFFEr2Hd/YJk4hqus0E5AnWEofwDC9svQdrJ1StgTBP+d3HS
eqMXFbMaFGuhwQFounalx54Lv3zGjvnx5yVm69M06IMwtKNEqnwpA6ELqhZ27CgwWQ0s1PfpoqM8
ozg6TeMF/L9Qf+iPu4uVuovaO6nv8SUEAoVyMxffLvUExfHgkoOQmYqhrD3jzrOxnevZas1FYgtT
KMmppag3XyZrdm4hpT5Laa+47qzQ9M/HRp7irpQYit5DN5fYpETKnUYP2Xbx9D1vEcO3dODbs48k
XV9SRp+Ztfs/1W5jRFjGfZdcNUjqOLP0BjKZOojNgYuR37nzTczuUe9s+B5wg2bfZbGXAzTRixAS
scwyFMX0HgO7O1ik2gv5FCMoMEtMay8Mf61cY96IsII6fL4Kcq4gFi049gpRjgIzG+ydp9QsIm+v
Q00WAWzOAUJw1Sdw3LqqOAVzBDPX8z/QFolQl6VrZcXIqWrdMcmvKuvk4AASHprj92WqAZWtbpJB
jou4Y5eBI17W1y/zlRclFIgAAqTlmzWq3TqjbSueFfGqOXgCNrB1CXtF6rekDlmDyrlbKM99Y2GM
fSh77XrnTrn6Fx8v38OgblLMg2MaeTa0PtWcre+52NhnPhBaUCOcLT8/rHIoVvvJ0yHto+Vb67ul
jVV4u5aStANaIgW0PCMFpn1LyA1nBH19gf7eUEkeeFgAwB+q8YJKIY8WZ12OrhiHHkjH/p8fTd1P
PMQ7W+iGoB2nmimG2WmiMYMIE7GPv1ljmTO4kMXr+vQcIS8YP4oDipGccVFXeaJCg61mdCIGFzVq
S6rZBvTx9Z9uWLHyaezgPAvGqSKxUXKfVva55WUP6gDiGcKR5AEcwcf2x1XS3pYnUwyWONAlIfKA
XXj5ihTdDlY7kHGLgPMcKpvvXQNs1AqPoiHuwVUy57Ixko4gxPrhaW5519aEj9wDreyt8ppvNQb7
EpKBEqSz8DAprhDrbgqbTkR6QQHurquGyaVDN3y6CSskXTFMLt+1ZpnFoTS2n5JlwbAQhTFa9/L4
IYa+UWg2d9pxUqMp3FwR7RRIVR3HNPr0ZnQQ8V+DD8mC+NHlQg2ouA8rTm3ekkqU4DTFfq3c1Ez3
8IX3VihJa508r5pn0MpKf6Cx90V99AGQ3XqgyxwATwCXHc6E1KYbFFPyXrA0Vzp0haxFCMP12Zv5
Z4yC24DLxAfMkn5oBU2sDO2punbPAfz2pVqTxDHmiNloCvxXn2l2W8825L3ZXhENhhVnAkz1HtgZ
6Scb0W7BOi/QTgysTzYUx2z7YUulXyQU9S6eHTVjEV3VbkQmwrE8+mIpcg4myuLnq2lpqWRXMqMM
YsdU2Py/TWbJt5osne/OXcwUzIRKO5oC/KRXYX6kNoQKuJK5+ID1CuZ6+ehnF7SyXF9C/yl8vPpp
9hd0QFE+ZU6E8RZU7/28wNqGo1Lx3l12ovXXRoEF5BfTvmWBPk1HwLEmYOv5p/c+5R7wp8KkpTZ2
v7aviq/D4VFJG6eXc20CKnjmMMPvkUFEOfh9U+aLEzPlSkxUpPX2FybFIkGMaRRCtq+u5H4Dsrc4
7GkcOkfxehBnNCtGR0FGSr8j1KV6iYoQZDUxnWvFtp0LSbUluXnE0KYKIlUvzIsmGM8ot2IAhxeG
cPGtWAQCwtIqvT8qsSeogyLjPb8G2VP7dXMXo2yKTfH4SL0Id9SMc027SPa2XektH2pxkWyoBa8e
J9r/FH4ZdQhuJCN7A4yV0loLnTX4k723VE3BDhJRmTE4C8LJMi/sFcWc99SJ+jrgSSvptYorFh53
gMB+ufl3s4XOjoR6WDI4hyjOASmUWtDCupkmAc4TH6rjZWvlzGEtMdkx3in9MNtq3DE7aVybyqa+
h+bn2lYQbkxCvLshgJSVb9eiUjN3lIOFtiqXaxIHormKy3G2Z9XZAy9HJ0AAXhIq/gN6ddm39VF9
FNel1jjfwJcA8YNV9Hg0rlZWvvo49iE4pNwmmGR1S38ZXIDOa0o8vz/8ITNZAa21UHEDxu3C4vou
dQDXrGmNsfoMzjyX+gdOAnpoSBH/P+VxNe4CBon9eeXiVLJb4Zr5eKiud0koOtrpIvYEyoPhZ9Wu
IntjGNrv1qNrGxU3dMzkd5RomjKzJOhnqUZYXwVR2bnMS2fUHWtVh1YjsmaoQkw84qBAMUH18Q71
EEleMuiiTmZJOw/+sWaQXjMPY4yhOw+A3ufEzl2wBcmkHJYXkQm9Mxesqw/GebtknSX3vTYy9l7O
2shAaIPxz8WGGAoAv4l2GBDsurSd176IckaIfAVHBzc3jVnQ9Zt8BeNiyndl0Ee2AD96m0KImhW9
taNw/pD70nQuRkXJRnVdvI4r2F7u4kgV0mqQfJZwKNw4H/Y7D03IZVL1z5TCdVjTOrLk5sN9of4Q
MzH1HLOvJ54jLVN4eFEZLkS7kaffvQ4+u09PQNeB50ZM+Mspp5j3lOzno2iomn9APQ0mMeKMMY3r
deLnMo0me1lkgPI4N/DWZVOLZdmtKqkmjvJmND6za14e4Nhi+++veEndYjQCIVIE0e0gSBnoUiF4
x/zxp3yq3gx1ldeWUMvbkB5WFCZ00EyK6gOazJNM5xEwiNxJ4BrArHHqLK7l0cKnmgPC7niA/F6+
+O71F8Xu1qHjbZObzHSoMNjBDJqFJqnnVHHnwbEL99H5X9v0N0izwWbjldc2mYxJ+STcEwmDPALU
WdDj9ccMz4pupdoH1JW/3KzHULgYOsSzWBYuyNAK5vBu5CXgP8DX5hUVzq2vUXUaEoqYXXsIr0fH
Q+EFmOankGwcmJDJPdBBZNOpy8ZI1qMld3nuDNrcNz3Or5Taa8e3MYSbeU0QqXzuuM6vCrvAKHqW
Ht5KNV/v5nUZvXjwXgJ9JXqBmKLoyhH078KNISUQEmY1jUuRiQPqBxBudzahjem8rfdkLC2gQfPd
9QDq0pHx5wXFVJdZPIAjLRc23qqlieA8B14Flv5RzFIQpoQ76/vEjMX9s49V4Lyg9fFYqXHj2EYP
aWgBj1VbOAH3RdDVQ1DRNSoPG+/afeotCKOTNUQvFy9k9RPUxAcqeOcmobY1e948bXiv7cdYMiQQ
rrZbcnKa8kkWnRmzGGDeJR+bCaLcv57SxvIqjiDebUIKPkKmmVKQzbmdKrTyNAV3ppIdfmugtiFn
99scQUF0NeM02aoTmNiwP1V+wviX4U1brJE07l9UeEDdDNqbAbr6lJcdERVNx6XW6S532mFOkfBL
6I9RNjVIYL9Ym/gJ+KefIN9dZmpgPQWwqYSh8kX0zRvMij/+2RL7TJFI4qoXssXGkyyH180JkEL9
nOO41E1h7R+XE3u+m8U0jyxO2YaeQ/TP5qE1aBtLtUZ3BvH/57tdfnhbPZFZG8EdAv1s805gq+T1
+8fQXTppGb8uRSO6RkTV05geX/yvksPyGXzIbWgaqdPDHI2viykGSDaCy2LNDv+YqmEMX9UWB1UX
buiaM4wJ+r/9B5J0yG5JC4BfiE2GNbMOrP7LTPXw7HJUZzP+kQsZPC3z4wY5UDIwo3dY1/fWUHo6
cx+pkd2dpRJBpmBC29BB24xfCy3+2ldpDkW0weH+H1StJ3EOUxV6ThnN2gSXWtmceQOiVA90x5DM
pBmrCHEs7NpXEoLOOCL/JkRmRtppz32IMkqI80ZZo07UV6MuDc45GiSGvS227dUmm+0/M5DQBE7o
Au2TIAcn+wAvNh2iC2uNan//5pTxqLfFiHj7jZkdmUAQK7cVMf9a2e3WzTRd68t7J/+0lEWItBUa
SwgxyyNDegXgdWj0XzMirtkYXLcdLv0+ptKYM3Lcvs/Y5uCBykmiqAb4ZsxZryQO8O1WKQPtwrJC
OvmJJhVAU/BtXMYpRTRLepXGwfP8RSvD9Gu0eHH5QEDKgkdjD6M0GtlH8W5cb8UM6+V4HD50LK/A
ST+KBtCYXIdyl/tSKqkhcCBuqOxKhzaJKBxLNjKRkPReVcBDX8TvmhzhZhYlQoCxxvsTowOMgxqR
WYGfrU03EfW6G6aVPS+CCEAlgTHzclmYjbXe5FdMXi7oM+m0SPu31uqNsJVCjBw2HSndRuVC3Jnw
8pLV4rQeQzNbGfFWXkr5F9tcT85EKhbJc5K1wT+ZKGiuFGA0OMDUBr4HniRyB7Eg/OnDkgxnw7r8
9+3qEKlKrM4/Sek+zGKO2qR+qG2DLNKW1OJZe4hvXE0xzPHMwjYOLKBUsznH5+kDRtKhTlLIjpWb
UALvWRv+aMzBxBIoLBIywPepx12sPsCPkpv/tu3iSb6eDJfqtl7G3QUPVviRsh1SBkcTTWyYU8Gh
S/JzD7vt+MJtinVbWw2dNapVW2EF5hHzVWTaBW9+o+RNRww2ZkCspuJLPlQMih63KHSXdkB/JY+L
ij8Z95VDDcayTcfvJVixE7yNXUnJwtc8Q681Fo/64ZoPveXZ8y1/Xg2SQVp5GLKpbK6bLCaRGQ0+
ygSLiCwmO3D1ca3F47BqExAU4+7ATyvrgcc0ASqHEDbV5g6QIbWnjq6yQyMTmGeQaq86uZbzwiKR
L78S9iOjpn6gQ7yNbLkbRT0RI7TD5OQY3U95nYCkZhBbc5t+/VItqWIl6OokQP41KJ/hehyKi9m/
IZHHR9MvJUADq/v730u68xnKkRuM1fQ2iIReovcoRiEnaKsGzvSS4GR3BscRjH5z0aXhjuPm7Hv4
KOXjB5braitQpR0nfi9B0g+QyrvDzs86AQIgCRpZvYK1qc/9GqCR74l2zHsDfnTzNOzfVyNdBxAZ
JK0LDrs2cpe18R5ImPTd9FEFRB0NOmUn4pcsp41Qe5Lt5NFn8hsKWsr8TbDM1+w8/DC1AI/ClpZf
KO9uBpmARyQl3OnBM2jjkVcKvmOY7ahtHshtVw/NWa/3KPUnlUe/hqVaJb3hXwGvji62AITKXvBx
5wilpt0X0dziua3X3u3t6ayRIxo6WeUR3UUc6Jbk66KWwiVzuwKR8opx7n1kYQMFKk6C3O1MNAkh
xzRpxwQzgDAXEG6o+Bq17PvdUD/U6qcAqlVZyjLyP3BzNBYGg1jeFwnonm/Y0Zwybe5jEzjCrGMd
yPkrSoluyNoZ3oQ/hK4R8YHcXSmCyYxP1cre2p4zD5srT/6hvDLf2ux7zwl3/1+rrPRcavjQpaWc
vtKCvas6AltzG2DtJR6w3dP0bOHzH5+4W6GWM5VvFNJfCysz66sUq+LB+gngTsTkMhFdC8x8RgRU
5t0nWGGbFxAYmJVCdt8jMMPZRvFV1EyjGmnHdubbivnVrexr06LOqQO9cfPGEu5B01XWLGqRSbwO
DXMLvvXbs8VEd8/ZXnNA0NRi6MYYomyOTB5IOxI6Ig2FXDixxQRy9GptFRm7T+0HTw0byGJhYzo3
/9AZiUXLOMaWp4w1XBUo4Y6y7IPgYklZZcp0oz7CeC/Y+dvy+5GLVb4bEM+c7y0HzAi/Kpld3ZwO
85cJZveln5murCqUStYNja2iwLlu/aJYhi2sVc0SBmv29gFU1R6Yvo+ZEcstsSwkbpAOTLphsj6/
PeZWJixSJCj1Pu4EoErbBtIOSYHDbSAnTt3cI18PGXKbbG1E8rwhSfFGhsEuCxvZ4EDPhFANKPTX
lUecs29TntQqrUfiF3lE4hdotsrYlcE95Vueriy/M9JflIGoCfrplnAbN4ZUzEkZd66PR5yXzOrV
bZ/zF828RnDjgXONVy50q5PZjQWeS6a68XqRclyQCinPj/SKZsHwJfa40yrmS+Bx2ljxbZ2/0CWm
z2QOJhbgt8tianfvnvt3YckwfvdtlEPPnrcVzB6dSZbxlou+X2gcaxjjGILPId+UviEgbrld4fON
VDwqiZ0O6Y/AlhP1EHrcx7CleCYPofFAuTnb5MADs2bBYTXeSbYIh4Hik04tjJeT+LJ5sZV9j3AS
TNx8kLGhi37bhL9rYYN3Q1th9/O/2zY8n6YCxInCUbzPUDhXTsVjL2VR0PKabg5OQIS8N5G7xkEi
bfqExccbpZtgrYwaqp9Z/lrILffBcay+66EnSUoGrI3O11iJNJWwMRhsQy4rWqVh8pcVxiAC+lmj
0ghEnm7RK8xYpLtkvmTc/JZOlxD51LSfjVcDX7JJS7lokmkZxGtKgYj/gOtdX4G0BjUzG+htt6E/
n1X549Lpjsodudp6N1ejABWXd1UoTSMF/poaqV6Z69WV5OpbecjEOM0pIb2gsfixfi8rl/KKgdek
hl2NnQfYoPqnnnGS3m14hyx863xfeTS9n1Y+NZm9pKfS1puQXG33KSVKWJhBibj/TjSXajODA1fd
+u8P0AAIDv6oOncgZOV1yLMNwy/q5JBp2EZa/DqGPeBWK0vQXoD844ysVOnE8UuIIfCRpw/5g1bi
5SzFO3AoCwo6RvcjSnBn1nAmbn3oPh3TCuhYY4T8QT+NiFOr8pLD7+R/9m1hNExPBRKe82uoFDCd
soQsJyU+hNNqIYnyZOggWjlg4oVax8mVJOzNEXb3LekbQ5FR50bHVjjuxfdevcG1Jlk7WCUJJ6aH
u4KyfKF2crXzTNRrgEx7sg1aCOk1Ux88JXWsOPcWNyOm+2JTJkhCmrLymiEocAl3wF/qSr2mH3bR
H3ZmEK5JGD6mVgcAfcaqTpY/GrC2xYNhaRFiyoA7YXLcSQyFYEARNbbef9AzHE2TvCM+gWQ0JXMd
wuCg8VgfQSDRR0QztX04jAdvwtq3idjURVjg8sLYMOzXD/lgGt8KNitx1L0uXhEiVLGVVlf55/sR
ITOmj9m//krdjba5/dTHSQZOCmawSzalOcmGYIt07VDQ/J+W0b5C4jA6auq1vdgV1cUHDSvTvxKE
402hT7coFAcFpucDRqWdWF5NltXAwmbPTzR7AEHDEvpYXanAKkpwRx3Rn8sUda0sV7QQNNOdmbzJ
xsQdE94gl/tTntpcyhaafo+7yN5uJs3mTCaZU8en7o/ZCnbqnuL05t1SKuEo4RWAXrdMJ1VebzgY
W4b6xI+FesAxSUIdad0VN2xnX3JlMgGbsRX5M8PKRhpW4nV/cIqRWlxwVG45BsrylEreJj4xmKZF
bq9A8bet60gcSyFTi4sVxfo5qcINf0oRs1Q9TwI21g+TF2Z/fFGMHMNhb0SEN9aB2cfKBcGN1hwn
1xz+Lw76/46KNJ5qoZGj8mmm7Q4KcZdbmSDeggPhv0+afm796lxMtJHGHrB9FSgrAPVLj69n/Ijq
7ts+mGlo7NjdJJR/lxFatF2rR9Sbqc341bQz8jP5G6NSQS8nkHsfMrXo20V49BYdibmtVkWr87cm
ZMaF4ZB766rYon45jgfK9k+RSW+mB7QoxJ4eOlf5wqEZ95YnzBYneuWUg0LM27RE8rhV9wJ8yaxR
DEfWKlDOLSMVHeXR2/LH3AgltRYoEkPryhCcjKNYT7o5j3XOviIDnzEJYw+zvNZ74iui6/lufRDP
RXN7wOfoDlmGp11L+xm7kfHfr4BciXmqbxThoVuNvnIw/R3/xD5/m7+h/MVdnHrnWk1ilCfzECxG
RY8xntaeEQBc9OYqgUCEq3i+C3tvp/fClb3dEYjNw+A69Cx4SRKDZ9U6sRRW71w2N2o5ml8JJWPH
D0D5wqOExbXs+fllXXlmtF58YPmdx67fvSB2vFBWh6RnrLcSb7e6IOoQfF0zsY9wCejDimG1mMgm
7aLxpJCZvA6/7b1x9jnBw6OfVOpQFnK63x6SEjGTkN6ku2hYC41kqhB+i45xyxroDTCb23XWDx/9
FZc/SDsGr/Ko1kOvFVdKqqQV+rH+S65TutbkQltuuWRvbSsNhy3FHa7Wk2Dg3zBXZQDxqM7NxZC4
UAZrkOlfe8558BVXiNfKL2VvoITKQ7xTOK4YrFo5T2BeYySaJgP+jiTG9vbeR0qtRQHe/NDQoUnm
QF4d6eq8ryiQ+9tZmrIMGg/Bjb/YkrHbIj8Edg4+UPdS6r4IK7ThAbjDN+XqzFkUDCiT9cRbxbnl
2FeHvByIwjOU/CtR2o26MHqqJvEj6k2zhxUe1P47qRuaRp5eutIEJ/+m9FD2nG5vHyiFw3Fxlcqd
R4WL1Vh3DS8RPMje4FLv1v8TBGS1UbF962ns1whyCY+X9o1A6HpbJVVeRLKhL7DWt+lv4E7cCzSg
wX/Lk2J6NCd0/hs5EZnn8+FI9pYwFur/5DorCxcfLf6XQNSBnlnwlMfNyCztjD/yrpIAMi3rh/vq
1XuOKSMhRjEweuaXicp0mHckKntsLo2xNjTD6eRK7jQPcJi7GGNOfUsXY9oI75JBwt5yvZ1J5fqY
s7ij+dVq/eZI/aCZApAKmCblQRkhE+TjzuKAg/QrpFhIW7d/1KgFfdt88CuKuPgyAJZJ0au4Lu8B
8G2nXe95qmq7YY5/2IRIhzg5Y3gJ6GPyevkT3OyeRwsDm9FvFZw9W5kw+s493qRu5htSwOgfzU9/
YdM9FZXXsiqPIE3L1vk7AJ8Z6dNYvpnX76Su4dUvdYSEMh2PY99SqJPm1fczYGF3pTUazG0EX8SW
22nmMAOMlVlMxYakZ4m/xwPGXrLLnadaEFe2sM9OaI1lvL8EECcKy+5npmCPau0fRRUOSSBFY2Ru
2sV7KX0N2giYcDVQ4lFAysHQe/tNMCPVbn9Bhs+7D8yoPfNXWHM36LkCmoJcNousGBaLbMMSeA4X
hmsvEF5NjmaV35/CbJQkb7CTtES3e+11W2bqamV/DVjCYjgay00Zwxb76moS4U5TlBspZS32v+jE
Up1LGctSXccBASG+dIw2XhPmx/qt6Ca1YiMnUy6DCrixCJ5Cln/8+J+xov69r2AySKQfINGeUQjD
NNK9QRfu4QD2ArhH8SkEC7kZWUEjcgB1+4RE9koIm3xyjaL7prPUZeIBimcNYziL8z50baFgdOBc
VWn9yiLUeABELcTO23HG1FbEYaBaie+OzkL7nmrP3GJ0xSCe4a2AtdN3eMgSH72JGTbcLzoaAkpT
BBWsvCblsF98fFIoQjywJcObHm4ulr2X2IDCM2NrMAnWrd5+Vf0EuOoQVl9LJ/nSOfBw9yAkeTF/
dOU5xjWajT2Jskc2Un9hj7HBIFsl9TxHyL9YE0CtskfqSROzfmBmNY3IrSAl9B/dzKGlYdmY91e3
8VSfkQlheuZ9+m5P4Z6TH89a76k6qnzH4w0WmAXs9NdHsOd21E8WMomAP8MUwY2PmDLKWUzSujVz
VtdxrzQo5w8+W5nWn7SbGkPIqCVCqbWl+VP9jrbv2eii8nVZwjnW+rK3SUQU1GEMfvzaMpBOZTNl
0VuP7q4h2WaDBAK5UMRoaTPY1hCf8eCW3ZIQWmW7nZaDtirK8rIYcmiMDPkChjAP9+47xLeJZEC6
NbcwFJUq3a6SqDLsJJ6wqJrNim8DAUue1daXgE/OdTgG5P4D8Z5lx6GmUj+p7OBpcN+UM2IZw5Vd
RccQ0sBlqJskuev0aNZjXPXkrpEcXUZRc/5xhNa3B0pM8wukbo3KAvr5A/EqScUUUO1+Agto1N5C
W1mHMwuPkDnZd1wws3Gfgf4GD8HQsORRzTCACfsFfztbK0oKZZ7oj5OKVKtjD9kjpCimrFWnzod8
PBvI3OBEJ/YLhpYm0YVIx4nfmGwgLWLJ2o8wuOwNduOkcsAvDDAHjQy2SZeKaiycWBaFvKmnbXJb
hbMec4AonN7ljVVc/vEdYLHqxi8o2kkNPDvoM7vcrl8bonTBFSZX7HOfKR5PqOEGD8uENOBDoTIH
7B/peSSP9KF+AiWpRgG39p5DTsoiFqbbD3JLexr0do1CKg4g2RoPrIT2cLvJLL4uN7bFtSMIPL8C
SrRxGJ/HqwDAMAKAD1wMNN/xyadQ25SPJ7zyOn7fe6yUPnvzvp5VoqUWg79PXN4X4KPADFkrLoHc
6pWzYHYu0180bicT3EpiTB1ZWrpOkhDUeClxmMaomi/04Sq3SZuM1pU3YpkAt/+EH1oQkUfc2qm6
ghGx5orKbBh7fkrCIcE6WL/qVUxzwF3qEDmBKKFvpIzt0tK7Ty8Qlf0mYNIaOYgcHqG2fCYejFKx
wPAp3KLDgVt98FPMBr9/JNKbWwsW2VGkNh2vynmvgrU6jhxj41gojpeZ/u3N6U0n2vlH/q0xUNhk
bZgdJA1eRP1JNQgZfvkAVz7268k2FVtS7CTgZaAcmIZKB85w6aVWPIakx5hoPu4YBz8oKUECfCBA
W2l05E7NaQMFL6w7csdHYQcRdQCzqfyFWLHlxjVD8aslje1B/FKVe2koftDX83dc5/bAeY4Ka5Zz
3EajwulqRFalVqfwxOpyp3CUA/M+zSqWti5J6XLbPjiCLI+sJla5FsD2pUPiE94GtA9Wiua8ZTo0
U4WU+gvazsQpfKQe3s1rZ8WaWgNqSKxkxyNe9JqheBQshQspKiDWp03rClFE6/mwgoD+17Pc1COP
jBUh14PyAESxaL79Ncd55XLhC8oQi2GmyX4Tz/moL26R0fgsx84ZYLmt/FkIWUmwKncAAO3frg+G
UC+LKjcfgzSG8tT4AM4vtvAfvDPEWQUL/SrS6S01QuQ4aAafHNJyERq/flxVESMjUXwQ4zFZjm0d
IzivfPradLS+sUOzCNvSQrioS5vxCHU9Udo1VmCAQhrSDtFdhORz7ykTmOpa1aOSzyOZyfjfKmNy
G8MQhEOpXNK5s665olekINHl9Bec5jMuKXrAfV7gGrfBbzDN4aE47wEyXcmDhew4FMCLZHonfq1c
sixPR43iQaONkzj/VagEsU+/X0iO+j1OW8SlcjjtdgDw0siwV7Rx6PlOvdA1an+iD2UqsOuuL7ul
KaNDbiDrHWzExMyovc5tRA2rifOSf77C9LjqA86ctpofgaHwBiiWJC4KKxUc+xwB3NL+gPL1suwf
+ByClRg7V7zUQRscpo3Tua6YWGuu3K+STIcX7d2Uaw72Uvv5gd6a+tAuAoksc41pFmR7QCwKTxu4
RmwPLt2IQnRQcRq8uVYXp2cmOJyxoHB16JwRmdxcBxuxkX7ImH03k2Lua8oREDl77imOy23TbnIb
w0ezeHz6hoKFs2lYDAT5DnJvMmYXE/Y1BzWd63w7cwvVkIUCorsABMGssKKMJDl9TAnOIP1M475x
n7FSh6LpBHAHgGj1XoyEmZJI8zV7Ieui3V8eN9Tn45/TuYWU7xsODVCgJeqoOUfDVcQhOhR5ajW/
Tm6joj7YHvt++upTJ++olQpfOud/DtXRy/TVTQbIcgFd4YuRY1NCIxpu0azaZ8uKv7N6rjFGa4M1
PFAG0uhxrLxoA7fFXR2dPdXvAhUc0mnF1+RNUuTe5UCrxXqbpzhLVo+y67Uzx9pAH9e9Gqd9yCPR
jiJXUxwO4QBL5Ogd6owWpQZ2P5iHHuG/BWRY+fQvXIWfQBWwTIKQRyqdSyHpJG8QMEGjYDFsIfwy
I0VfubVNVC03EZmAa+/XM8pLSSd8Aj+cZI055qUIUZJRctiSflK7uRc6aO3owVlxrf8Og20XY1Wr
IWwbomPWj2WXPu0dvfSKqNUdY0tgDumYQmbHbcwK8HrMl9QXdIDlEMcEIACO45r5KgYDYoa9Y1Pe
Lx5SfdkWuaqPtklcJZ66ep6ckQIOxbFtyIPLZdvI2eEid4LYqJn35zhrY1AtGCB4IXY8ULj7RTiL
pr/G9ZurehF95uYl+D+iTjaOnW1cnw31Y0ByquF5XnoQP0ebPN68I7tuOeTDpR85kbpsvX47aZ4c
plAk5nEV2LBcq0fosIscKdbfu61o+Se4YSUjPSU251VgWRzdZEaNfZ5dyEVdO8LcgHzH1rKEZR04
ejGqykURBMy1S4EMnZCD+MD9JB2qgx7i+7ZyEVFjh1k8h8ZA+WwyZvepphakSyAu+bc5iGTqxylP
tzGPKP750/Yzpc7T7ChU0oVCrEKOnhe9yUESPSm/t7Ew+JffFORnwJfu1gE1cWsQMCCVLaYmogQ/
U7e1w1fppob06cNMyz4ro2yWb8fOzw3feGodWdBthgo/YX9kd54QztmZK7w15W6EGfpnGHo50sjM
C4ds6qtmD+xmq8/9jALgeomcEMOxxhzbUwBPoCPI42fYn7zMHxdGOEbWIoapS/x/5Txu6YeXLDPq
6ZnovhO76PnmjCKr4sSrcU3xkZaUxtGpJr4ZG8R6cjh/sidM4YlGS2WbEDJ7wc4j3uOq2wKRiqWu
LtdLiYQSnKjvXNH8p3pcqi4Vf9I8fQ5Osk5PYpcqoDwJSQtOWGyIlZC7wtH1PsWaWzckZcaZo3ck
VSCogVJ3vUovvxeY9DSL4osMO5YH5fan3yt3RwAjWkIS/7Lwdb2QDPW7hQKum2BncjtFozeZI3Pp
f+DXXnrE+Thgh6SXRZa4W2N6v0E8HD3LTUkP7sUsJAg+wEyCAAZmRZODHNFzZm3J3oHYN6TvqHH3
/EmEQAc36ptYBWHkf2qolcldzH1QKlJnSvtiywNrLROwaq1Ucsf6udTS2c7ww+oPaux8A8DZgoG6
0AfoTWoy0J/Mow5284366+up0MZOncH/YU1fLAF85lYuYM//aXnjn1Hrg/hKkeG+mRIO4OfEAoAP
7SJmDO8W2N47M2Vmd14EK5HlaFqqKFLV9lUvT0leJFVYGT+LpjkIv9UTnURnGb6P/e6XsxAJ2SBa
3exQIOPJb4645K23pFrra1xasYvOZKdTUyqX/VML1u9EGcI/GXL4k576B1XE6PUgcrST6JZyTim3
M6I5Kvkh+gA0Saov8T9xNDMrz671EDV+gUG+n6YJnHKpAjGvdYi69kb7hqi/wuRvbqFvjR+ah6hq
+yaeOShXjhyLVGChawpPziWCtVQDDSJWZz7mJBUiZCCqbbLz7OKWYWnd+tuFsWgIx7C5lHV2zEAg
o1CqvOhCc3jdmj0QBgqd2Epgw1kqW7z8vii3SzFIbsQ9KtNUJP0bSxF9/hr+rpwIBquFmgnrvDY6
R63BP74IGmgugGW6YpeUoU0MIOG5Dl8lW77Dn+Fplc3a8Mvc10JZRwUzsPaVzwX5He6C9cSjDH/i
PE0kT1WxNsR3SAYIndFpHXMLlyY9rKXMyLRpCgRIaJ+AI0eNdV+sG3yh3XXqM4xthLyfmrorzrsH
iLaJEOSpTg0RH21vIcH15ibBeGOfNNlre+fN49kY5OsnswO/7vuJ7QJ+GJyJKT160KWrVuiibV8b
hVHIer9Tx3IDWlhZns/Ss+j1MvFKJSiyu2wcEN/glzv2IdQOB3vkExbvMLWu4ha113F/5cACxflf
gJ47wOcydBirahkrN/Om6p7qJwkt3OCXriUm5ss5ONSadViNbk2obbEcOyzB+nonpMRq260EcoDx
SUqMj2d5GD1F5ollQGHXNLrL8X6WRg1iYdSsLpbPg55OwihftAseNX3DNPjvIrojLNgI9jHrV1VL
0WDOhOM0j/yB+Esv2QH2MEai7n8mZydFMg9Ix7NTZPumOIiZPLWO/5dBzCa3mhIsozSlQd0CsrFM
26VLWSkAnUX/pKrpR0V0fK5jJirfgReEmYstyZconpmswWHIk6a/k5G1gEV2l4U2nVFCp1u0NONA
g0UKdQyMLucm4xorN/oFv1BkEdzvI8IVxN2xXANLleOBkxVxkXQ3iQ4XZqo8K+Zudq7a4ST3rdPg
V7bnHJ85JOZ9rw6Q6fKySeNXJzxMQyDiYgUo13XVnnzLvKCKG6yN35Pc14/CwoaK/pOM/ODiM2z6
qpxFI//xvgYJPO/sO7m4BGiOCPHUurmHbmxebB1KPEDpPbtAze27ToUCvlFoZeX6a89VbD45JsVu
VDvyPNyyGhVyasUtqdQSiHTh9IOOmF+HfgLvv16oR1gvyKOFDfnsCpTYNkDN1ehoNsPxSurRUNev
YKOo6/GVeUqi2k3egV2tll1hAf5+uMNayD/z3WuGg0hiEOpESJzmE5NhayHaa56pW/1bvLtWh0ev
jv2epZEyGBYkIPbiAO9LBCIeySpnAx6ACF3kW4n/SwxSGiF5Z72zHwe+6LkYmIYyKWFVyWI9gOFs
0N0zLmrSs3PjjSYgTs3SITOkgFlOMiYNAZIdIUY31cwu8Uh/Jfg2yMBUfWX1ghaLnmdm5tHmSRYV
7c4EVImAb30aDvhUzoYVBDeQilhMCB4vop4fGEENMRUxWNsvZOldiLu1108vJZrxCeJ6DoXpt7WQ
x9cABk/+Z22ghNSmOjRZyapptjkgf1KM6e9ZMLrPDzP8kSC2U3uKMXpp0GkdPPezsp/HKFnJi065
os/cCGPJaj0DzVTyCIFQRR0K9fadgsZcq/TNLTrmbkWf3CuCy7dDzloTMrwrEnqopZbxW2c5BPSx
yZnecw+72anOokdWpa1VVdHP1IsUtVQN2BbhOr1XK7hqMwxY3X1NCQA2ivli9uNaVI3u8jgGu2JO
BqK4b7GwYT8qEkV5p9clxkwf+GzxnsD10RVROxQ3nnhGECh1zwSQMS56/WhXzVDmEg+UroORzxYw
HamzdSD014hKQxnK3vcILPSPeik9s1vnPzXBErsCfEhbaGHUFN5l2pRoLH40MIZw8kSiMzd2DMZV
rc5S1PH92d97zK0RU9cZk/WXZd6qY7Jm05n/ryF1X7vY9uzYaEc8xLYMrIGpO4Jgez0pH9KjaFlv
0oL9vKPL2az0pJvCBIg2fiYJzP/h+toG4fY1Bi8WYTzZM8aUrmOmbS87yOEw0tAU+5qCGHFiNFmy
jwbpnE1K+y9CMxGIIZq6SupK7/dhpXLTC+knpgIztfNaCqZ52qPTDgOTbBHwtCjncs7L+eQaixjn
j15BkU4Lzay/wK3O3P1GO79IXR/rzDjSgNJpT7Q/xTJq2XT10NgJwkmg1YSvYVFXYhFB1pSeSkOR
wWOV6mGZeS/KYgTokRanwhhNTrX0imSdb9DhAiNgPqkt/DYsOHsvitx2uQKui+njjQmvevDCpgj2
lJCsOVrlYqpnqCBGk5kwhnhDTjHY319MGSYBARiA6PJvWGF5wk/94BUIvVudWVVhe9OtwtB3iQEe
yOhmcQBbOlTEtmnXt2wqJ4Cczr2dYHNbm/wGFmQ+Jdo2BoQsV2jI/BxZyShmL2SeRAqE3wm3BQ3o
Id9dJgWbO7lIlK1va8Z5DZAaFqZdqjkEV6P1EzZ119gsBvbCo3Anhj/INZXAtGhCzIYxi9Ufni4a
tN+gszkJmZFxoYj9UjOVTDyKRQA7ejFbSK23SYWKC0cTY6gA2JW8Q9I27Fae1/PBA9kAsWQdalEZ
KpbqrAz6ikrzmoRepY0YkPc9bnHHlxhGv3aHvdVYS9VRrCB8NgdzMbYWFBdNk1ukT1gF4T8dYj49
y1UzWHP+/C6oGqWtnO/Roa2k+jn//ViFhnWwILGe8kAtAdB5Cqvarc1PpHlidLxyPICeHLYgwtWt
g8OHwM4QTP9W6tiE7PuIwD7JK8spaalOQxw+hJjV4Kip5eFF2PK6+jBLKkLZP0nm+alEigXrpcPl
AtFkscH4Pj81VNmNNzMbZLRkijutzC2Mp+EreLrwWTV0TPtz69F+VUCmqINeXpCambTyH9oxv++O
u75D4aa3m8VLYXEZFC2He5JPnFelnZrYGO6XqOmrkM0OS4YBclGqeYFpUUIlUpEZKpjtnjcxaMbG
OhEuE4eDBBx2lyIKLwjZrJ4ZkgakywvzD3nyUO5bvxd8JzDRtR/CfIJ8eTDAN1LjU/Q3tqTKrZmp
FypQEJXlXQtOiO61qxBK1qoO6VxstoL+TNId/lnL46vVqKO9Cr7d3jE5E50QDsXe68lVpXFxnwRl
LpIkEQhhoHDSdgAECbv+71uOwQS7babjpfbmXv4lpQX/hSgNdX/HhF1W1iKpV0gNn3WP1lOPN3/z
O5ZHvJziwPRkMH4cVgri78HoiPlI3T1Ta881DyPUxChux9DQtFOXAvUfxc+odVJEb/TzhKn6Bd+0
HPlr2AsmihcYoXkEsJPQlHGfyT2+CNwVXLP2+6Kcr/+XnunCZ2dejOS3Xd+ub9Xep+2Vs2wyAAvD
BSqWfnF/zEMnonsPwT3ARk1KKTtFeHVbu3m1Jk3/0gJCpEASTbLZqagjTFnRJQWOpAXYHrhwFHsS
BSvBECFHM0B6oYCb2aoZKrpjWJsySFIuzfwEQG7jQE7UzfONvuUjvV23myHj5B5zpAYAVvGnwB0i
3FNJNcftps6eWCiQTyoql7wm0limw1NnJR3+hr72dkfVEIuydc2N2CTq0e0PZVz4i7SAm/T8ooBn
tkutwU67phlDDGp4FOxd+OGApTlbcTQXzofis6O1++4crwe7Pg7jpEBHBmxv/qvTt5huZ5Az6QiP
BvfZFy+lf+tvTBhCv04pbWaWkHOXFzmHZevgJcks1pILasP78GIla4txigyJrb2qp7aw1Eo6u3Qh
1wd/YLwF9yJRGKNDY89xKo50JBCp31/N6nFpUu5VCCGD/zN2iSBqaKrMljAXzuOdvd7+6TUC/Hls
5hvFoSZ9ie9YQlieXiD2Jw3uBhkSFO5SGKLOpvgNRbi0wfvwChgkjvyDo1VneRiCTSak4fB2U9lQ
F7vuLycx0Dqm5dXeiRrpHjrxOsGY0A4Z8SWtZdF+H4oX/Y6tQrdy9S6S+C2SzO4QhVmP+BqvaRl5
M5z6/gpduTS9aNkaKn4S2bol+FDyQizh8xc6oGvBNXFSFl7a0fLGUv6JrVlTycvvkSKJarQjRRP8
oCaQorNudh1f59cA3l73ZPUp5xTBkdiatVbRTBh7QMEqGYBbzgxNk/JO2JpQZsw1vw26pEMm3Yvz
epilpZWxmaSlEzRywPuy7o3oADvYH8Qv3Rowet9q0otYMezov0Bjy2CqwHVNBgpjcC0MYvUX7qgg
Or4IhUxaevL1dlohEzbL1LwEpe8eegUqXCyxqo3MkYo6XoukE9tX/p+xXrz84tehOLiiGo1ZzZ26
cKYeva4uY3pUeHChBocup6+q88giV9eqT2tawnwkJph25rk1dVoNE1WQSP9UEiV2CcDJRMPYNrdj
51QtxA+QiOwdQ5Fv7MJRUvS0Nb+3cqwQf8fEdGy0hW6b7hJtIJqqz07iGYyOSpBAlIPYjdGWdJiD
MCRpCHlQ//Q/FubdFXqtR++AsFkj2+zc1yZ3Wm7CbEEHP18APj21YGKIb1zkom4dUqOXI8AMLxd8
p704J8C+M0/FcEX0lcz5rCWae4P5uTGHA2/AH+ng6aIf7UdUuW+IJBX3Ddx3npMOGfUVwSdAtqkR
7V9IMCOeDvkIVyg7/eywQ6PgYrdSbo3xlqUt+0LOK3nINN/PkwBMU0Ftg0mHQF+jMgKGq849Hkek
86gMtYlQ9do1panEOoC3J7kZELVaOrRPse/hWn78SIceSJbfWNOF+nxxNd5F4Ei2Mwap6BqTONG2
HOVDeYPGgwrUB8bZX33Rn+gzs118wXmgbQ5LO2vJYVeMhhszed5h3sYMbGISNH6yn6BejcENznoC
u4yrFmc1ESv/4I7aoErvo0+UQcEs9ykimLltRntES+LaeXJdAfHGzw2WZU+NOwWN6d2cP0cYoLjR
soAs4E8b9XpueZETqMKDt6UYYwnxUWCV9XylDT/FM4Wk3+rt4LMa4sPx1RZFOlWZX3P7NgeXh8kS
yQeIKghSgyX1Qz0g6Pl1IB5knq40kgp8BWGuh/OIGFRwH47Nr9S2hnxaFOHO+NEnPYz0D+UJQ9GC
F0O6ehzDXoTiRTvirVWTfHYfIdjKkNULcKX4kCTjptNfhl4W4lrJvfBX7S2X6/dpMZhs+b2uOGa9
QU/gHG5gKacydCT2bUKpxQwUXFsONDawyNBcuE1M2VSNJRAwptH0L3CWOTYQCb9wmdK12QhhmhbK
2rp0YICRH85lm/rjyXkzDnu67XLxxyyhkSn1zXsyLYZzRCPWUMJL9MNV3UEPeKgjHmG6qO3JbcxA
XPFIHKII6vKLQeCcVRdtSuYDOYMOnx+RwOmddm3Js+Yg7HbGYyS/FX/cV/KdV08AawauXS8HETs5
C0OskI+iKwIfgybtaN2kgWdy/tYTrouA84lnoV4ZAdA2ae2Fv4DB5qNEa9pIISO8HLwb/UREElR1
YKyzgqbGdI+ZW71CzYM/Ft3406hPEpEqhd1kT5mgYZLmp0mm0zHoGn0mQr0Rlh/8ZTX2JQKHbBuF
aT+QUq2EboukCjPd7jwAOZTeHZe91fZ4oUrM/Mhr9DhOH0GMnPd7ZOEJmeDLBjmbzXE/BTQkIajV
stVfCrk0pfCImpBb4v4N1HykSbI8Ho8GIY5cixUowxHIacHj+ObmQ/QMz/EY1ib04HWMwXcU/LwY
mdDpNo3WoHuiIsPnG8rHTM85cndAzIOsg9ufK/DMXokblgQOEceblnWrb2V7U1f48X9EcKCG/KYq
SgP+o29GAaEW9n8IvzYHeK4tY7M7BQlVeGzToztGpBF50FeKDPDAvgT7IaBlDZWWgHs93t4gz+3S
SzrDiY4rYEmlq0+lvibO4qLfWqTXS927LB5eXjVR4vIb3vVuH9bF638ZZQHJjXqNOh/7YdfKRqIa
s1lboQMLHpHHgCq4nvez3QQfUTqhzoNNg0CBZsSxNQu6HCmIlTtCsbxiaqaQ1CkghMO6rHREKplv
874UNiLI+PWzCbboj8KWiVyhRU3TKRfb4BzognArvRwZNaaFsMwARw8ycOd4IDbmz2c2iUB98YhC
U/E+c7dWR2vKo18MS3oOjtiV5WVabHqloD8EUNkdH3gKaYDEycRR6zsMdnFv4wpAuWjacxW6aNPM
6wq84Ra6J0/kDkvdP4lCnQ6rhDcaiNLd/j4UG2xm9uRxblUlrmFlR3NuPc+h4M6Nc4c+GjZtxEhp
d3A4r0bnFRZ0hoXK5S1udbQyXD+tXul4wLuZEdcDr3qLwjSaRImfvJ1j+c7E1laaBdDl5lm8WiAT
pM/lGgHmICuD+eA4fEHhNdM59oKPt3QtYu6G0DFZRya11L4S2eAl5PMSaZYgz4fvkoqKMiDIGKT6
M4NLQ6mU8IOrxtMORxeItpPBYbIFdyU3wbQGRt8iFCH2/DSPVoLT/a/VvPvZZ0lhM035RSRmvbJ4
cqEnkaANhAn7l+vThFCackY98iZBDF0rVLy5H9aJYhJP1THPoaLUsBtWysjX7NcVDODirYGPSz0W
x0sBHtqFANjN0nTPw/UlsKWIoOiL+UsnDZDUBV2AST8Isse6v4GeONwEZVM8n/T+DYbgd8KoqoI5
qgx25GeXmtkEnfM3IFQMKORSYZosu3A/Mc6mIoJfK2/XF4wTO2wxwUZJbYSMyXtZCVeF7nU731Bw
/8Q4H9k7Z2KbWEtdzX8o20/c54r/3hTvxV4cWULFOiXwLUSqhDJyTCnk6EQyGl44V9Vh16b2PNfZ
PNZTpwHU6adGxLd0exLQ7CGm2rblZ/bsQgeglMZ8SymmzXCXqJqpcYX5UA60NRSLA5sExA/AYTJO
6RBPxIixzo4dhrEpEgbZIPvbcalzhiLuWCrTPIhaT+ebPzdfcd2Ift5/hit64gZpIEzrYWQxR4lz
+0sPt1/+XAueikRilDVOV0Z4Hu8ycOmTyI/sDHHEErQl5Y+FaGlWbIjJ7aigxaFAVtT4cC8JZj22
ojStcFDZYqGnbqVWXvT3PKpJD7i6BU1bSznpLHVViYGEwx/40mzgXNaLUgj3Q/Q7ozBonzttsyeI
EW6jW/syq54q7f79Dt9Gwv0qu5vLOY4uxWCj7W+CJXW05m5bWcX0FhdQg2V4bLIQ2QLLKu+Wdkde
jtJL8FIJZVu3snYc0/pjhc1NMsRC+c8aTXGKfRFha1mNcs5iQfOks2ko1mda5/z9HCp1XpMXfN+0
bMtcVVydoATiZLEGP4LbRykWyylydD2Aw7sbGFmUQSgL3Di272RsMOIA6PIVSAKwhOxOxwEswPWi
6hsSPQs2KBVqdjBvSmO52jrd6LKNTR88ACf2vC+nQUGy0JGkYM6pJy4As9078s6Q8oAzksRZr6su
Nrqzxvbba3DBB7ou9s6ETlyU0YJO1XqzZ2o8W6LQ+MDhUPXaELHvQhVp5FDIQimu/2fVv1FG+Mha
HfyIeF2n0EYNm2/rURUEc07WkB3pqS4FOvbE4hUMrijB/mw2bSWy5FlOUa90Ij7YTxKK0VjTaPpN
yyGpq49ZCRC8DukbZ3q7dj+E5doKRdjIQlYsJRJNq97/VFotEZxaUMmcruCrjmh5Wgolngd/JyYZ
r8uNgLUHjiuOF6c/m+7r3rngnqGgNg6I/QCu3wJ4gUTl2Ms1BC+4stakXTljnDb4E4aHK6v63/BY
thKStPv0TVtkef1UUOc1afWiQoQ+slKJf5uE25hjrVcjVi+RmYmKXjjtrX7OELhfu4sq9xgkRBZh
coi+bj4xx3pJaLbVOUtuUWEW+sb2nG7mst1pewdAJH4HNODDBs+4vH7NlV4mM2uXbrkP10nLVBZ3
JCKVmkmUrKlki4JzTsrBUTTTaVfbLN/PSEG2l9kPob36njDcO/5Ko6g+yo+FrZH2MJVkuHNCTdx7
im/aMIW7nHpPh4ughzoKpiM0vMbQWDTbGGOWF0lKe5wFuksGaQaAK9H+Ix2VpbPG08pXU3brQs8K
BYmbHqXa/mfLdahxavKQs5oLbPFazY/gPL2HEQrytG8KNAGh03PM09sxGBVZnTtrV4p/rq5DFovH
Bt+rcxuf/RdMJaaXNinXEewuMZfLsa3/vAvVwwtbRDsrJSPjwIluExKcqxn4WXF+f88W9ZaHXlYO
cQJDaXOSN9vfbhFF55T4Kpck9VtbYV4jhKJUtZXP4Lux/V13HgnFajSgf70zyT9bJBsS/pWhMCUX
WyjMXMpcOGbz+V/sap5AnHVoAgwZFAD2xS4UbrlA2F12oBJVm+tnKWgqe8rp2MMAjHRkYLC6zDsW
idwkAXrmvfZnLEM3HYgoksMge611vFuBqiR4zJptOtf0xnlb9nwdypkiaK7sakuyZojimQchA4ni
9M88Pgb/RkKvCaRSZXgNziJ3n5BX0MDq4//5sUWe5GLCTIxxHk3Z8uLE2j1rVSegdnnKn6/YOZ+Y
gZVoPc1XtHUYu6Bim8O8OgagZf1OZPaKRArm3oUwTDvciCMVj2DVs/ohwQ5Lr3p7W8Zu4l8SX55G
JzmouDk1odKV7CFArX1kWT2pSYJUtfbWIzo/VnQv1bOv0T3mft6HgN7qZtJPBXgLn1CpC/NBsHjF
LCP+yxm9bITHJptE+uHHJ5h0ZhtDKiYozkPFmqEmNrt0HE2KmXs9cwpThXk+jtWLoSKd8CQMh7gH
XjHtZ9sWXren4xjmj57ALnnDuv9bYyfNxXi+zNANyQAp6yDSf87cJ+v5TufnUUUSTgQEL75AOeMH
7OVOAfyZ30DCWy02cBuLpBJuSAXQdxwizPGF0Ezd88duJGOQ67HwTIl/Abnb45SQt1EbBbvJrNIA
762ESAcucHA4TtJDQmqNtvvtItFBGytEX+R0Z4E5gy0xGO5kV3vFjXiNVbfO/CcfsRyVdBQqJuYE
5gCiIB/MpaHjVRtYUNWdlTjckwBIjr/bcFr2LXRwpcZwB1qqDi2SB2tIxEuiQBwN+WhPbI0NnqVb
GYTKf6qux5adhu8V11DEl8hFR5AEDpSXziGDiOvfnoXvlrhcy9BWWuN+r3uhyqLr2GNPVaMcwEms
pmoDmBrAMruY39j/E0T2NOhsvDqte4co5NI+B/PH+w0U6uxlSpr1vZt+Ry5LKjnge3wQtI8na0um
/pqPJDKn+shBQHuHsnc2NNfNCMgFQiCy3L6mZ+8c1sAwDatLUyVAxR4ZpcFgqhnHn5PXTcFJlLHb
XUSmXr/ZWd7W4TMoUWaNpTE9g5RN/7GwQzf+iYmhTT+pKL93AiyCj8BmpkreQIl3dvoG/pNMAxJm
PdtyBHmgcSO39xfUYKYCld4pjnbMwcYHKMzpQdQFbyge0ghf9Wamd0Z71sJF0SAZImpkrIyZFYiZ
qukyD9ZpJtvbfjlPDId4W8uNnyr7QYkXchg4XbokPxIjFm2vD6fLPJBHqsdzbLC740Iy7xGrIxNU
/yu3rLO9isdur6TIuWeamXEszc0YDeaW9KHcGlv8x1TfC810mUlvswwy66jkY6iTU0D+Bbf0imPe
PNYTGMnyjnrGEOIYDV9xH2RE4sXUxVpcrcKAP4refvdreJZkMuMdzmwKWujS1/vVCn9uJVChMvIA
efTXsGOoXOVPfdBB5y1wn37oMKNx7YTIR3X07nCU6sJqzeEJGH5FCxtFMjB4DOENRXWL28D78DrH
wJtv4cMkRPHfy87jj5n5iJ0sgkuVQ4lU7Ic6Nc5FLQh1lcszfoZZBoB5PkYrSwXOfcHwMTmItXyh
hK6qvRVOaZAYIJk1DrtsF5a7MF9jxpYoZDSn+wMlCqdDsIccYz/k1lAs+wd4hkQk9VQpkfQbcbSK
9yFKRna2Nl9SEPHfv3ix+5dKf36SuTwoKQK0MbY/6QApXIAg8uOI5VYAsN/GhdLLF11YZ8oKGmgZ
TeHqCMRVekLgIsCgwnpI/Q6KbOsHBeKsR/6X4bk51GOoUKXWXNBn8K8CGGrZzs/WMKY5Rk9uuVul
mE4rRkNsV6bkCx35DH8odjNH92R12/NVF1vn9BspqxNCDnObeO3ifpmlMqW1LVfVDbuYQ3f/U5u+
E9Q9DqARrNvv/uKHK7dX20AyNspOzVl/ieE6Nl/upy2IXf3Q5zYTj08g6ES5RIfbWF5IlHYOZzB8
y+b7QeW0tF8jdsvNUaXsnjcI6yLn1h7Vj5v9AWEWpjszjLxO402x0F+Ez148GxmHXdaWFHdIyPbJ
DwY16U9HzrT9LopNLGHkyzvqAWcjAsdZt9XGyCZX6cqGWa8IYOTUKEoXvUdUH5z1HDh4iwy5ZBpD
OpcjiOcoH9zwf3YGnzDwV7umMxRtrDXKdg9p8lcCTMZdSfwbP1LB5KFyJZj/E3KavXCX8cRy3hrA
JN/QRswFasjA58fQIx2ltYu7L6Wov9kGXC6VILuT2EJWTHQZ49NF6bo0voFa/FNdxamwoL9n1sPI
g1PnmijBYjvhdOdoSymabg3MDT08X4L/skf/8Stoc3GS2g4lgYzphi7jnGd9D/rau51yDfot2ac5
2FUOZ6GV/1DmX1Flt2EGBxVo6h+Su7vU/NUgwuw3aXuAjjTr8yrW8o3Zfywvb5jH+EpWmOXc4ZEL
SNyh7VkFSaMqutB+Yw4WGydtpk+4weyf43MGWnG1m8Yo5cZ7yBr/LMTPtA5ndLa5VSGLXnezG40A
akLiTknx08TNzEGhHlvwNTz4FkH3mw7Cl0A50icFgC6xRqlFZz5dy+N5qGdVf5inxATptIFy5ZZe
khQBnD7QtwVa1bKtanZF42vH1EPpr3ZEhxWe7u+zVTFuVjAlHgcYnRO6g3lTStZveIzcsU7NSlvw
ITtqtf4v7nD8ZQc1CXaoeq7vY45wq6fMCiGSAbhfIQi3t1S00bPhQ3xuC/3z/euTLQEbDMjA4Nz0
3tW+w2GxBIDNikpWRdP8of0SznmE8PkMo+jstaJr6U9rcMZV/nvwJUdW8XJpJOD3ZkhybFb+20Km
vwZEXYlS/B7yjURQhORLz3GmJQfL19F6hzkQXZ7K/8TcjTQa7OA7lmuYSP8hpoL4XIKkvfRsP0he
tbu7J6EOtc2B5iVl/R0/oCGE+GdgHb0ww1ewODinUDM+U9SvUk86qhFaI04hyUmOERT9SJGGt/a5
I2FZ3mAQ6yQYYmBHU7SHMyxvg7m00EMQUvNp9K03Q1O5OVVBsRx9Gxmu/guEFbCzmMRCJkSZHwMi
3KCUg6Y2tk3t0mCBkJLqwhGgWLAlDNMSPgwalPoe9NeeeR5bgfm+URq8E4XepLDFrPBzqK2yrByb
zg8O0pA8gmUYMGDaY3edGLvgEYkMEa0J0Vb0rWcl7aDAXUs/3Y6Cl0VDcKzQOgKnXDW281sSzljg
oeVb9ZnupZE3eS4IqpR5TCXGcFtuWqDBeflhw7HNsudhFXQ5SU3r5dgPGn5J1XaKYPfhaAnJGLWG
CoTzNUt2bxEf5Ai00S6XI5mZGzWNqKvO8imWyXyEvAsjG9mHCCRjbkGSP6Rw0JZy8+CI87zbLza/
osDp6zkBLx4fBZIp9QjaUiCFg8gPc1xHzSCz2VYTBnbA9Kt8Kw/AS3RdM88ANT0hBIVfV0eGPnSk
chIBMAQPsmy0NukH/kqsOiR99AxjuusDtWU8yk3FMD/WgW+NWhUAyj9VXwzDk5MGcmBmKvzZilVs
zmUDGgqL1LT5jaMQogkEydZN9q+CDmLoZIEa4KNBGRJkJln2vKcLbrpN9sKlajO03zskzhm+0Uu7
9nYCdWDj+d9VszEUFIm1t5kGinuq2xj2hS403V4KFxrMT6mPuPZhj/mMG+n/hywbklPmukX6U2tF
f7pDcUznOd5zF7p1OuwXUR5pssPszcCSuKN+XnplD3UB+RvpOx2s0iPeCZasRr4W9ufzi3AyIIkR
CcLVaLJa6woZeMqnbGHCG3+OFE9myQLYX9NQmKWXormc/xiNVHVdHBwgaixdp6w3tpbCBT5MOqOK
nLHICYMKWvSuRJqNP/dFoyQyRSyhPJwWywI4pKHwRglY3yF+J/a0DCc1UwsQTUqAnY3AJN9eFYIW
jRdTmg1aqYF4okKTb+T3vNPSTEuIhG/hoOe24iMRlgiQxtxHf08YS2pVI09+dlTG6v2/Th/ijJlV
pEJphYg+tY+ARu8GHvk171CtZ6ekI8KlSARNoAulvyzuwoDxQy2moc2G19VVHDAxI6HdEWcFcpI+
gtIaiEDGZFQuUtwwdC6MqamxqzKXyj168T52vvUGPhvuE0t+n64fZaDqwd5OMX7+pMStVB4Sno7m
U9TstMwYweAf4sYR6XtQ2kRjh6IOGqYbuob5gigPZk+VxMsJzkfMkpwu6el5qoxj+ZHgqngRHy3I
MaoziEDOFmAXQeC1eqe1tkzSUTtnMlF4EkhS0u6LhyHNo/O/aiFWxCQF+YwH0EGjT1UxiygF+oBs
UTy4RQiZrSvOwOjaGIFRhPrZzCtcGo5xJ92ygZNtoZ+SUatqQEjfjIyyC9I7RE4fSab7dd/RBUvD
CYu2ZvoWzO0L/UNNneRFCVO36zKEXLLbDvI96z44t0+GHREXYeUhhu33RUVcFD3WIJ0KA3EG4gtn
uD9zeSF97eVh7yJSzNUUiPN0AFca++c+AUOU7y/1GfIKK4Ifufpr1cGjFX6//Yvqp9B8fERd2v+f
ZYA9GWyDGFV9FK+LeigsWRctMEra8LfUZvDGIxAxOT/Sk8l+QGpweTup6C3Qz1lCHY2W4sndWhqy
44kjsUrHkAfoIR3j8y9UexCyCph7R6FQhOgie6VXVVghvUXUFgzIOlANmUOB9CQ68sXi0MCoDWtf
yCcUeQTgMfKgOM2vLPw19jtO90z6Cf2tYCH5sJADK2ZUtnN7A7B1Pj+vq/FxQjwH07l/TYTdoIky
GlFJgia0Xat6cTlB5hQ1bffS9Ns4hq73nL29UmUxn8lRRMP8OK1C1iff18bbXq41usfb5f8eBfp1
T3zcNekOZLSJRco+6jJZuY8kEp69/0TtFvNgqBGvk4e6BOqEebToEWVWdkqzkmOIwrQeuZWHyHRr
tWtE1DJ5BEvUB2hLU+RSEHBCfxdzfG1zSCtEnJ2NekQ+nZXKwZlvrmCI52usnFFSdXyBheLt6L3/
l1zsCRspFGMG0MiEvi/6rZtsvp7KVejs3CRcJcPnlJ+xGS5kYIaI1yb3P2N4XuCFm+2VQJkixflY
lexWJrRa8oxcs3uBLeI46Pf5oPXm8G3az/rWu/pu80AJicq2idHnI5FOnvg6+5/3z0bkZouhZcPD
9BfHIp7Z7Bll89YO9M0zYHMPOJ3Z78Rpz1Q4A4jt6CN4fYB7z+GvD46F+wCovAI2g8L0RW199uTZ
2lQz4jT2vPWOAd8iCZVTRVRqKCbhKLJwKzEEASVF7j+kp+Qn5YV4wTCwXxU35PAO5s4NWTFwir0N
rPW5eojM1at6sKG8Luja799eR/O97HrN28Nka6PmFmYamwCNMZPP7l/HCCnvc1ck1YnFVKMRi3VT
OkxXjl/fo5JMHF0xLoxC/JoOstvUa0ulEW7bB0LCMjCQ88oEVPGp4+eVsgOPvaqutOFTzW10lzMh
G742PN0wlSCEgW26EY9viQ2XmBrfXzy11l87+LhKyAisOmJ8BcOS5OMbmwR0uSuqcnW3D8uDqGc/
RoL+4h9Um5fwbwXG8Np2zLAXmIUX4KM6zEKzYyrAOYb3zkQ1FxckBiM7L9yOTD2Ply0K/bhc+X14
+UxeRi8KTWIOB7RbfmiAXOuZvEiGnKIe4TuTsZJR/vFm9z1YLXKVGJasL2DR5KKwXfWoAlKi+KPZ
wSoEylqtmh8gbsrWz95+MgyOw2VEsqIQd2tzji8pK6VHRALlkxJHH9whXGAKXt8c0wnrYIW6rfdn
5211UXPaA92FbnexFeTBBL3sY3kbun0On19GRCUivyS4nTHy0eMIO+Kb6uonYTHKJN/uM8j86qkK
9uIQE3bxXkzzFNTMkCXiql6cPYYdxZzDrUZ+V2bICLZKpN5Lj4ek9WL1aX+BwEpDlSyJ0XItzsQy
LHJUXmIVc3b1VCWY9sxMjft/jpMgNKrbD78fMxVWKA3kcK4LrWivbxQCzZSYSOu4w99uRUe3wu2W
imxA2njnHvIchIV14AC3QiJXBRmo55UxD95P4AjdiH0Av1T0RgEUMlrEh+zTxsdmwt9eEDmwW7Bc
KybJg91Uxfyt9+MhGiGwDWpP/Vj5l8SGmVQYXn9KMmlG4xqlDN400guEoyjEtfOW8Hzc7wKUEbrZ
RmLG3N/kTM4HvcybuTgfWhHrhVHobsGg4bRlOPpsROL/9RXsT9b/XTViWCap26IH/nySdQ62/hna
Cpzl62rxoq2Gg//5Xu0Qbum+ZVZhNzIDkwVqE1fzSuo0G+RzMw9+CQgoVSI7+qgzmCExs9reetBj
tAUeB4RoWHzejBO9EmohkllHhDUgtlHWJ0UG8A03BbRAyn3uu/gg1d+572dG0ORMcpyKb3V3+4YD
cnXfMeRBoMmrNVFzuT+Xdsqg4PeWj3Z/ReKfrH2/sUk5e9esCBNjJ7di9UydvBqHm1d/USETx9V3
fC8hfLIGtgMgHDMdMUTp1eL7+QJJKJCCww1ye1raW4BzjGnZO6ZXQat3TGJhJCKMWTGz8nwUKXXC
dE890EcR4udksh/OXAwV+zcOgDBiznSCk88tWgbwG8MIuTp3danH0vrwOFP3v/l2gvA6+3SPz1LP
qoDmIbQ6Sieelxi6E983FKy2gBKhoXKWWhk3PFxNSqwEVItFrI2pBrYXrvJnygpc+EHKDQMzuzpQ
cEmIV/NbVqRi8JZOIC4aJf0L0dKMxufXxMuq2bdS8KwYVR78FDdfQZDQ7DjQx/Bd+RA/OzlJe7xT
emRqjriKIxxjG+VeXsSGipuJXm6dx5d7Oqv0RPnuvfcRyCsHi0IQkXfYng7mP7OXPLCrpNVLdBPZ
2NKPb3r8t+wm6t8SCpSDepVgj40HmApdgU9+Q3ANWDeEhyuUzopmcnS5K9MJgRCtAy2omdQQORQw
NPPe5hSHyVn6D2zNRPEsQQBbLILGpL815IFqVACxNVrDaFB8VSWSxINrXRo/JeKCoXztSzb1ncyq
N8Om0c6CboEDeZH5rn95SEsGf/rZZEFmnlcRc2dAU66FB37sdviIiUN75L3gWQC/7xBpKnWsXeY4
IbG04/b+GQS0sPNHqR69RWw4GU5gww9irFrUZ+GcOomm8hd13HabTUic/xfuU8LeHd7xZHkBf4zc
lSgAtHUf6NwkYlflaY36pqCOMcDtNo0n7uK+5D1+g+3UbmvMkwHOh6cJVf2gZ9pJzLWbV4Vkd8oW
MEC5ubMWcdcuyOfiwLIh8dChjEN8B7aW84qKW2UnrCIMORFeX0aS1j0aIMewwZPDCRxZxFfHaNs1
c0HgJHImPVVKHLqBiBjgIgo88U/lYatOYTmR+PWMHHRabL2f8tfMvllw5Kzc2EZzrBt2w2HrPNG1
pGOqGqmVInI6fzBLx/wxNeK8NT4WpBMISxbl1GueKBuGxqTSWFzuaS7+h5+8nX0HRfESZGBXoGYA
hszAVCZq+h3ZeYp/brOq/M3gskJLhKJSBt1u3AngI677hnxYC2S5WhxE64WVB8mulB21NquJIpKA
WqOQcrl91aQuqbY2je62jt6uX5Sx6zghNe/Yq9dXU286aMfUbFkeWscsSqfYFRtYPVGt3k+pigJ1
zbW5/USTYxpkLpJAa5fInNeRgpmgp7NzqHpXeyWA2qzEG48tfmC9Wdd3rHj1qmd6j76jfWTr4elx
X8qUpMnLgFGDaWjh2I7LF5s7lV1999+6sm+Bny5SlM3knHp4OJ0LYMIeu65QFDxcly3qSQb0uGkj
DmZn2XPDB3vQ3L7EzBwl4k4xOkcRyvlpWVk8W0PJITHREFMRDJRF1goWOTa04a59wjnc/mm7fNE/
pcBSbQQd8ayljcElXEDkYUf74c0cZ0gGTtaG1OvkgFxJJInLxmxpELm05VLJNQ6ejv5vssBu6rB4
DONB7FXw26DIjWZ1jcPoKBAOO1Lf5xQoiohL63oyhI9caH0tVtXGytXyJHHqpsDlHJAZM8WYfBP9
Fr/k1WFROiQwE3fF/POw9j6Vf4ebONEFazUDmfqR7NhM/spE+ZTjgjSjKU4EHRVQGXp6sD2QMOyA
CDuIDgs6jjDPqZY699/p4ltQX+SiKmkmzCq0+uQ1mlqoLjo78u5exrkefgFsJNkkkWaZ9ZlKcOkd
Z0LeQkv2px8ObkoVSkCwxmg85nPlhXHoYsO1YG+R+mcaN5uC4kgxLucwu2L5RpsOzODEuXXP8hKc
/0c+pkeKlyBEKOs0u12nEdbVC7LDhCbCDNrvGZY1CEmPD8Xj0oyZ1RWhlOSxYF6PSxahra8wS9Ty
3p2B/oYqVxR+EJngRxHJ/z6RXxpnjbComZf35m2cUm8zh52Xgw0JF70uVohBJSJxQMfQlFvNLfdd
XWSno7yeTuVu1lVV2xegrLCZHbZkiSaZxj2rbgx5ANEbVbkqXZlBzzCw3FnMP+/+6T0AJ+6T1XNm
IpJ7npspQJiod/iRIjvsppit9dU+41ax0m1NvriLrJdycgtZiagPIcPSqvgUN+6UbuydTZ9LNK30
HXEMjCMaSDahLnAL7+sBFNFshGcKc07O5CSNXFE3dCfdRIjUDJ6WBEdJHXuCnpCR4PCCg5PfgNDh
c6hqDtuZ7kSUWVqXIiDyyqCCEWhzuz22/XGfyIKM0oEadFYqGnbblkKltAs1Shl9frv0z7gLf90d
7Wo6LN2WkxwbObeqE3JRphnY4LCyUuc7C2np/bLMlBJsKV0CuROIPpODMfx33ABDAocmVpeS+4kd
Vo5S5TjnLCyqOx+WmXlUCa6oZDy6bJXabqKyBB2pu14C0Gm9fHETOuAuOTNc0TscVIZFA/s73zAG
Zbx2yRObr+C9mdveqdLRMpvfwk7qKh97eGYzDN1IM7qq0aqrm5L1F91awe5rN2dYy5bPCRn43TnP
Qi1LE5XrBDSQeWHCK/sSrp2Yu++QPf5tionCH0VrbOUQ2u+Cm6sFeKJUV9/1IixUYqtmc8tWYXxm
Q7n06NvlzPeg6EKSIM5JfHv6J97oDzwOqStZHj8EbmklHT/sFdxS2MBQd58jDfFFb/tgB7Dg43uJ
Wt8CjKba1wPNCAmhPQFcO2cag5iP1yqwPfjRjNEm1uFcD+h6PLp2BaawIhjNKSELjDICPDu37ASz
0bp/G55Ndg61E7HtrROgtLRkAGsWjcSLKjjytvaQkEBSaKznKQJixwlvHt2CquB3Pvevy7CkMy0L
4M4znVKdFha2exhVJZbrjDjo1NRABABBvkHAiq9+SnZAuWz0BqDv5ldml8n6w9m2clHYGsjZ/qiP
BzKp2MvFz2psyGk+TbgpL1bjtfG7ZJxGuvFqexBa7djrtNEWgTITaANhutl5nbyQOlvXBfFJ3NFb
oJVx83Rs5kT2kr9I+uvXNgiduCmXNvFp/xr/ooY0ty53JgfgXcAWoaLyCSAnyVwMHqPBM/SAC5DQ
JnrIvKJsPN8uVsOHci5hQAHRm5/b+S+Gt3pB8LbGeqAA10XcapZJZan+Ux9LM7+lEDAGIEXeEOnQ
ffTgyuV0jc2+GwogNmDEiPyA1/V0wNA3BNs6LXzHpnOJr2y10wWkcmFRE8Nex5GaQn7e5TMWU4+s
L9yQC4wN/8f7pyus6keA1trrkH8+TvuaXUBIKsHo+siQDe3BpTEnMlU/t2AompCuGM0AvFuYlZJI
e8qqpByTd63vLR0Uq3MS5A2Y8X+7gy3FeiKonsL3TOxhj6esp0/clQyehY0CNyNwAVrzM9KOqGZE
IO+gI5+r7XSziW76GsJdzIXFjKjjeapQpki2zIbNs+RXRxwDZ+sIvahinz3/fDnEazIb4KIk1UPP
R1SA4OlMsnHKx5j+7ein6hUUziWF6kZ9kh6I1GJgJruPLqJ0fLMJ+rLaEu8G+HPmRk9lDiATDCf6
5UXE3m9MeknVJkF0uTGTIv+DRct9NNXf2BFF2F9QU2CPue0gsq9BhVpUQjrmbh3/KfDye80WTckw
TxObOmebLkEBrrQGYfvBzCkveraCr53m8QSm7aTvgGR81do1+ecJvBl4w22P7rDeBKLXria7zZ7R
yzf+6SxFu2BvnqkCqxoXI/MdQqpC7zX8yXcH1Rart2OewHvre3zVfaq/MRUnRJSbDKNryKB86EFX
/2XJts19UQLRjG/mGYTUHcz3IgE3tMZ3RSvnrRUVcr58sxMDsrYy+tdskJPJrTBVhTbJRorIB+sX
KNafA6kTUi9MFcYRvdd/iTH5zXxAQWsWrsbHvFE08YbsWAvL86kWzKVehwDyWfp3/d9SLlg0NXie
6bBOBU4wKrGDXjKbY7AAk13ByBrUF6TrwPoHQ3vOPbwbdMMhHKiVtora8mxeiYF1DEoZtjJD8KNS
mkbbJWv+Izf4SMCVmifXnOhDjDtNFejJHpozizwlfJH2V9ptkdy6O+SAs4p8+nRObfajkIZA2JM1
m6Kh0cgJWvWc6Mj+QY/a43hXSA2ju7upvIGiYUA4x5AEJjMxgPFwU8UvKTmEf97yRoSH8Y01kZ8+
7YLOkmnRC7FAAEXQtNBj1yWkJWIfiX4ttBKQVqxJMpIAMaSMI9jM4LMkTyG7q5TYLiAsd51FnLcg
cQdSdBtK87FWrTV23oB7uXxJvq+Bh3k68YSP9P0xIZRC7u5u5DJ2ZQoPPBTX0fptZo+MACxHICD4
aspGfjyYd31GIqBSrspAwS6XO7pTOmgL6sGPi2abtSBgTDNGy4avDHEMUnqfoDE5NGsT7YdxNrW3
FMs/M9rL2ekMBX+DSFFWauTXpU/5jD5XFO4PxYN0uXLtKFM2AhBuaFRKVICkdV23x42Px9Q6yKxj
ificbPHJIGEagW4vFBP/2M6oiiEDw7vnDIJrmPRse1/n546sE9rnCJEZaxViUVWg0ZI5YWYshOiY
io8HnF2pqP09NdvvS2RsvXT7iyDEXqkzMEgafZ6CZ+ollxUTuw62QKDdduichv3hVYzfme8rjPbe
Dx/5QYpRiOg1S1vtdiTb0zVzZM3Ku30hzNMY8nT04Z0rHmLLw1IT8UtoN8mg/4o1Ty7FCi6V04mk
ytkUmBWae7SD18rS4T7WPXk3P12yMCZBx4B++vgIUpBLjIqJeNVZz7VT1Nj5Ojx2yZtGE/zVByIo
plrVgTQRU/BToCc5J26oEp7ek6lj73vL0ZC/T63lbMP0eVMfkiJEJkeXUw+/lzyah4v5uIj5UTQC
xBvK2l0LxzbZgOJ3T69ma9gkzpye+Oz6fil0Pa7/cmKVHE03xVDVwzxvAP4WcU59koOSGLFAiXCb
0AM+1vutBpst58MtulWWf+6FTk/W9ey7zJrbwME4AJ6JagVgARLMIEPe0YZtRuse60C7X9fhGAvU
SPzjKCyO/b5CqgA/OLMzL8Tb/kXBUcUHvGfafzHRlTBGZH/cy6Y0J3PHX5bd7cNvDXRC4QinGPE2
qmWtHqlJBQKa5LBlHRIsNvKgL1TVYj9dwfophCwI4F/FD8k/neVjF42crYFTnu9EV5T17TSxB/22
6RijCCKF18qre7vClHI6ka3C0UZtXhrppKxV0NToREiQfhDRp2frv03WaD5TV35OLCP5D2nHVreB
wxGjT/PqjAuXiJ/nBN6fNJPA5pUKT05b0DufPYHaocEyC15MzElyxmQokfFhMRSgkQakXn1QkNhO
rhWNtTPP6WOQ23lloYw74izMNSjvYW6w3INuL8PY6X3kuBi5PSfg6SNpCmIEuYeBIViuqzqiKCdO
1R0cc7q3hO8NNdPcWvPtcNfC6s6goWGOJPqaOQPeNhwIfNee4dDeyJWtNs9WtaSTVpKhUon3fZ5I
MNViprt1cI8kndfYeSw9irqAap8G74/xW1wQUXO2lc3Zn4MdjJ1vQVdUQa/KdQh6Mz8DtRO7YZg4
3kGO0t/1NuMjTLJJoP8v8S3zlUUFdxMfuSKMimF2KdiF0em4/eu59AHauP4vQJLq6pquVta2DwSW
fCJomV7yME4SJN588vEVNFbmtDDH8fXnEsl2mjrKWVTeQuzQ0iPBnEyoU2FJ2+J6jx5WeYcup7iZ
Rq81fL3s8uZqCJC1HfZwS8EkzT9F9tSUB8bKfbRCRqEfKwwszqq4dHvGlnt532nSgoA2uCB3qv+p
hSmMQb1WsAno16dFmS/E+qDplJMv0GztCIt2JxYFQZTv2nKEgA2Mz3OYBLglw4W6N4Gl21V8fqNK
oaes49Ixzff0wVUjUJdEWHe+dVrUSPpy99v2w4KToIqUnRnmv/8sztG0q13nzj2sxBts1uMgc+L7
aJhugd3tKHOO/rRFZYvR+L6bhRFfFL0KD4UJ1p3Zg+sWyoSursUvz/ydb0fFPddEUWAhqZAS5yHR
RsmyD0KujC6lt+WMdueYiQaiUW8PRVjRYKywgwxxH9L30boF8cGiAZ2MiTEgL6a4NXqeUi8P3eK+
uAfpbqKwebeTgAkox3WegkJYg+0herpxRvjOdak/c2VygH39d8zsfT5uXY1hwrPHM1zqtIp4A+GX
RGkmSerUArJJYsmoWSx2lZpL1yiVL/VtGDmqP8GWvGajkWZUKI/Uvxi9qwO+W8eDU2eMp2CTiRWh
oaLq+iJRYmUaNpc2OhxEHZA6ax417h+w1pYEHmsx2hiCbcTR8rYlmcCSmgHVnNfXcTSFiL6uKCcX
TNw9OkTB5zTH7gwM7tHcuX2BqR2y9a0nsKIQr+P71maw5u5eVKocABYkDajtnhqGcpxnX6kAjefd
3XgHhbLFlXtO8f4GeJ26lYRtii1WH9JwJv1gxN64vd7J3Khf34OF48TqIyHLg5Y7Vum+n7ZM7lzA
wpMUm1SHLyiceR7FaCbkhXRiRPkIgMz8ZkYKlrZwDhabFdSc/RB8MWFJ3K0c4kJmKC/NJJnCNqcp
0jCtAOhVJoh/4qI3qCUB+1VZRKlF/lwf9D1NFZkEr8kLs8NRvG4ENlnTLDpjp87QLIIfqr+NRUvc
ciK7fXdf/yiNElFe0zqRBXsCwQbX7gjlNiIqBKoz7gkg7IrMR0MGIX4TPsiDvUGA9Qj8zQLBZZW8
KLCAjrL0QWSAjkugTFKL9HGLzW1IXx0wbomqpv8eMo415hk5qQTOB34Zvqs0TEWTYB/xrPOW/mKB
Zu9tA1e7ff6UvwoiZsf+5/Ha80dNj9OgpuHkluEbyM+JPWP0ZKstMbgLAbWabaaIaRN4RIgQQClF
cnSeJteLuk5IYEX0MGM2JDjXxbU6WbMesKLafpb84N9HIYpghlfW7YWWOzNfWkFICQHovFqNolML
3ZRDYEk6jBjyKmgBsNfmP4tihWdM9LBdzWajQNUPdokB3PGpkWRoHCbcM5iP1zPyyLfQaGd6VtDC
ItJ2CbYbkHOWhhhTuON+O7lEe9SzAJuv+hKJxYH1rxUxo800QSQTagWDGGozKCztIzqkYCXFT56E
T2VpR6tqdzH21QnyQ6YACn9pGmGvOjj8ycYXOxnWUjcRrd98cj1DIPZiA/zVy1S/SRrcECjgxOMV
hY4Y6tYKcF47BDs7ZdRB1nTH1uWO0gkpR9x6/A8T3XNIGKe/EYUDwy8pKijGT97w65QRstmZV/M6
T6OwSKYcNeZt8woKeOQvZvG7S6ZhVeaGuSYTJ3Wfy0MdV8sRBpPevPx4/RGR1zWgz60qx/qNfD6D
XXdD29cqXRtU2yXPKYAy2GeopEM8IVIwbQswtd6jyrTPqx45ogU744chtxOf0iIN8kfPJOP+lrmD
soiYURKuEHt8AoVFNTTgUJgGupPaQ20CiJHkI8Pw/Q2iwDnrF2aXfWyQaYFqCGIT4MYCAGdkdUNK
4HfPc/vItaHU4xJi7s28XZFGT/91T/tYZY34P3fFJBXA97pDz1/IaFmk3BEdKoazjXkHJQY9VSsg
XQWIPDhssRYqNbmfNsJlFVBOM88kwonJbFB2YUM/5ED6i883wS0sHtYNbgiIAal1BFqDYevAEZ/T
kQewG+XTx+EdX0rG3+yJ/kVI3fERbHD8yh1vVImYlEJxgbMDEh756VJcYtZi14JU3S2otYG89Q0y
HAh07PtgmWmExu8ELZTU5QNZ9hCNiXRrE4N1slO9gxcup96xJNZuoU5g03bdbqir4b/L2kZpSBS7
nlYtvaeAP1aUutmO/um9w4syfewdTSvkVM9snWs6AW2m1nM+9j8KKi+p5+BBEoW4skxaboFKS+jq
nbYe1ogcJA06Zs0M4ig1bru31UvtCVIm318NmcNYNR7mqE2ABsNzg/2fFdJGxn+WGvcD1rI4Hadq
tak7n9GLZTXhYLVjhnu1YA+5p3AiKQhsKLAVl/0jw+Gsr5sKzFPV59hFIp7ky8+v0Ka8Xx04ObpR
EFpdfQB4gRlmksL9+QSgVLYu0MsAH1sOYUzjrM0tbkC6h4Ep+DDchCAy0fL5xkhJML0+mMp0whUL
4B+EEwsHuQOTxSQfIfZCxhBZMaiL6i4gFymWaScSCKAWoXtemETuRKI0xtsQkLhNTF8w03abT6nY
gvUvUq09TF5MusjMzjQiauD/WjlOGKxLn1HOlMQjycYOOVwj5tOdBOkcJ50fHEHDvSX8IVYjk5PI
F7xSoNS9hBWuzAZFxGQ34q7P6+8N5nGYRHfHyoCjifApuEnNKAKgb0QCpc34CzG8rPXRLMQIz2LF
rWJw1HuEpy3Wcu8ZSF23RO2vLT6VQmpb0Hnnxx1veS0SvH2+hZHEjhCGTulY+SHSmmUYeBO4VZgj
3B64pZHZuRvlxiv0tlSJ2zRzeGNd+9H16w453LlO5CRg579760cWcTkrV4c4/GhnGeFpMG9EKct5
DXEBWDX9I26vHT5BBl9rmWQo38XFYiRaBEmTdTBfLcGvwJVQcFEwvWUUX5UZaLp5uUPeYDCiLQEq
hpLXGp4AYYBot+OpECgsDv9FR77YJ0sGLWxAJr8YoqxAmYJOYgyZ1EbGh2tAkTilahaK4jfnzdCF
kmxmKFnMby5EmHh+ews4tSwy+FD33uyYqpMGOMlzYYE3QyCHCTF8gCfcnTH9SBNLmS7ioSxWXx4p
bfgUciENruWdKFx60DGVQMfsT+0r4aSEOQAi40TIUlxab15TlgapiFqWgbl3dOvOxaXTdq9kMxt/
cAADp83EUvwQfOg+rs73/uYpNycZavn5+EI9YlPgvHAPxl0g2VDXkc5LAfGgb6e67lHeHNO6zQ3q
c2ew0aCRwdlwjVxO7VMNpUvU5l2XA/h4REupCXApQasDmguiCvHY4TGJuHYZMa6JX/9ShFhL5WJY
30vK3XFu5BWwSWFX8OIKtu00Nzo4bNG1BwmUwze8fSpxGZiSpmx2X7nU1iMA1KeNay2zLiuDyFQP
1KIJxq7+/YaL3FojI3cw71k6//FqsxFomcfaD7WxCUhIgGe8c4XQ0Cv/7WhZYV1H/S+n5c6GrWMZ
6ba7OqQQdK9w3r4KnaoziDjHfcvA6GfCwV2knBGZvIqrayz4qjTmWXZVoa3PQCPHQy1fCoGFE5so
OFKLmVbI9A/XP0Le/GUHJC8TKmxYQqTbc10IRBduz0wpUd81v6TVSZ6IQWLWgT1AVaFV5shHbuAk
PpJs4o/VFuMdS5dE2iViWE/h47nbi/8VkFxEHcII4Abn4UN2D5BYmdyJj5C5chF8EBse00LKar0M
xMXNyr/V7cKCe2rdQy6cXpMvimlLRUsd4318bicBOXHyBiYJtbLeomk/CFG9V9pZyfK17dycgB5w
wPN8mCL0+puhhGXm/ct8bbRHx5XIX8wJiUBsgVIFwH1yE9RFOzJHxcgNfeSgiauGhWo1lRKoo0um
Vsf20x/o9+OnZjOiH/Ueor03E6iRxr/DZmc9lzMpFkg2jF2yOzFdydgchcxS/i4K5AvihowQ75u0
q5QC6Ssp30TDGJlalIr45oKKbzzq4aQ3fkVpr19N3mtNv6uG67wPmI1Cji87D5v/m5683/K6Q3xU
uOw0WFfjkzhTz9uiedyCCMfDMqtWXUI0ujxflwrklQn6bFmpbIIZf+5eRhEqzVEDPAdiriXqu1lE
jqmj3hhb4aadp/h3Ypm3KFk2unYspxQCTCnQdlBWa96V9pqlPCPf+BPimmqVSZDyynZ6i8APr5fn
72woirnDeM2i7ZTQU229+04RViInTl1WO+7fG4WdGt+edpdbuZFNq77H0evLlE1c4iIy9Aw3PfSN
0rYAlJ9Y6UTast9IwN5u+RNBvyYBEA7gvUB9S1xVjmMg0y5b4TI71Ps+ceex0QV9aqbOOf/siAOD
CvdUhE6Dl+Lyn554ta1pQgt0gZFazU4Na31B4NxenNZaZz7NqQsYDc0zfdF5pflDK5J7kVQVipGO
LAnSwOpYe8XosT2KCXFX+haeRBAC/CKnKTCOxNap6wvmupxG/Yt9XWr/vDpjvQCQ06AceeBeOFMH
BVKSwjsDh73RshF3BvX0VZrTo5hWB4PcGGU4pUyNwD9AdxjLZnlXja0xdiamfKLDgfWhak2aoQs1
5nkGYFDBrX8N0xDZLB63AVpPeFRBCAyjhHTm005jJNJhj9vCQEeKoldMDUmTQvgTDe6XRShT5TKQ
Bpcngx/BwI/KZ7UvOFrs1QB3zRAgfZDYHJKu+rMiQ2NiRFPTyUntXYJismxV6/Cd6sTrFBy19isz
z13TkFyBif4iDAd1bKQdImN95Muu7XE4FUpGtSL0yncYQ65oQI6cOMG013b1Mwq7EziCiJ1RE7iI
PZgicXNdmZ//z8VsFxvIDiPf2g9wbRzVACqM5NnmuvNCnp98z3msVpIXYjJ6lFPQLfh88L5LZf2q
j8patlqPx8koB6R0T8RjwRNeXf9rhDE220H/Pt0rC0wMhu8ie3InZNRFsVsrQYrnBjjtH+xHpu93
hA1XgUnOvcKNq7+gnWid1zDDon6Q6TbVlx3VWegWQMXF9w10z7ZezceNp9KViTfLFIr6B9fhqpZ0
CIdHyIOMFfX6JcfiRcTUUHfN1DJymyL5156Ey8RgYZpAfVpqfVjMXCc0IYFTEZts5hoDESbhdWs7
qHmblRVte+zAuzCmO2U3Aj7rQdzOFNh7TJ9fX16DNHTd61HDxpT8wk5VS4mGR6ySb54Fzj8eQeoc
B1qPIfzfWr4ee8b+FAdoPKvenVGbTueVpMLMuv697WHzIX7s8iY1he3Gv/7CzbgmqHobytQbxUxX
9iZ3fKE/GOJQ7OYa5KhHqOIdkcI6MsSG2NFuqw9MKgJkcbWmH89Nqx9a1eZOL3tDopNsn2Ownt7a
aXuWRWeHkqUWwNIPA5NdN0RlTEYKH4Ia5cdaxIxSkBTfkcXTya9H/O+Kz1eqaA+Is3VlG9yEALj/
K+kXgkjjtNZKyfAeflDvbtrZMtydfWt6NYslLJA2BVabTWPRazbkHc36mKwn8rTaEcVYvQfiJ9Oq
2AVZZ7SWO8L9By4SkpVMpL2gAdvSpEx3RpaG19w6kIuWm9xA5vGmnHSYxs7C0YIwsGIMjQTGVWQd
PbRWA89dGoYhXPYOow6VHUgjmiGQhM3HpcFALTFYPQ4m4hImeyGlIyeiXaOaExOEw6tTswa8LdRO
tD1uIs6UxLXu0QjNK/SgAKD95K7v74oGRUdxx/YIdsrJXMTUk4yymxWMP0iFIZZZhxSO4FOFNWiq
OqM+mCw2M38MrWiKsipBiuPPb6qF00XoJnh+DYmU4DnpsRTZ0lUj4nV7QcMwq3QPyE+swwiIJuOX
cSv0PyFQtta5a6bqMznxWlLk6A+Ltr1urqX2bPIoYmAvu//T6JUnnSPcrS9PHgjHvXMZFNA4aJPP
24QaPKNTeq5AWeJeF/8HfyVnirgqGAKIqd61gb7l0IduO8A3MFTYSPLu7FF50ERlmCCZIlIEA0My
WJSY3IR5hr47WEInXFA6m7p5A0XnTpQpFpxdpBVT4NEMO3qqAjfhZWmazVK8qO5ZPJJO86imm1uQ
tK4LzPAyc/3xUrNphqqSgXmMR1ivITPfx7HJkB1vosOxiWPujIHW64BDlQssdvtHL2k9hwdsLdmP
c+kIaY5Ut0Zb7VxeOUgwaCL0/B0DPOCuHsImf4FwEHywutf0g3fpkc4tO6u/qvQR7+CXHdQb2l0b
GHU3lHji5g6Z9p/LcLksK7yV9kBNSx4m9sA+4JoZMNBbTXdCT+8iezh5aXRBUdNm+xpgmESDltXV
WshOl8OL5Q5348ZU+fvS2l9sigXUllFFdO0c5t2u+NLF8uSsPIqFs3bJFXM1zUTg9PGwNfr8rk52
RdmZ8ShYA4GhAgQzvvE6uTeil5Wi+FGG0grc36U2wtj4RC9oGQkD/0jlwff/lzJpkPILz33SmzOA
LQ5nVBPon2aBbe93AgFhoUXWzFQlF7GGtCM1i1kx3fq3ccUCUhIIvm7OQZbKPZlX7TTR8ByxkMzk
sO6Xj4AE4sltLqS/fgmw9A8EoL1BqlAdGpp5yuErUbjZLO7e3+mgswubAbLkYUU57qCTH96vUgWD
Yp/Z9w6WIYyg+REGNf3NbtBdoM8KkKrwfa+Ez7Ch8BeIEX0/xp2FA0Zu4W6Mi2ZVy5MhIeI+gCm6
N0aW6LUdDV9FrxiRKt5vrC7g+MGjB6wrsODkkXYagpa+w5qTzNXEIRVe1RrMS95w163psC6NkAW3
d4sKgY99RUTejcgfE889UzMneGlP0uxEBilKd8kTcvz3ueOItsmcCj14la6a2K01OI0yT35gG/4/
Hhe+79iKkmhGQRkAXFsXWlPTjx9hxPpank6v7mkR2CkjTBpUvQO7a22HjWSQP0ccZ/tWVTQQQz8x
4zNcotlhnbgILz0uB990I3jfI81WWM7Vc+Sboz9u54zZpUe+AWkIgmDBnrL5YlM1ThJWWdnn84KL
jCVQWB4xFfY2h8Hvwj4HSj1vgYL0XxroD4JmXx1JKFzQUo0h5BT5FM6jC92qMRzUek50wig7tuHo
vvDGGUIbCT3Z9ZjY4JkN8K/welnIfsd+IsevMqmyBHY6oR6f/axiNwEJFdsXo3DJ4e9pZoJVPPoK
lSZIvMRcuQ9PNWLasoiD7fdSy/CqKYkWlStVLkI5TlWxVw0BrcT9dseT5q5Lt5LBsq5tOxjr8AGC
ua7pAz/mWEOu3YGb1zzFP4Se/bY+IjMMZeeFb31U1wh1I+BvR4IFyKMe796QRjxDYiMAd9deTqvs
qwiJjjPmk7HslnxBNtqe4qbQoBJXYjap9gSdWQ/Y7hsYCYAEU0g88i4Cskj5A88m/YczdVatwQ8G
yybPjBLtotNiSQHhFeymLPvLMED3VRTYJDWbjs52s43rHRBGVmEjyRlORh1whBbgpmiEJttVpWtB
6nZWGJ4EhT2ZVWx13zQxdry55lPwnT1bI28CmysuCsaHWk619b8+RB7KuDfD4E4/92P/I9GXo6+L
PQC1PU5mn/K0vdqcFSIJxzaP4NJM4w53F+5wfiIPtHVPtGCqjoiZ9oZHKZTHEWXrIL2eL0XOug0g
SyrD+Gvgj1OOX0LvYUGKowKtHcm59fiRbG9ELixnwXicWWwyv5mqN+X4QSg7GQQxuuJuVTZcyBZL
PqJcxxctKKfrHEFig0sNUE/Vd3UMgm85mHN7ZxOm6dAOqKrqG3dVp4IegLbLzxcR9nptWzrINubN
TMZiNsjL0ij66iDrLmI+6CxjUDYPQD10d627xRgti/ODtBLze0VYTDM2ilnJhNm8ginRW3gomFfl
dnlkgJd0E8FGrz54SYwSHXik6HLnY+T7BTqyhtNycoGsAk2GW7kHytJjY6EgCbWDLZi3G6z0xfu0
B25ls6mtAt0Br2TktzDTfNswJtwDmtNGqCXwLTMAxuf5jKvAXAyw+PF/cwrb8fuaYhW7QR0W2gi/
3/U3hLWHknArpnaXas8NV1UIg6iEOLqzeaxTTXBJ+LAH5/QlF0lr1GAN+8FD8EVJKJ3aYJjLoWWl
uAYJ+fgSf2x6N26VFZeh6gG2gTo1cA90DAkhwjoBwTLUNIkX+Vk4VT7Yz1lKZqQdZbSehE2ya28F
Ur3V4sz8l+e554WGMAS07fqMhRrgsTHSyLfknDrmxF7oIB4S9l1bI1nvHQLC59yW8ohX39LDNgQU
JW6tPxj2Mq4N3dycRY4jbPmzJlpN0z/Z9L7VYSzaHvCLyLi74k7NE1xQb0m6/YHvoVl8BHTv0hkZ
kZApaH1yppmUIh3ti3SZ9FFYFWsomZLuodHlLxefjsteoiGRkAmyI2pRnTGDxXlA8ceAUHOKZvv/
6BvT07cSt42u2DFjk8lgZs16e7bl4l8WZ/hXrHUOkoN1HjeN1OAMIVjxjlg75e5cRqeJ0nvGofxW
1sV6I3zjURJNqDD4r1+JJV10QiQDmadv6FD+3TYWworY1nIKDjbmmAH4P6osJc2IBoJ7c5SVx9uK
u+jMILmAp5jnAkBe7h/T2tQc3vbVVwQVlMvuVKkGvdwjsHJLAx1ttiDbkxqwd/Y8rh+QIaZYRSQ6
6uxxASZm0Rb0GINyvf0Mgw4qorIIXdlD4kc/JmMV5J3eRem2b5MQHkbhgXcfEGtDfCSF1ucCH1XL
zxQsxT0j2Xf8v4RVF+qBgzGqbRjMmxaxP7drzVSZcLiihzPDXLaJvCtOFBUJ2p6I2DsVzKCRVi8y
nP9Ogyg2Z96kzwHk0QBKzLgxamXoX4TSA4CNkyCRv9TJLASsP7xYp1KnobCBZywhfkuxVK7RDBJR
zfbDjZ9dismlNJ5647WEWRn3RjPAwqQxqS/iuFYQ3alUjL49P8B0hUS2MR8E4esglJ9xnzoNqD4c
WnmWNuVMebAB5+gSRQuFdDEXxKgIgFPGxD3/zOHMLbxgB4LR+KjdLTCIRQ98+HlnCMSz+9PVky8o
0UIwRQgh06m9vvS3ea1LjI8i4Xl1Ml255Rjdbc878I/SiP9j05Q5taorpmmC45XOceRrj/Vc9UZ5
swXskh5Z4Oh/3CXVk+BYVN32hdDT63k0SZuVFC202XHIijB0l42Uph6qZCahlg/zsk1w7qB3ktW0
38z/VdHjNC+aDLEcUS+gBkRSKLFrJjf1xDY/7pBGYmubvUmZOAK372hdL2IoCDMf6xnbRaUd6+tc
SFrJ+DIa1kWdBYHavwsQ2cePwskoN0yD35BQ3o36tgeA8a66JzxJRgqphtYprZa88xpY5gT3gX2R
JRkChyLXsIpNfVf84p+W6H7gYv93N9HWUYu0fKqdXU774vffnL2WNJHzYEC4rkRojeEQIy1ec8J0
eufnqO5o+WH+HbdJYA8TZqrc+RG7g8MpTr4nXu1aQy/yHKjGL1yq8zkllDEouTAc6UT0T4vQzNQ/
hIPgYS9U0WatKxPKlm1wBmn6uWKXfbGNnrkUFcSZjlblynLhNno7/ciV5HNU/fnTB8f3sSiUFElw
Kl3MV+6HQRmHk+sT3YivD2rszi5mIteQ1Cf/lmL1YGoAmSfNz7JiwI275MRME5gGIOAw6wAKyGIX
8kvP9WnCZK1hHYzPFxXK3qHw2SisqcpMf4+YtXGCHDsxIdZqVULpPeta5YfiU9MYVAwwACeCSjKe
l7n0Dku/ocZlnNp83wxxYTC+lMRSJNy9EZ4O9VanlIb2iRBBcScvA3xhuArl45crElbKeFFYEczw
Aa6FSNYeaiKieWXFu+MAbeV8p8bPhtTWyLCALiGmUNqGsroBxbTte9tzRt2qXkXI88TIDRhHR/ti
3/je4Ad0rruqQdvzgbYXHySTsm9DkEM5pfxDb3S+1lrcc76mOu6zFvbADJ21Puyo/Wfj0RHzJ6IL
xhiTzEOtydmxcyB+AoNHpv1ngt8BDQTT2YnPa0DM1lZOFfR35CPadg5DcYawZrOP/1G0DrTTSS1T
Zjz7JF2HLFXMCyLjk8l5nvyjlFY4ZNipZ0F1QTCSMMh/6WSyHH3hvvbySrg+rSyjPZ0jMBBsF/Cq
u+ImAa+dSiUkhNxTYvoLwFnap2Zn+kLDAY0bwBTN7q1hy8J3ACGGqrkMbmJhpXn/FOkN2rAUFtr3
CkhkKuJt/tWlfOV8yIG38NYaWgRNK0K5tjRjGwpSAFxhkzxEokOctSC15/O5+qun1HSn6mEESoOp
yDRFQwEp0B11Y3Aj3LEyscLVZX1uENAWN6iulYe/YKKJ+kTV/6n+IcnLQEcVmRGOBPGLRjn0eBXd
iE2rYd6lUpbjPKPggjzuUpU7E6B2jBWA6QfZtJQH6JmWrs45BSlkby7nDLgrfDRksJidAXVoncSP
O3h83YV1SwUnzdz448qcY+E5UCvXR67ORKbLM19K1K2tiSwXY/TJUsM+WfxAmg7kw97aauBl+VJN
/MbxzaZYl/7oq1vwsX9NoK8Uz6M2Wt82H/PhibCzsHOIrrL1eRs40GExDWOIiZX1Sos8aPN0zFlb
0mSyNfC3WI0O027ibIyH9yRGzhu9TGQrIHwAVlfrSgfaSbRhOUPyuZb/HgeXsNtgWeZfJUAA4/R0
n81spyVNEsbfFLeTQ1B/5tafB/0XjUCRdVeK9kVEJ076AdbiNOI0yqwHcDIzwhpiTnWf4kvmiUbl
GmAFqORWuOL3VEg5Hzi8HKKMmYh8hUbuwnx3ozhe5CTfhIMglZkxNdUyjK6KbFQNSH9fhrQnojuq
mIg7IPQtrhOkB4jmF5vrfPIFoasjgFeGGwpIGEgKcx2BhlRMVakBpQDm5tnMzY1ef/FY0GLIsi7/
NpxjlCogspqQbcMJuiyXSkPmJWICOxnB+b1WpN7I7TJzWiy2xW7zmGjYY5dunrFYHGTf4aOckudy
w7IpuOhN30Xi8fz8fAX7FEKcN39kZiMgucoDVCsPqRtKqbq7VY9bRGMhi4r4o+RRuH7HOlHGBoDe
S5OVjDxnj7QNQHYRVtLecaezyEFEtVbSzIbfwG7WMPSHy410tjl5j1qqbXOOWVC8X8/eDtIW6PZG
+WqWfG43jJTBEthyItIkhVXur7n0XfhyauJ7+QXJM+k/IIXdHPaAjDVMJNjRxhS08SdbkfFUul6a
hbHD6zYxk8AYk8Wo6QKK6abdMriuh947rU8IEWMG9txLcoBZ5CHGk2Dz4KshcOQKahrdLDUj9ZTp
U99qsoyGWiUfAQo4qW8w0xUwC3MPE8XyredkOopKVYomCgh9kw8TuTX8sa9sn7CGNT2y/BM79OTX
Gl0yOekqJ01YIUCEVCyt/hPfGHMIuRkm/hOmRHDiGThiZZ1q2FV4rR5itG4DGXNPLZaNGEOH9OD2
9eQmu8W5f0g2a3KJu19e0nlODh/YuQqLm3cvVM98NUOVWpNPnbSHixctmHmZQFWG4A09Rfy7n9dJ
oOHwqmULezHwFhSsnvFEgz5xpW7CqcqSfS9NvepZlFm5S8/8Y7stDjNezGiqLjVtsaCzNM0EjJDF
9omyYa4eVwzdh2kec0n9w7o6FZYtMkyRuAnmkV6k+p421WTwaOfKYWdmwRopniqw9SZinMl9z66v
ltcFjgy1kiY3d8I9DhLUQ6nNwv+a/YXoUsjx2p0dW/ZLihxPNGfVizAkbSljh5g72gYxizjdjOMq
I4jtmcmeRKlOtGN/7+emIVwKrFxRI1AJap/317fvC0W9t8wlyNV5t0OBbHL+W39B66Zj+Pta3P47
sfYkAQBPaWIxJ7R3BlKW8ebZ6TFSLmPHY+Y6edEOZBhGkKtlLaKCIp6LHW6cGtpziil6SuDCnoF+
i+OG9x9mqR6EbJsKXi/KaUn99PGy/Wbs9rFjvWYRrUF7c82wSM1rMuwV2GWvAOJw9QtZVAavhguZ
UWnxFeI/+oOcxapnE4MlSCAp2SCxkJ2lPHn1KLjdQnd0lO9Jjs2ZoC7u3vjkrrQHsXQ9YFqLPcGS
Ol40XSkeTFGdqBxv5hi4Vc0otwHBys3aHe3qmqOKzcL3u9T62gQTHL1UYZBpXKfqm0Ddk3m006Cm
5QoXUOsgb8G6aXSMnfR5elYxU5HT870L8RHWQ2zMwl3m6aH/eDfYqSdxKKjkMGFzd92oxNWbb7vq
ArpPCZxT4SL058F7f/ku9oPgLNEaqZbZXLAnvatxicii1HUeeM+v9N4Yjc31kB/wrUS5LFJSS2d8
TFP/Oxb64J9cVFXBNWViWvv1ZbhzRO4jKPKCEkfuX1Lxs2UfqWW0NLoI37Ivvp5Y4+5SXwinE8No
rGibNBza8Z3iqn+NteMv5pFdav9/EnmNocx+J81M63I8jassmBCvsbr7xkdNQ+l5mvQD9nFrf9Xo
sF0Nxl1st0wvslG1chqZ1dp0riS4ARW1Qns+i/XLPgWzc8S0+CszNx8ZXi7eiVjWmNoKl0E5G/1v
Pl8XcFvAz1acTPdp10zOfFQo/lpVKNhA948gnm2agVH8kHLucM1pWVgXKVqlKKeaCWwHxwTECBz7
Qc3qO9K0LXOLqOoPWjwVSD1CaPT6X28hORehcoemyslUIWX4Fe5nkbLdr1Ymg0FnbiPdBYltG1Xd
Mez6nOOOfimGtj46T9J2ZAJdxGlutPfJcF7fh/xncEjLdscCrvweKRKfAHyhFRuRrYn0zzuk8RDp
4AoHP7WcC+Zu72cs1xQI6KriINjn3siKowtOCoNEGnGbHZgDrdedABhbZWujs1E/SzFPD4s/4Het
zRoOZZMWTBAzWH4gZPJ8b9oPwm4009JRPTtD+IZZfjt1p8X3LmEfi42gljHUP7n1KFBOD05ivvfe
C2vQgF+11kukH6zZe8X2pGR5fUMMYy2kOkKFfaRhC+V7ZTWvqoJCIPCwMQXq7Eal4Wb9R5eOduZI
R3Him30aDCP6Q+bqM8/tU2vkwkDDXpyWfh8qo0nZ7KKhFOP2GI5VRC/dFlXQHWGcQjiXcBOTYnFm
721Ha6kN7AuDr3in8vnFOURW6bzeyymHVjIKHPWND9JdeL5ICRW8AQV4o9XCI27OED53XG7DUTLD
4EZb12dYfCtBUhNWemCNkxj3UnalmJAUiUIaCr//D+PzNdO45+Sf0nBWoO33pDAHIxzAGc6a42qe
d3gr6J+oUVncqRi0MUqwxmXpTIEmzYhJHWqZ+rzYasp6QLe7ZkT/osMOfoT6tIQ1IL4pfvyukyaV
MJmSY365UiKhLiNvac0kZUgYo3/Yf/pBzdI611BjyumL8lFJz1iB0/KxfWNebO/orzzdMwjTa37u
fL3RQMKYgtXQfcEpCoZFWhixTwb8hWw2gam8A5nl8/h+sAWW8Lfp2PHFjYFLhdAJTZf2BM26Tz+X
BR3bb75tll9uHvYWmQtsIYiR2nDRr15K5q7Jl4Uy3gfsZpW2ZXLxb7M4isEw033+Q+ocEcSswIR0
Mu1w1IDBb8M8781Y34pXXIEW6O+/ACpgXRPsu84Bbf48xh4eSwAoLYNtfIyKogwpTSzMKarmVlny
wnGf7qV+0Ujke4De84JG6Gxtlm3g7wmx+Zfgl8BJrkAZ8MIENzTqdlHlNH7AsS219HJi13WYEoa+
18pd4VmwJ9Rvz3HypKfwpxvsC9diSnvidPVQYBueRPXipOqEnhs6NbZsEBqddb4tbUZ4OjS1mkf4
TUcy+CHgj6CmYwyDY3yzqy5flNb9mlWS+PlYoi8lHiXhF6iE1GQ4lPoe04wXBVwDhGuVYYNhRpfS
fBDvXpR/reAhQ73dZYAnpk7Cva2AZ34C4hR+qb5v1JqpKUX3HfMhmnQRZZ4DRqoHymcHNXMAi+6V
uyUzMRIQshq9fanx3TTXGM0cqMFfx/M4CYe4YkoATtCT/k/JtwCpp95zLC05iyNTob9ysj+wLQt5
N7+oqfitbWt2iUjUdNDwkR6PII7DqKaStTgRc9mQfbWSdjqWjkKKgqvXc1ofYE+Z1fKrcVa0In0u
2V2uY74zH7kf1TbZVHGCiNcI/ATnDGJRUM7wu2/B92I24+lrvZRRK8+xRkMY5F0z98NVwogrBfbe
l3l/08nJrgEaatQlipc9On1lt4djOH7EA/dqZDaiDYGxlKDDRV8MXQMBeBB3pwCdTvvEOF9j5aPr
FJMz5RAZmpzmC35So1XsctZspcQ4x9aFoc1y+aFPBNS3hWZTDonSh3+GJO7gr8wHoYyOqLv0eiNK
lTQYlJtgrFXgwf8k72Cbo4g21OiFYfaAIZQCVbgr38myAy+ffPuWuO4MYEikWsV0EvTT7y/tIIVh
agIvqanZ45NWnhdUTipjgq9jV3xnCLjfS8Nj5Vtq0yo31LUgi3sajklo1rLoZVxqaYixDgMGsfzc
bgVvAPeV8yuxKG/nSabDmMPDYxg0LQ7U9V3YlYai/STYT7oS2HBCHLrla02Gp2//WlqPI1smB69g
OZRgwPgDLYTcMMEMg4yKmmtgDPtqARSTqmwW1jXmF+MDkGJ/kCWj3JTPuNB5i/JC1fEaNBi3aXxa
wcztNHElKrf1uS3jNVGwk2WSn7o6CS6NpdKMe6OcNEornSeYKiQguOVdSE7JYIb8BGF+41PsbYRu
sIwcDbowmgXbCK0jUH8+vRh3YCeCcwTvU+BmI5g6t3awv7o9+pFmUPa1RClCYWtFyh7Qx02XZo4J
p/whbrLtLae7kikkr4Xn0gIVF11T9tZTxQn2aH2MTM1fHvsk0b/vwDHMFZQcFEHYrf3UI2Nr5hoX
IbC6qk2USu5W4V1txLsS/cFLIDxt7+BesoPxFpku2cEq5zCYfRn2kzs9ydZiRQgYBkFpzIZUSINY
NsBPBfKX48hYl4pRTT0yvbB1YH8JelZMT4soFJjzQV9cSKH/qiUQzMD6hB/kj6KB9xJ5ZyALHZox
aW28Bx3wRQBs5vS0coovFjo5iTapmkSkokvTij++AEMaRzHZlaLmL7CbjghySGVDbfu5QNNBG8/3
CvQ/6BJYbGhnsZbasK8CoJQEUC+hFGxDLGtYKSYR5HuC25kwGpQF9amdqMHmvvjO47vsa+XuS20+
yMJpAJ6c9f9J9Gr/lnGSzmVp720BWeGaTilW+giTlXEb5mwZ2X+VRypB4/Ax887oAair29jJ1YIL
i7XJS3OrgPLMOvc4Ir1qfbaTb5HWAk5FLiV+AEy2hrOVHVjI3iDvgOTWEDYFQbtWywA+bc+VF4tU
uO8JU2lvrtEKrpvPhympbfMF+Y31B/M9RNA7TOLYhcV2TmlbVhFgXQ/1DGlNVLWT6H0Osd88KkUx
uhzmw8DHHpwy86IdpdxcIEo4rUV38F+GxfC+8JSMvZuyFu2H1Z0nl+O/IRAfdJTcyP3hGzg5eLeF
c8LqdmOC3lgT6IUJahe1xz9aD0I3IPbSNMidNx+Egfjl7DYSO/TJLqNmnYi+a64b/f+fn/QujeNy
NKra8uda114plGr1V+beceO6xmz71Ic0MaxbmyEmpTiAqCSexSp6k/tCUuLuZDmOfcUB+l+rFPz7
5fu24DDb89O6FvIX/7N1UNaqFRebDl5XH3ePUb/9GOcZtPg2cIK4opXK47wUKd3hGGmVQKButscd
ZNlHwvAB6o/Gj/PgLbW0R4mSzQE+MtBRru6+EqXs0WjNUhsyQSGmEbzUit6dzgviS5iJczKhZ46H
Fmsx+gV3VGOyaGzvN9yzMu9e5s4RqflTWscXsUJqr/2v7eU2CUWMv9GmlIrMXXv1pTN/ONiUSVbt
cqxym1Nsp1wjIUQ/ffG/nQS7qtg3EFxT5u7Up4tC6zDsGDQFUysxfp04x3n86Mn3Xo2zt+DQPzO2
Pq8bpfjgnNQ2wGX5eFvx/UY/ZKDcYlRVovfBLAdYzw8VZsw7kaB2Djxoy4yUUcjQi2KR1BOsTCRK
B29Ixw7ZLyR7HDSvBe9V0GVMuy3MoJI7jWBhLqIE7Hc+usLQ1cn1qs0KFztj6dzWHbI0oDIalhZt
V6ie3lH0a2W3lfDRNCw44oqNfxLYQz5n/OzbBEdrTI7KW2wwP1dFtaaEGsi6+XJzdBsoQU4MPOT/
GFS/pt4iQh+pjgu9TnXd/ymcr6xR0bTtkOtPJEU5zQHFhOPnV/FUiIbFkdccB5/bCi3E4p6W34Wk
jhEDoVABTKzh9165xtLzZz/SQ4ucfD21SGdb3w1v2So6mylIuOfiovKZIuF8R0txVlgbWKm3D0Rs
joxTltHUjXayppzx07NsZYLPCIpLiF49HqWxa2GdPSGErdLOnIrrt063t/TbxEDMohUnhFusoo7r
Dmbj8eE6qhxcgHiFYxfyBWKLWa7kKEDOjwy2Picc0G2h/8MjA0iA9+xDYaJfx++FQ/zU+e9pOr45
AK5BYF4q3n5IQuHxhzi5H9x2yuKFgEkjQoai1lzlYs4K/8ZICPZD4nWpSEnNKX2j3r7cdBTUBzKY
ohdLrHD5n23Ap0/CgtjuT0x0azL8WUpyT1XIKgfLD802QQsTtvNdQ9kRqrvMUU6CMoTqjWKLD+6R
Bn3nfmgky5Qopq2xkg4rv/Gb+bAZsOiabcmaV9OBPqz8monvNaiUuhWnYyfRN3dHQlTFCFm3PwSs
gqMR+mg/0FyRC6Cvo2KVqq60llZ8qiFvS1rtGamWSlnBCsKWqeyznE0fUjvXruzWOSIBiDfFfmy8
xJpHZ/w8cCGWoYYcptM0d73ntMDed+bE7DsqODsNPmfn9A8pnyCAx6gjtWKXDEYgiupn+/zFl1Zj
x1N+a5KqiX3sVS1Lh4+TkaOgul5Q0tyJpDIuNtVu4/EQxEvgNz3Hv8t5/yLKGS8h73ByNjmbB+yC
wXyIp8N+vOPYtByZhp3e7te3NtdIac1pVRSHafygKn6LsD95pNdXSN0pUO2mcUIk8Z6Bp/44CwAa
ydjermBnE+LWHQcrkGsgmkgY/igUiPzunSwzbMrNYbtnQGDERwJIKRDEqYQ/2yliwVYUDO67mIz9
OtnzNOFQ8mHfTpEGZDUWy6BWpUkBilpAoMDMM6T3/Sh2pnIY5/8NX2XBk/er88tFvallrBnW9OGw
lM/ZNIHgAzm/+AkPG24y0mTrrC7UY3oH24F+WMiGBeCpfQpG15ozhTlNXbw4ICdJ8rrHgVD/6SFZ
TvK4k6ogej2Ed53lPxDm2D/4zo4MkRePeWA3rM9WktbVoMCHZKUB2PU+g4nNNRmSpcDwiQKSs/E5
FqYeLBtoH6EDN+0GlMCt9xZS4sUECaTQipQHPX7Ow3TDALWYUX04xlUes3QHBgft6Z1Z4VOdqyEW
Xa/BtaXqxF1jmzGteoJrfxLk7OSksh2r+noMfgsAiGjynlMmcloLGTbzGB1rOItWqrBxJYj/u0qr
GL0BwBl4AnedcoqufSqhxbuVYan5CEYCQmJt9XdSbWWrlnb6qA5Y16hF4vFaVtvgOt9USvrnOPTq
9CfbAqSZiibYFdKExPz/3aDNe+8v9Qn13zKFrKIvhoz+BH3VlMfnl+aIPnvqdTgqsaTGkmgKYnu+
mL6aDQTRYJ3S9LWtl8YBus+KqD+zPqkxRyzUVdAc4dLghawnLXar8+GrXrNl7fATtERtCJ6UMzf/
t0npTmADVUPx4UUqbKjs2Xd4PFOlhe01S6vt7YSNwc5Du3jfTcKSG55MeLizyK9CghRkLnBa2WgT
U8VDMyJJLnVUwGY3o15ePJGHMGMAy8PdTYWDLIM0Acpw265uqT6N155K2IyqxuRhHbhJQtZKBIUU
5iSgyRF5U4eGTNZRA4SaU5Xbw5rwbBdaGe2NLQV0+sx2JM1Ko6T2ebd3OZWY2NTAz95CPCIvAMwa
JCHMsBpNQTxY9bMQ+mTHBpHsIkliyn+jbRLnXeUwSXzU5dOPjUbVlntf3aB6dsQQpVcryA+8UB0A
Ea4F3IVyqFFAw9RywSq7v+3e60mQ8LCh/CT7Zk9O3LPn2ekp5IrUpha0vbw15bBRzQg+jDaFvKeI
GK1ddOI9ZV845qK6cwxDnDbI/f0RcCo3dHJhtZU495svouoD3SXjzNMUgYnNQX6PuG/NdQx4B+Nm
CUZvAUiYtD5G4Sx0u35SLrXwCo19kngeZPM08hBQDRZQlWkayC5wWfp68hAQTLDGQFGC8XUPZZPh
bgaJFKuYv2sD5qvgyPFpgrS3cHdws4cb/V2XxKjUfO7TdcpklhCKwqvsq68cjy3nlSH691BzVpkh
B56o+Knjz85bAF65+mgLNBwD+8Iq6tMPPma9PPTBr0nU1ydqfaUJ9kgjl4+OZ1oLg/WdzB1gHCxQ
rJ4DHW5jHarIGboiR/kf6v2RQw3D9HZeVYyqGVYfcGNVI25LtzXl+b9SwcXrWlWm9EbZxsP2DKBo
YlKdWg9+c8S+RfcR5yxGFsnUDD37YJW5Vhex7xE/4TZgcQ6f5/CQ02+AU1f4w26cGtxViuourpjy
9YuYYgtiiOrL+XppU+1TwB1R5q8CsfMflOdRXaWwTF43N47QJJjZIKwibCz6CN1LtnrdRqkPfCAY
6XnGw/eAxvAf2Iyj7XpKtWmgf4EdpHBDuy0wg3ezCENDbRsFoaZZgsQLHPzhvFa3ptV3qkZeFEpF
7F2VjOhCUYDxPF5d0WSOEvRmL1M1i/wPm3JxoVed36bI2g/jO+HyEeuDVpn6/VDJoxAtuog2XEEd
ldTdSV5cAHHUwVnWxH//UpnYA0IkOHyOROi1vxwZKzIEW2TwtZFCm3BV7twx+RtPv6tZOhERpcmT
69WQGxNYSRfr+J4qP25AU/4eDbB/aQ1MLzxK9EdV/x5YQQX0wtCZCJIoMFAUr86ch+rKo4HMuW8L
2BHwFAzui3xFPxlVuanBBOeLBTgt49zuN7/ph/5D0/8csH1d+1cP5DY8WpXiFooDesScCihAEM2d
lU6xDufXgO2H3gw/JKFwWnp/u0oRSdgo7i9jfHAyP/NWs2ySgEK5+9xKrdj74LqaykOOKR94NaFG
QIVDXEt/2pCI2t4DAIWo45eoYNV/o56IO8xTvMfEbKqLHb6NrdY4hBy5UQov+I5+POzViPQo77oG
Iv+NE2JpZMsys7VkQYIkc4VcuRySQbcsg5wF6HeTecbuZv9IjMPYB9Jr+EB4yfHO33da0rLBacNY
lRqNTH+sX6PGyOmVlIXP7wLexeen7EzCS0Qme17c9aEdPkYMqRzjX5x9xqxAkaVvzfrHnBbK+8Zg
Ui5F/xAapiGSKPhf4v4pPUcgc2Zmwhcf0DRzEyb08VNyA9uHiLCuXDbzglEQZ/XPAoMMDqBTaxLv
4wdLMuKkON+zqtxQRosXV/9UUn9gzjYZoDBC8IYntZYg4yJrXLssJqW7in/ajtK1TcCXNUMWlHrq
zLK4AdnHKO5UgAHK8cHxp+thX7Zo8WblYBHOD767RLt7wsy0xb3UWkIyEXYDhiAcTx1MwF8HFnoX
PVUsLeldVTeiCzHjrwG/19yTck/c6cHjtVv6jn5hZfa8ZsdGB7OicyyXjRyritCPXuLe4+PMmH3h
gdRyoWAeZns2pFhXpzt7dyXIGzyXCUJJJEQ8qQqA7FWZcZdLWjHhUL7is//p4g4/WKmxWfVFxioG
xmr34a7yqAN+qZ2xWbYoZSmuanJfMMXveqwPhZ2wh3Ua2YnECVDklMjA1S6Upo9u4+c1Qb/htSke
ig3lizvAAvZE0SJ9Ev2o29Qrq0Nj+itQPt99/P5edM29TAo3/aQxD5Y2m4LQimcrwP7L638XqqmC
YaGH89LA8eeyUNI6xjQckK34qbpg4qhkYGNeBIzJ3pJlAT6xncvNbbhHtQmA1wM5KxujTkhzrHHP
LxTCpTa3TzmEY7KHMSxXGKh1iO83EFKC+pwM6I777NhSUvYHLPSbBbFRRnyLLJfGrW05LC3sgYpy
NUcE+noYy9YwIQTMkoUrIIimt4TJrJjCqG6GyVe+065UnZ7Tb52hvNLIVLLF3ETJwMUdaq7XSRCs
yDSO0RqEcdiH4/SOLnIvP/tacBnqPgclZB+qMn3X+AEhQ2k4G4TP9qZBTBoeTbxLcdCUf/FpuOOk
FHuILvRpC4UGDN+g1BRfKDisZtGNzkz/UGIUAZS+vImrdU2JYTZZVHRsMxzRlASdo2vMKTb9ePii
SbBzQZ+6bSrJ3nHDlgdPQyAxa34Cr/Jb1Zxbj9tfHCmW+6W9S5eiA2dZLyik2L6mJQJiAZuwvWA/
0lfvhohIcwRDqAD+e2hPA4FRasvBNZPRZdGHrEhFUjObndTL1cYdh58R2aN1OPPbBoKmoYKkhzGR
X8zfYDmWYfl5Hi527ZEjJZKAWhmCWFEBU/Og328gVhMyUfpJML3Ah57D95ryjJHT0Yw4o8FMPSc/
6dSPadPFHZHJoh5/hhGVI83JvqEhonkmHdMt4/KHbYIJYBDbPqjpmG/WCEXIm4FlcVieEz4Civb+
WM/uSadoQv/qu7qmT8ZMAGqUbDsGtPiCUTxqq+BVcj71Amub1zlysD11JKdRlK/3xmz+2b76Gwed
T1KA2K6X6EX4ORkfNORLHI0qUvoPQ/GdeBaEYO9xxawn9Tb1VZdkh+xLou5BVcQ17au7KV2HlbpE
YQi9X7JMzwZ5ZQ5tZodgmQ/ogEGSdF0xl5q5JzgilRgyxRn6bLiyxbJGYi/JBt8pWxMnSdXR+3Lr
HdoCtY+Peic2eeLOxOGx/TDiyqSxfoxMOaFkf6ZW015v32N33ikvQpf77Z4gW8za4hgJbXa/1tLD
IBZQY3bWVr+mXyWAnC553TdIf/c50X1SZWKUwGbAz3uKPGRNsLkYezsmfpXoWLzpk0mWbnj/Fgq2
HTBzV5Xwmmka5O3DqN77ZigQoX+DIKp91NCvREd5IbOVvxiHA0WrBo14e8e3Nn8qBD0QSiN81bin
6Z4lqRxKiv9lZefZ8amPp2I7lP6/rAk3L5IQ8bmEXSkugsm+P0qIJgv2jQtSM3kBx+cSqY5LizEF
zq7gers7Mq/eP+OmwAebi+CdSO2nh5t+KKst5crI1UNByqAUoiVsEdYDJA7vNIU15n+Idalho4o1
RTu9VGSp0BLLjnnc/NWSLvdyRgNyKhLdjZTrZ4XcDmChW5itxpOKbMsy7jNR9Sk6CrE407w/gVoD
fPUp1AlXqIPfayeLSTLimL6rH1QWZvYMK51d+jvhcFXMKzdR5tQ/bRbv39rU5PCsU4o5B3NAgS1L
JSRLSTI0oCk+KyiUyuA6UBu/wvbIaOpgKl/BqOPGsONmKFdAg5k1ejI7oi/tJhVsiIQjITbUn1/g
uSKnZrvRXHTwQMGRr1mtRGEdZUTWg8SUoOgDNSz/g1dJfXUcJ7p7H8A4I2lQk2N3AdwBeZNdPOE1
WPajLDK2cuystLzqWHvMtEUD2pJGNVNYH+cVFuNz118Uiicw5nAh9GVHMRu3h7AvQcpAZRTwA2xK
G+DEPOwQAOZ0VgiRKbvVKzGEykAsve22hWi2Mot/5mzW5tn94vPphRarqjqLbFs3CeTyfH36XLw7
ybe3QmHZbMbNFKjDRwUyhdrIIv9Wrb+Ve3TZFiWX8nEBWfJDIePN0BA1I6u/X7LCl0e8UafmWMpU
BpO5Wii667ROdRLsC/mJ0AcMNY2UCbKMh5bTKKaTNr8s8Q3HetcZB7+nWBwsKUPF9lfZaz8lGUZI
84kr4eVlFMxTMVyd4Nxq8EVtkx6oj/JYufyxjEniuC0gYlfLKqOVg3+kP9YrT/IxsjoCyRjkZdBk
VpgrpmlsBy0aBm2ZchYgPYJZtQhcv8WNRKk+FgbjCy2RqCmv22etOjmJzbH3kR4SUrVRQb2oL+gx
PeE240pjZ3nYSxCl4WbalrJ4ekjVOpQr0YsRlp5981+CLqw4hJ1K1FUcIi7mif0pkHgtPnkzCB/K
SYBvKobGoMtjCVpoWrGKIFXPD75scVfHsoeyvBD9QoVddprA32DdhPb2BkkG54fMfKkDczsBC7CS
CGZ2ycdSxpOOvg5a7uoI3C7huAjWRcXQvgtA6H8iOSYkcKoIBsUQtFU5QcbNKAfcofun+SI3OUCI
C9QAgr1DObDSalJRy3IJe1e4ap9H9oHrkk5a8L33N0Ghwq7WemnMjcSA5I7ayeGui9kNXcQcd71v
VDj6M+5Ln3IPqkL5CAMukSSDJTsg5pCVmZ81FfFgi+ND5Msc6oRt228e/43x0XVs5mU5WF96VzG8
NE0kG9oyTMe2uKwGkBmslBksKMJdP14uKeffBushjfz8+ONJyv6JQx+WWR/rIZ1XfDTv9c+WDKCB
JAbU4fW9TZVLpJjZYSrglPbaGnn0PvaXgLyMkwXLt2f95o8NTHl0+Mb3SU2N6iDU87n2RChyYDYS
/FqT6rKwZYQa6efQ8OBo9BYmMe27g1E7T9EOT6OGMr5+w5Dr6tE8q6hg6u3ckbhGwHPJ9lAX0HX+
OKERGIJpnzvC1twpASIg3PxuDqZ1maK2f9uK2ftV35yBRkOcZZQ7edvVs1Cn7F4gyh+MoFdymyyi
RcVl5EUjNfNsB9rwXJPAnlC+LQacSrma02n4vxuL8Zji15q1fBqhZMS2I9O1uW0a1mBp/Hu7esQP
QulSNqvYqoJaNRU6EpR0InxtS1byE4AVbGyS18HyuSn+32aRLE2bZawAcvN2Kv+8TFG3t9gU5U3C
3wkdvnUxt7GUpDUoyT2FCEfY/FO3ZYX6FxJlHme2a7tV7GaAwPZ9m1smDE6/e3uuxOeoKSBarJSl
x1OAcmdPE9Wj5bP8cFjblPROUXYjL6Z+ImgArkTUjjMHhFtR3XB0hQqMqB65v+XLVnuf+7hXfz9r
U54x8BboKYMC6HKXENLI43Uj5U8XBiq7+Kl5JtSpyGV4ZX5p0EVaUgmmIFD/t2XLQyZ1/p8W6lIt
EdGvhxwqXPvFZ4EJAQjcjyuYakqpt/QrgK/miAelsQRhgjroSo0P/Iqq9p3SXvPlN4sYikerfqHG
EP4ctQf1YI+XOwrzkMobJZMF8GEddDXQDHUlMa1YwHBQ7deRQRjBGoawG8OyCQ5mVWSEip2vTnzY
pgiS0V1r2fzbj8JKnXtQCP1GqPn+H2Uscgxq1WG7GVgxzp9nvrOHHDpD+CokJzAXEmyXAYtvrzTf
S5qbtJL/JAl1XpsSVsZp7HfxEXTlnqDjVUyBEnXIvOqNn91zpgrcGX6v6YIqR5wCNApAUnkhBclI
rj3v19ukA8s4bGB6er450ZO0T6Dcik9bsHhxwSS28c+0JjAlJyOL2tn3LaqlG9WmX+bf2yv1X0D5
waBjFg8ZyDq7LQFCtj3HOh5pkw5xYOe5SVZHK/qTmOZnvyuzESU8jFiLyZKv93hbDpjinGbJyEtR
/IHGcRaeuhVTNuasEd9ZMAFN+93J6qh2rtnTqb/Ex0mLuQxTZeo5G3NReu8kaSv1EPddRDZuZd4x
fHZDc5Vjanc5gm7UuPdTC2e2mq1+466MW3lH7tPUcxQmwCJyVu0eAxQJNrUhj3WZ6O5affEXDdnC
fYE+mqY1xtqNwwkVtNVl6EPRderTTKvMbA8i4ke4GhAAtxcljhYaY9acqiJwV0c2CqFxaNiqtglr
BL8r4u0GDuIQ8WlqhUVHvGBUlnWEGWIPfL5IRsWVifNiM31/6uDU8g0t32Xy/y3rd5vpEN5zJkZK
xPRL+ljrTijo4sqKT2fLtKJmwk0wH0ahgQdS3+UvP/VMu05ju8loYcfZy4wKNVyNKEYCk2LE/0ga
N6qeadOvohiX8oDEeSS+GQyQyguNPDhBz2KDs6iZ7YW7WtnByDOY7FvzwyOpdHqi2x76y1fpCzJi
QRILUu7OGpk7JmOQm8tGBH28MxFQjbpkQIDU0lD8hfcXkslWq6HINYg1KGwWmLPLw2pQj8Wne1T0
pq/Kp+a/4bYECIOykuOPOpCpapXoIErYSHlnf5QTtQMTWgI/kw9zEHne0WR+ME5Fm65d9O94ysVd
eDa4o43f+cVRrobTIwN3xINv0aExSte0epckMRBzxnf/C/Tjkq+5oeUE7NYhoHjm5hp7cizqxqaS
iW/D5lA+g3E99SlVV1xZBJUHeVSiiXCzrksigMjmG3dNbT2/U+kcFBIYxoWIl5lWb74XFLUPPuVb
UGH70oYhQZ0AfpY5glF3t6FkcKO6iIUScJlAqbwXe0Z7cDTWxlcuwyKQGOf48WdLIncgjQSDrgkH
5GC13Vdf//4ItqJOv02ydRDiO4JaTcK75op9Txb3wKPIMsyzrs7FwgdppMzTOQGx8/zmeF+YXF/U
21+dB5JRD8PBD9+z5ZkP+b8SMG6f7jX6s3cs9r8qZlqYD4FOcwNzkXvx2R6wsk3dgDWYIymQQz69
R0MijBlzNIKME68baACEXhHhoCUGjuynvSx15ArxBq8Ow3hch2AHzEMx0cQhoL0VrqCEmIvQZN9R
vceo3okjn8ODZveztnOtWFrgkW5H4nRwqc6bY4oXJCbD+EVs/nTeGy1Y05fRtP+1WPgDs2szkRDe
QHrnGGSlEmkHD2PT+7MHug3vaeiQT13WQlGDN8IqUfDePtUeyXR9VtisO96OG/7Ps9luOdDcngZN
s9yhHR//0iYWeCykyZ9pzJT07nD5/qETe95/ILeROBJrSFl630jAX+89Di5IcgYPGpqvChFPJYil
VoZoqNmKvMcTPNqOgtoZSpJHitRqqZnAQIQGGRtrVkXm/ASWblGmG9qg2uVT752QXNM5fePcSQV6
CR2cgSCiNFWe/JzHzEXfyRo1PgUny8l8a1TXbfIorB9iqBVXFbmstGYAg5VX6V2satSAHbl4Ds7y
CpFEzTvmu18s4itcC996gIAExv7BHTopTtE4mQpKwEIZ++meywI18OzmW31CJoG221/B7SjeBlQ+
IhrErx3wkwtmWhMvor7/XcowWXKV0yhmmeln/GcMNbJFKZjtv97THvITdkxR33Xxxfgr6s9UqbEX
LUVVYRNr3UEYJ9WQ5d2j56Ug12YXHGOIC9mA+J8KeSFHexPEDsuVN3zhS+Xqqe8no6uHRoZH6XZf
MdybyO6FKrkro326kgKEXkef39ruU5QE+AoLPVdTAs4O2BFI/cA32SgFD0aBANcizotqpqz6WHjU
e328Z+L24ZkbGbpyLiMS8/KJK4fwaxuYiVfMNyaydNdo5ln5kUWTqv5niru49clSKJdJKcEcO6+b
PiayttM7BqENN7VAUVpX+aiJIaMfbzRZbxyBEcL0qDcYetKe/s4IFexJ0ebmggf9UkbLsyxjFV89
qOhMSrWedybx7bfR6FkjcY6uEql4IMY1nrlMGKmyOur57cANcNyGiCF6e5zLmprCHYJ5UOWnfTgu
+Y+WnDpRFCq/4249OhoquOHN87rZuZ+57rjzp2A4l7YfsNuOwSem3pvCcYyVL+JiAm1xLD5aVJrA
a4p8UiyI+LpDULA7VztK+yai6vguQubgyaBx4f7Mn9ILre1jhANBvGguDkPVjGIWrZrct2SsE8Bs
LnMnci4nMAsGUSYLdV15h7sY4FI0U4XVUsSbVOHr/KZatIEUPBGUC9uJ/oy0IMqPGUBHuegEZtIk
L0S1UgD0RIB2KseAAK3npShKCsxSC72yaicPGqVzAqMZhBaAb0DHxFareU+OXRMWeAn/YZRWZWNW
wM4WQ/RQiriELziZRPBEl7HfU90dpRQcTPNHfHDVZgiWNqAMQc17608CBDLZq3YzLRzLKL23d9mk
V+Qvm4tHxGjPW9CQ6rjoFw25smO82C8dtYZ4EI7w9KNzVVFT/f0ronizt4i/YYG8uJe/JdQ5lYP0
on38omVdwJwChSIVp7H/eagXzGQFtRMvAXk5qgeN1IM1RxUJ1+I35d2twqAhm1hbmzvzEySffgcx
c+HzG2uPZKtxieyupzXlRJdyYSiONZJFHaeD+pm415uGAP5W8tx7e0khCol3ipO7AEzQBgRMnXLw
Hy6PE0kIqJ+BQ2OTfyQ9yHxYfCZc+NJ9bJtm8HQhAONqHpz4IlCb5cDjWrnZfmohf6O+gAus2tQj
kHmJ4s0VOUXiXPNQKa//93KaLhZXnup0llF/XnGPehBa/7YlR9U7myRucPvumXpEzCYeiM4AIW2k
SIcN8qXdxd2dc2/O1j+D4yB9ifZUjBb7DmoZiwpuPrExAQLb3FIr3SQfb51Rs9269FU3nl5lz1Om
b7OBuD7Gs2uvARtzj0MeBKsltIH8LPhAIeSjD0ncakN3UYNY2sm/aPhF9AITswQCwoIj8MDzIjZ5
mWm4DQ4SZ28rSm5jhwrLMTk5CiiO9WV2ZQrqk8e76KedT85AYXuqjCQcZ5xPAFy3oCnRjw5dwKe3
EzNjxkuvVEVUgn3t3TDAepSpA+VolxlkxDova0Q68RjvRdcTpG0k9Rn+2C8llUi33HwA81g45mDH
XmAgXMOJ70LdOqV1rgYlGy9cKXNliDlSBpdadfIUwZ3UPEXOwYDP7E+DNvlc8k5p00+GFPmIxD2I
daaToZJNhRAub/UaG/fmGyzj7xfeq3F5xDPOSPqxrrGtWdVQmlryfpXswIdVl4PKIaapdnS7COsq
gtgE07tDQp9kyjkVAKocJDMK3tZg5DgSVrmM2vU9nugjSQVX+PV5FdfZGrhOvKHqSKTCtUaHcxV7
3+zg3MVq9gd04lan9RK43Lj1DUFNOKE/qLcohp62C7xdxCo6Up8UD2vomQyE13r+xZYuzvTpEkpe
OJIy/xGuEpZ/90FJx2onQGQghKu2CewnDB7so9IDjtXP6bIemukqLA0yMG4HLFlLimYIAcTduk2n
iJ5jI/o/S2DS+1G5kjJmQe90/1qwJwiwmGMyN2+MyAPcBr+4zQG7MbtI/p9e8nV1s6yK4O8bsHX5
KQXFOW8jAxnCjwPiGlVEP/N/tZMRRbB2YMtOrbOvgx+Dy64L6uqHmr6QQSJTMXJ28hjly5Nd2WZa
cp9evrvFeEK8cG+XLs/1HSdyYRCfSURacsneMFHDxA+FG7+FprALEKbt2wKki1WR2ETV+/2sCuLj
hTydjVIlzL7iery6ja2bccraJ3hMrK9yTRevvuWG0AKPR1MrCD2PP+8hlLPOdFfpQflo79BGQAVV
NMydMOxp6J51Zyguc0Pm071NfLcFr2BxhvqYMYdFCYnMslKFBGn2xQaJ1cc4WnS0Vq1/3qRKmYk/
540he86Xj9i8wBNpZnFR4ssUKasFsRHvfDa9b81xsu6lU+2EKW4XJCXvVof/0FsI79dszZAWzrYP
x2edUSROjZ/0FyYRKXPuMSX+PL9W8a6pSGSLb1T/exH9KlKGYSiQMcAs3+WDzzBEEqX1gqLlacpi
NQ8djSxal7hzk2IJKPnV5td3M2/qYe4q3JetO5IgV4Va0cFW8/A/buvx5AzaQWZSW6gAAk4HH6WH
bCA/Y3DrIk4ywkiDl1S4iUjDs4EeiNwgwCJOzpPONcKpQWyxwfyMa7yPjyYxpiqTJM/siXuvpRQz
cLyO1D78PCjhnWFRcKRShdRoVKs0ICKK2vl0VNjejQU3DNMnOR2TnmdqOfjj4L4OFK3SrtvCxMMZ
J8ta1dVXddhEzQudtTrzIKXmowfmYvyxpZX8iyj5CcfbMAcTP24F0uB/cQU5BTPzqLQcA+T9eQfT
apyW3K+RTTBazSlo6SNQL32hgjS7iAY/d800LLjnp7X0dfCBF4vcxjDaoH1lKMDG5S/xP0zHWx9O
nOr/mK1BRx/5w6CHur1e4bAMrqi/yFGov/CFkuPnhoA7ba5wFV9hebG47vaZ4aUVTdi7S15jQ/+p
h4BiOs9dQWeU72O2zjpuhv++TWhVbUwA2hVr04AzkXOHpTW59Uhs/TsREy3a2GifJbXtSpCG7J5T
b8uK3QI2OQWQ3nceTs34qI6sBivwzo4fismygLO9piDoRxUGD5HerjmV8MI50UYBtCmBJv2Yo86b
AVhHwRR45iE6dHxJ2pVkcekH/PbPqZxCDWoYeXQjzy/FeqlJ5BXCYqLHAHOFYXQG85kqY0L/0obQ
wE9jc5EOxwpY6hfJmcYlqeq/OtFZI+x9c4mOILX+9sRlBLICAU98v288Cr+inNPizS4nHqkThgnP
7YI7SnoNaLHZskc3hhYJ6V5LlegKuHu37bHwGujYD6NiHbx6t5ZZlUzLG40y2EwWqeMhiRTtcdQ0
YF5uGFGS/TGAYkyKosJFR9EAFKVX0h25vRw+7QXkjkHUu2MabA1lpTc30OC/RJdcPMuzhKzVFxPt
qPXKUXaTXeaaAu6hscDazp0l0PNsfv92aDVQzrY6qFG9n1vpor2SBIdoM5COi/2ETfOxX64e/y6G
EdHjYZyGytlGGnQSEwLk6wBH8vkPCj4+VmP/xGjcpI5bW+zA8UkBnInRjLfM45YfIL6vooTVrh7N
V+4+wMPd76Px8QNGVQscczrSRl14gcwf5/6+XaeeqMYkl2Ly2+p11Kbf2q0nD8GR0kFyryztvXVV
zNeOize4OGFtWWPW38VprlrYSITTS3PNT7NUhl5nZ+/nJ8zo6lEZInLWzCHppiLRrU6EhjWkgflx
fhm1tLPbQ/ppa8FTg1XsrioJBud9ErEVe+zyn0qpFRQWvBSU4a+zfplYI5comdL/e4eE1rNC+ozC
qy1qBmz/DlapBGlaQU5D1FZtk/Pb4cl1aMAWFCKpHIYn2egTdj6yihkd0r9Y+2BigIQJ/Ego7qE/
9RJFGa2rRtqruRffTMRnkmxd4AW4Qf43SPu1iROB6h68yj1dSl0GyRf7Ik24+W3/z+VHNpGbjyfA
k5JYip2xb3M44t2uyg3hGD/Db4g6FXdMTkTbxN7HjAXBoTDImHfmm/rV7w3xuyATnPy5FSHI9duV
cOldNZ7uEKDMYZshVNfl9YVLASLYsbOUnh4KHo2HxPOMHBxJfhqz6GA1x5sOB1Pjia19FyHCvZMF
DDyWRdm5RBQYbeSaDFpE2dk9YwzBddOoI71rAPVVsDU4nWjWJoZ9v9u61Y33Gka0ZH6oTx3oj30/
SlBhWMOGFtcDMD0/tS7mzQgLu8NXS8qjd+n+F7p17T+QlVk8QzW/WOvh96gc9294j3HIFsBnQEVc
SJDfRdRdKwHAjAhVC+bWfgfskfAhWs5TQOnKe47Ga04iKp/b5i1sTIDmIrac3Rv5hoSjaRbNI01R
/4V5S/+vRQHAJj27YpXDIogpKlyF9ulULb7KJceqI7RS3TUbTjkkDC9MJy/nwIVlhOgKRsMc4Hdj
1WQdj2yVml6hnfi1nd4r/KEFRaUJFo4Ebt/VD5sXPmBH08HfWTGzJBZ9GrdQ0po1RyhXaoHsZh0x
lCWM3W9Jzr983OcFSu5mt+sQbUkTKDhvha95Pl0EVGeZJ97FfupUkcOLjpDnt8RIy8YXU8WOE+JJ
ROEgNh8bJRcpt+kxAE0gUph/dlwHl+Tm2jHSLl4GPjMt7+/VXPLFKMw7Ssm0xezDHo1AMont15vQ
UvwkGZkZrdwIInJu78Iuupcl2r/3/7UtIawZ3np0HEZzaBNOREq1rKvALV/l+jL5VZDnW/boeJM3
Wyd7iOe9P6AsCzYi7qLjyMhDCc8yAKZdYNIyPr8lWVTPiAyJDewAtI/YKgLK9fEIXg5aGmn04J1b
cx+SQ9JNCtlfG5/OmvD+r0jfMYbR1iCjqIVq8g9p5stFkBkpKaTHDsF//DryXJBZWMsAQsn8Bxi8
YunqmhaHRMwSUQXq28QeGUBxwDrLUkFREEU6B/c0pS55XuwJOgnuQsbik4LQz2HwYz9IJ0nNs41R
mPsJ94HV0i1YbLJOVwEESIBwwVoMTxSOe4aX7wjzzNDIUk6ZQoXA1E3cVQ/JYOnFIbH3A2ZMTLEw
AhTO2goeiQ8d082wIqtsojvSZv3/dU3ossJPf1lqxxnGTJhhb++xAgruoxFHk9rulXbANWageQz9
BlSfpXdUf+grFauAHsMVQQrJATI7n++1cU1Z3jySL6A/5DUQ/L+siOPy2jlTVN/odPwkl6MehFkz
oimPNdKFVF0ow6qmEKDzqq1bUu8JLimuEOfR3WP5A6YJNbzwiJPON/SQPyD6rmaIP7fbX8+JQrgf
PyHL5CSkhYxyq8vBrZ5j52vrm+6JJMf+n0qjVz/z+ILi701Ncm8pLIljkM+aD+rBgg52kIXGVvX8
/Ehk34Go00g/uVJDj83OlVMV2Nl5s7Ww2OZ9pUn+cUU9T0Mjkj/tTSJ5NZDBLCvhLtc5eDjrtJGz
UvR5YRv4MPPZgVF17TUeW0UfCi4HRB6orm7r8WaVAALAfT6I1HPOrptJlTZJUZNQa+y49plvJ5I4
HYgpvF112r22QMVJ1v/RgoumTBiZxlRl8biRB6Lm7bquVfSouLudA58Ds0kYGUrFUaH8AvnmQhRK
oy3CtI4MMkI5JCAW+lvc1votasaXyZkQnsgMsEfN4wkbWAOiz3cbvpXYNUyEfrK+ezNE+GmLJB0i
skFiCv+1NjHGanxb3DwVPTfIFkOe4a+iRhdS5j/mecijsrHzoD5G/vpznqjpAG4hPewLXcK+5ZY7
NXU0evltqKQzLXIrENT/x5GBUbRD9QXh1UIxSAy+VhP+4uI/zAWX7OTFSurkdOClNIhFmEzpRj2P
Qb3E3Q5R7WnzreMcdO4cIbs9vxRuO/Z1q5gJ5e4qePwO9r5PaxpSD3OCBtRywzC2iYgq4M5PBaWK
NlVy2pnV0PRFnbSxXJndwFLypnHHYwSYXGdalrh/k/QK6AQ/khlFVqL4nNVUFRp3I4MhLMIRh2CO
hXZfmRZ9bJYTm6AosN3h4YaBY+mp0yja+Y5wRkowpGJJGoGVBqCRwg87qK1htpqu9y2+ap4nHC2i
uevQE9CLJs+5OjUcwiV4GZz1qu3gyMQztLcf8Aqz46i+cTn4Br/a1fDM9fkALrBLkB5S31m2RDCa
yWUu7QYX25JewaoqsdHs1zAIPjSa1yHHKiQIBsRgBg/I6APWt9QWV+1HIGh5MKs7Xn5TcOGdzlNZ
79IXDm8BgURa/tRcMDg2IlO9Z9yHoz0u3UUwAZN++5dfth2mUYpoTOAXj7fpxUILAF1Vj57TK25f
S3zmy42/xCGoeF6hfiXdQzUwc785f+T1qmk3Xo5x8cIB0KVZ/w99vUJNBG+67pZgBrtJBiXBJlnf
fRyim9TMVM1djiu/ytzQoz7gPt/MHs9XODFbQogq0GXo2WLjfeRXh2D69ywUmJZH8d+1LPJKILEU
7+UvwF6f4Izwrmlgn/llfmHRLWdYIA8m7Vh9kvcmYheRMYeAsS0cWHnRQ89QVXWWbfRXnKxmb8q8
USwjKE1ZlCvetkbHIHkhvOCzVADtCIbspkt3aA9vFDWq3gWfW0bJzs7zvRcFN3V+0PLqdrc35dru
iZdl2VhwONcsuKaTwuwp4d8jKbc9A0mfwhQ3MOe1HwEKSL37n/KMabbCdntq6afGn1nHAvDiCHVN
G9XbmMbue4ROJQCTK62/jxmSHdGwXf84QP8wKFwe4YLHjJfm2STrWMuVILNe06vHzW+HH0sd4qSt
GTgQTc+TDSPg0gKnF2sZfLS16Px4WcgakeIy6ZQRa3c8m1ziTvZvea+MzOgslVygQZ1IZDI7FNyU
nqf7I5uQ5HxC3AdCwrRqbwHG/Z3jBvI/B+6Ia4B0j05vF3pmR8kz46QPZWnJb9MPHouNSlAk6S6J
0pKOXjVwIIzQ6fd3GYImAKoiKOpfimtuDPvz8O1DpRG6zKq6BT6VeyOl/wMkJyRj8nlDq5pzOdSV
Dx6LaTphd1qRZhDJvIBadUWdYQPx04GubGDifAiQ8EuQAdrGnfj7+HRCGkJQm5S+JJQ6K4ZZKsjA
6aIfZQAD0J3Pu1LXqC7L2Lc6WcPWVio+NKd/+iIRLr8zlcdKLkj5dKunnUSFygnEUHgC9AK9+4If
1hmuiyRziUkoc6wFK+lBenYHUV6ppN316aYY76osMPibfAt/1ne3i+T3Qiy5yy76VzSbVF25Zmv0
6VbOfoj5ISm3mf/lhQ55CtjB3WG9D6si4usorTs6TeyqYx8sNuaHyezEnAqyR2ve/5R2G9qjGmCj
qRtelOBwGr42MelYnApF3BFcskeYrvfrdXPnYOHDtG0MWKWgnn8aROqZiEoW/eMX1JdPXuonD+SL
zqjtrnTxHQspFFhmLaUoR0iOEvBffRTmBE/jOPp9+XbjPeth5goVO00DCvrnmZz6s4qRVBi/HztX
yBdtDvk44y90Tu+CgoBt0zpOm6euWl2Dp34BDXzd0bS+ay2fu3HnqQnryOsdZkF0tejkdYUL8QV3
4NZq1dcQZ/y44VZkvb4S1vJifC1aVVtnTt0TXQQWD0MsrmWVaAWbFdjsBvK6Q8Abh2MEpklWDPFj
OYx2tClwvO45mv3UqhQBbFeJR0UGLmr2vONKA0Sb1+BUHjGCXFrTR93VmeJb8QLcwe7ytQUSR3yB
qOc+RSaY25N1vNGETgqIMGv72/hqRmP1UCBhgyfYP/byRCxuc+lnjxqVO3h/baex1fFBISJc5ZOA
dFANtkHSAHU6p9slH+1PKdSUrmc+QcZ7V5rG4eYeNAF2oaQnlEOZaaBEzpidU5TJEWTttZRrGSWT
sK7Gcy/mZZkxejV7buMHYxtsCKj5OpAsDFiffwdr8QTY4O8OwF7ffUhicjtVIhrCeVVAWQcP9dKr
tdqIwzToc6tYHQGGqBe99yF577lLPXpgTdNHD0WVwQXVRtQRLpkXtvpsJVxivhiKSlY0qAjuK5tQ
hPN3XBsFFEJC3DJDEQ0JG3qMYX3k7pPmD3KI/Wo0rtQaayav90GC+H+F8ZCmSgY5oiptvvK511nM
BAaZKhQUfVtHa3ZURzhGdwfT/eiGdRg6op6aVQzNnbsIQdF8X0wDflYfrluthKhKj9Z0he7zwdvY
2SGRaNY4LLTg+/6e5MmFA47rDZ1DjaxehqB0kNAMV1D/ube14yRqV4NK7NabocWgr5Q559pLiaKt
oIY0+2iNfz+aNNjL5eNO43zcMM3xuwpwBulQrpaAxCI72t7Qw9LCdkdE4UVS98mRfswkIToLrzSQ
JoKAg8tayTFh1OHaHdYIEbGSPkfemrl3PcPPuhrKa+tRZHtHEmrXZKTh23aC8dawiXohGXr2TWnz
0N9mn5MWIVz839swV5gkXRz0eqds2FalnRsvhu9NDNpXlHuaAzYtwyKFWm6JE6oFYZtJATK376IR
1JOaluCF+25ttp+OCvfUGm9Vlcp+U0/6Edj6DT0byOXzKTJeeJeHZuaLrsnreQ5lwOvFJq5qvOxq
bI2uf75uc2gbPUsHm2swf+lPGj9qe3IqyOe/J3MNPWFv+kseG6xxsQ3bNsFFeKsQ4jJzHTdfoK9d
C+YDuFQ7DxwE8Co+0xSJd0ONC04OmJUhlQ2FOpTPrwM49CmbZ/O6/eGPjV/GnBVbNNNTUgM2v2dh
dqvxdqUXOuJ6mTFmzrgPVcb5CDG/ORTeUYp8xyegW8PXcQsqhbERZymHk8gheShK28cGJJ0envcO
B2Bv+rIq9W1YTOcfDgG9rrCCkXIvEKknZeRXsr8pVojePFXOsxzwi/skfvvV7LqVelCddM/m1mkZ
Bp2GjIq9XodF/+kB0X2nPXXUqVh/0fFtdXCCVQCao5Z0SXzQAI76MQQZ0y6WkQJbG5cbr2+q4NHC
jGyukdTQAcOp9O0qAdMBX4xfvTC+0oOFJmp/bPzSJKoa2zCBy9Oa1awy4vikDVH1TtPb976XyLJY
1vrf++1d6vzVQPPlOyQJBOelbCwbfNuMgQTZ84fxV9/4A0yMl0qN6NGtgIRI0AW44WgQwEgdTJKC
n6vKHmDL3c7Xw9lNxqiTO0lU9JDAXcblGfuX1qZEF+sSW9RuYBBzBqLoPAp47pXz7VjnssVbRwVK
wMbSE6efRmSYXwD68It7u+jUO1/c1kXs/0dOkUx8j3OKyDgDSBfbR2ipJm6UBUAv61auarRCX9u5
Zndf+rKVTjXv7IpG9Ga3L1katI7l+GJSdcROyRyzS//3jmrPUtqE+68PFm+NpBkLbFm8g+WJuwfm
g+b3lRx/X9ZT8MUOJTsGhXJ91l4oU0w7Ecu0tGhW9slJrHePSCEOi2aQ4rRxAqr51i8xbA7r0AUr
lsGQghOxhWeP8C3cH4TuISMzzgKweOeHea7O7JjqsnTVcbIu1pxiDkrgMhJmhe2gCKZ9XJyx5k1L
tcv6v6nMIAlUZQPopF+66Cepak8VZ+7g84IPTDWDF6CixLoMzuSdytYHjXqcH9P7qOhLAEPKFtCk
mOgqybHNbYR+6UiU+zM0tv5UtQnvvcHD7wVE50o7/FmeAcDfEUjMlKWyXuyHcKvqiugFR64WiPFK
ynjx5UjMgqKMdsaIHX0/vS605iEHwJ/bpRQX7liUD9Og6Ro+qEZbU9fnctSCU3br/2cnOW/8bdPe
817HI6ShUj5iATTer/jnnMxhXqKogUFBli+oO3RfDq9E6SDCWzoqO4ZrTO7ZDgSkFdnFgxEpI4LV
Jm1e+p4samFcV+w2mx+P0qYHVvEWMlHg00KIy0Ls9bSd2MLx0CGoQ0GEd5Iz1jH5xTOEA0Lt9mkB
Sa9Qq1zdviovluNJ6RqI5Z5ZeLMLBRblTFiI4ZjW+kUJ4lwg76qF4Xfo+4TwcQputpEoZej1xQ5H
fE/ckIAIGeDKUQfG3if2SeFBvAYMRo/hc1qzCSXm27gpPJD/RlNa7DL2CsnfcUhnJbDyJyNAhy2T
uPfM3YLcP+McQX4c6yvFHmMJ693a7ZKFkTF/fppf71PhKGKQC273QsAaoIunYl6VQW61G2J+hqsO
LUHaH7y8cIsvWbDy5mQYUASXz4F5JnxB5Sj2PJkXtiBWEAS+EQkLBDlEfmm9gtokxWM9oL1xeRX7
HEHhmDQaJ6RmPl5Vh8AD9yhCqtUkTEaIIH8nhiV0SypolSUwnGuCwp5KVTwHCWt9lBRU+W15Hdwa
9ElA1Agir28/KLhIhdu+lN7QWK4Ng/zBYq08uhY2Lm244ZDF+pJOC5Joc/EB97DS6C/dFePDFs9Z
1e5Y1/hK4GnacT7MOP9lOKdDFtWvaTeF5SJ96MJ5AQXqhHt/obiXIT+G8gG/DXPg9l5WptuP27Wh
+17vB+NxoStan9ajVAtPwOq1jl86ZJJ7VlfzfgShDchwcW5eYFLINR2C9gXjcqxaMES2Qt7ab+6Y
IEE5WI8gShx5GHWBT2ps+356SApR5ZcrhpJ3u9A0N8zWcWs5oPaz0Q4L8cIQYmryqAw9s6ANVbbp
HceGOvp1n0+R8g7+Tg4nt8zMPZeBfMlSMA6zhh8b95Fm9J2U5GpgPFPSGl3nr8cU9SAQi0cbORnn
XKCzeMg6Uogo1qj2ISHeNjHroITIiZvQtGvp9UTh4FK7gR/AHFzQ5Hd/MLkXNBDLeodbFTERobAz
L5y+2ERGOiOwCR0p/Djbgje7hfGbBO7i/02f7No++qLhjn9aCRf41UxEP0SPOFYtsShaZg8ulBJ0
5+CbKjuwdQkqmWQJgxnf1hMNrbosZXlkSG9MFRuMzvt4Xiv5xj/kapemOFTi19Gb/7tm+s4RoZ5P
StPl6GIvMQMajuGUkzEC+0y68BBY7b04fFzZELcDlmW7rLFGSICZME0kVHvawyrtaFKD0ThamsFV
AM+rVrGx+XNL8/Iyy7tTz7sLYwE3EgnnnShCOzz5LZwo9Xi8olY497vwy9aNWQ8vmODSXI04hFuY
mqNmwv/MXaUbQp3JSbY2TFQNavFUfECjFz+m0p4nuISgMshZrirr4enH9PL4hFrfxXDxSWXmBIoj
+6/TjcpN+HgKNR+YElDHGZxh7EpYAm0c+0gY3MQV9v6064/XHIjnl5Zgv4PBJW9Eq6FXDdUmZcG/
GphdPcSX2bcDTNd0v5NMlWlEHPeIHkJ+pLajTcsNui9qbczDU3W9OGj4jqGQA+vaIUBqLlm36BYS
WJvOQYZSPh465SGe67tuj7N/Ljw8fIgZZ0dYd6+rjegCYTmOdD/JwSsFFq9b3S8ZkkoDcNFF/pUI
Igkl2rWtmabanoLh7+sB7AkzMlyJ0DY6Bti8+GPo7nRN1RLVXBqfRxdAeKcGKLQ09AVZ9L/ZTITO
a94oOfhABaL4L661TciLg5p5It5mlFOw0D+FH7o7yLcj3gPs+xVSQohEG7nNYIipEfoGa1FWstIX
0dGTaA8UTqbja4zNXtRDNnk6OFBHJquadd9jccwBlXXdrAmfzkkZLtalmqKGw6ATCNvi39xxGJcd
Kp5gNkJAHwL7EkfYhn7aYYix1slDDAdVG57ojgQttTP+3DhMuyKR1V8PhzdF6GBT3B/zxiksaqH1
94coMs60ZzwPcPdZz49EKn9n3l6c7GDfyDIsUwjD208+S755pTErsl+LtCld8NCLenu7HAbBPJY6
OyPt33jE+3KxBma6XP8/px5yGEKNpwup9uyOgoIhEIG7oRzZ3USLoLHX1Lw8lRyCFdXDfrnU0SZa
PGsEuX1nBJRX/eiqBNZTb3OoUpkIqmYX/mF0n+3ugPJf/zBP5Th7aBMDH1d8gjne4pwgobL2OnkO
Ds452nwJdC+w06hy3KGMYIEFl+Av+h/AXklCPrgE12XptjtzccPaNVuvzsxe5tNfqLYjgwUaBeGp
qzVSUhjLh7mhpfDpptIObdnYeVWwKeODjF/JvFOiZppsX/YRQUSG1UEkwG9ctKketqUwLIADtKR6
FQ87RfilnM0j+gKYVqLRad2gbU+z3x/+U3mUyo9J1wxyisvC10n75D9O1jdu47/f01Nlzi+jHzjX
7MB09QW8klbgVFz2mMp2VU8YxH/JMPlQh3J43Vi3MHruxE9p+s1uMuiC2Mukmlq6EGmiuSV+d2CJ
FC60/HBHcc/g0MnykTdYgOfZ6HXqUaiHmBkEtrQ2ryWI9MfMTjOzMLSa7FxSCQ5frkDjwkvxJj0w
GLHGsWA+vKhWkRiGziRb34J1v1fZmCcDzCzblGZ0GgsNXww5gMlNZSAiDK+qtdNvcpzu0UCmq8ee
j3fB8HgZ7wKSGWJX7QadLN6R2f3OuXxaklCrlU6fPI1kmuoOUSBZF4rjs4u5s2hqEBOtTcb65cOQ
lHscvc31zGhdrPDVJLlqzOYKFrhgaIJCvdJketwy/k/87+fXEKBi13YPHvoVIiPFSPpHGy9IJAgW
MY1wtn8PYyn+5jwTDL959QaaqeQQG9YqXdRNWhVjVT6q286y1N6RtgAnR6V4bUBLTeI2X560ba+6
RidGx0jGGoQBBck7jKHmHyj+h5RXLTrxFiS3SKOcwTn7jVVrbkl9k9G7CMdUbQkq9btQ4CJIKU9N
FjkrZBYIw6c1/TQZ9FU0QxdxQJHMKjHwUuCSFNKdw8kIqNhUsyMwIPAwbf1Gq+juglB7hU8JOHp2
bekM4AiSdmFyBlKGz1Zm6JeHECuTevmX9Iix0MTO5QJeUBxNO5//00tMYNFYL+ESpSIDpx2K4kd0
yYh61OVLXND1D0I7IQvyXZuYFpTdE38lyt2aO1NeNEwVK+ItRLKckzmBxyffiTICnjOtbt+y25fd
yUOLRFIqHD2dDZPhZ46mLp94RoAYKp1kAOHaBYXuJyI9JzV3kDERpjIiAOEMh54a8K2TArhLHidP
BflyAbrDxm/4PRzDi/64YsGjD/mBCULHQf4ZEGwgkiONyc9rVxCvXrxfPTJRbSycdeOrHVDbyhjc
0RPYBbQZ2kIsc6arFzZjDqvjFC+LOP6Bk1UBOzGG//aauwr/rLEJfEfEb+A5+00uLibeoUMLJ3kM
prcsdk8QGoHLNQr34ic7xAf3Wp79EQGq/8guoG6m7c08rAk4dE327mLwkyYVXEnrKq7MU2yzXdh4
/1EYInk0umDkqNwdmXSpBqK9jpctZN9qyc54gqnt/LQfQ2sVuCfZN2BM5urdX7FQ8kGcx2qE1yPd
JFSLOrwcZz0prBqWTuyi+xhDoQJl9/MdqluWRksqWcsLJ8ZOBc0p9Px24DoCbx41r+ssEKCcH3X/
CTVn+11A3E58MP5TUSC/inusjaPAP64d5+YlvxIHWWaX4BiagcQMbJWOiyZMtVogRKpeQ7o8rHEP
A0++3oiGs6bhK5THImLkTEtPxqPfGURPWUbpBI7QwybG9V4YgOfvYc6HjIvZl3RbhI8zDp3gNxOr
W0snoDjfGHJkCJH4GAdU4IIO41S0W9yGJ0pr3xmZhcy7kEGH4pCl49qPk2an7juXE2BAZXPopLqQ
7Jr6olufSGLc4N6t0G2vXmWICBhoMnDk76ME6il0bNdx+kAzDR2S2PpwkNdglcEoI9SX3zsB0S8I
aI5o6RvZecvTn8lm2Y/ZJLoDi1KSLC8HFjUCYjdCqe29UH2pWHHnMOOu3nSbB+FhMwgcslLQS6NK
NqF6NBzWEsHDE9heaSxZfL95r49hIZXwSKHzbFwJaM0a9M8ASRTTSnAxKtqfSoRY9/FCykOk/a9u
dcEhPlbzYfn10BTLH15FelmoIb77+WEkWZmq76sOVz+TtZKH+zfE9vEcumQFXoEHJX0SG/baQi2J
pDHtGv04m7J7BFjzGHecHBA0Wvg6nRQSaGEa2sWFPYXVlP/X2qA3xLyspnb8UX1fCGT13Y/X8P9m
NdRXmqnDXVsazVmAJXmvbjbDDN+3c8LjAtHyNgbfB0R2YHk0ZqZW5T2OEpxWdipfwypdWarTE9re
t5GvCfw3NKnxHcc9075vgiDF0navFci9pFZ6wl/0zlQED8WGsvPHAdTNsXpAQyseVF7gVUQREMCF
1emBaMMdKAPdd8Qg9H2ajxgYE71oGdHgiRtLcoV/utw5vahpDmFzaOYPysGDL4PFS73J4yvNG6eK
B+aaLShFUmTXzFf+7KxHu8vwC8U4JjHV8JYP7Q5VGN/euSdzEdHTqQl+g2zFEg4ejTrudBW/l9h8
9OnYF3p2KJF4gWc8s32kjYBXsSzrIT5+zHZlm5fwFFdUlnYir7vCjcielfRT30vEyjydLVge2REQ
PU/VsczskfE3MSmPAaERNqFXdsyt6+sTghhtcKP/WzxEqL/XGGFAlIkxqKYRLONpj4pqipjlhhIN
OYV298DXsYyGCDanOQ36ClgBurKWH7nVFMVbNN39zvG9vuVMBUXyRNCxYnaK+abZqCbvzy3KfgXz
Ysy9r5lqLH3Ub8k95KwK1zJstrgr00VaE1tPfK0r74KmB6/Ez+bKFtjq/kfb8Pe9MUAoAkFYEbHB
b61SkSkGPDgxh5NaS1tWfZF7BHNhK6g+3t6o0I27l3/7O1U/D95VznKv/MywmF/3ZhpXLOrizxtn
NqYhCo1tTAWFmZT8g6FZt5JBdeON0DyOLSyEQp+tnfujZ0So4UR4mK8aBaPoX7yWPWrhuWzcz+0P
Bg9M0snnlGx5OB7Z2fixwjX1gRJyB+JYKVSD3I4eYSYWKDri9KleB61tByn+Mz8fWk7WjZq+Xn8v
7ZG1veVg0q09ANqAcjxdiMunYov8526Z917M42Uyt2ZEorYsCDwZXLUCctUcezd/IyBM/t/9SHpL
pQiFgcybyruNRiFDsftVXj6DfGTbUEAiwJJv0cxCZls9ZSrcV32rzv13HMtdr9nBETAF827WDX2E
fzVpglCXSMqC7Lscib4B/iugEsJ3ST1SMF6S2OdlpP5+4vayS4XaaCKiDoKSaemjANjjxDCtZqFN
zofZFbjxff76VQUgEtDLa7FggW6rsDr3s9foB9pkRJrkEIW5xwyy9ajDv8/C8Q8tgEyEiat4L3rg
Q4tHSxiWMn6MRmHEka7oMbpTyys3osD4dkBXF9krqVAwuZw2f+TskdIs3hkwo7EHtJZkzwlRAvrh
LaC5p9DVFO4JuNUSv3Oe5ThFaroy3unGGXm+IsTF7SL7DNoxqkSC/qZXTXyVkhJBfy4TJ+uAtdpw
MyicXU/8HjWH2n/1EvsIb2tEGBIZLTog7ozR5pP2E9EVuqqgAxR9HwzEe2uUQzj2wcgIyWuOtVk6
b03WwRtqJvJN1FV8zVzEE/h7UoHjd4X2fs/Fx20zW8fGzL6oqvNKP+pAy1YccP8yQhez9ourR6RZ
5Rspfi9lFPmZFhirgvip3EfSbXbT96IZk7SXqM+2JwYJP/uPi4eFNZ+hLkLyWW9ngeZEu+QErMW2
fRnSqMarcQJbP+IcNG/rT8G6kPUrIGAJmOeBY45kwbM7Xdv7A3Pj8muD4/8J2j3egpCcWublPVgU
d9gEcw9IsVnw9gkllMVrwT92JZibyf+UF1wmTmhaCvW4Mrz6Wyt+15FRo9q9YIGxSXiR19gm81e0
vGTBr5C1x1Rtiiv0YusNf3B4pHk6BaB2rlF8dwUZMN25MHy9WSDuvYHI7s3T++HU2zwp2dwQj4Wc
LJ58YqF1PV3V6j4nZm2tSxkcF9yMGM+3IcSy3BbxvoGNgR9gkYGC3pF1/3tNFZ5ImT949fQBQhn1
SgzCjIQfzFl0zWbmG5WlgKIyZ2EOETp8XSKQ0tjfkLthAVmBiC6/2VJW0wcQo8YzHHdsZg/77JZ4
EwD9bK/m0AaDaB9OoXQHGq0OAl51s5kxMwb/u0B/pONy8yUt2EhS8EUjjnqRJdVKZPAXNN5RVe4g
wJY4CKAxU8Sm732I03l2hhaROXrBIcR43RyhW4alw+N0Gz6CE9SwMLQDkEh5z8EriN4Ndn9N5KVY
h2Ew3rN/rTUWq35wQWdCnasXnP5wegmmHal+YAEmlTqtk9eETrt89AkqNjJjKnb4L1kQmoSXBFfK
e6KZuimCqleKMUFcPDyJbDbJTGjjciwESodiGZc/ORvELeP8ldvWU3Xyk8RG41H7WaHAxGNK5Bmy
AF0v1hloYcBA8fjCkvBMyMFgQSyZkbSwndktw5UId6dfoIq45MK59yFUJtEq4/tHO9LmupG9ob11
ReX6Hf1KN5fQ2gG28CCKOzxxjJks8xFSUFn8oUU3SG22eEEEuvWxHjlNdc5MaJB+KrUXob2WLgtn
4y2EbdCVhw18XX58VLLJPfxH/C1LERhHQMODHvw/dvsQgvjx/M17J0zENrwN954mMW4C1RMZlYpC
8Iw0rwEXgy77VOiAk7EGtnCYlQaen71CUoX0HHSUjDneSoTDKuthkNlkpb+9NBxX32g7MUnW0RW4
2YHudfa3Fi5t18POFQu2LKWOXC+AkAgzBbUnrLA0BKeOfSFmgqzM+jltF8JYh/QrktS0WLgaN5uU
q7bnf1Ps2cvCrnTEGKZ2QGAQnN5x9fYZn7Nz02lRBkwwndWau/VPeqk9VOAsK1djtTr0G/Q9FGls
ZLO+bNGdwwxEx2G+f0pamsCf4vUMjNT/1/CO7yxSFbT/EyHJDUe4nbReW8OIlecli/+IZilK8Doi
AG+niNAf1MxIFsLoVYyLlraF61QmV+AmWjDHmqR1oUDqggzpLtpa12ztPnBq8hUdw1b41pwgHtLk
B0vyTb0OzFap9xrUhbVofIedymb/+5ebWMeJ2clxrDiQH5fdgZ7+fLVWNEfNepc2JIIyFeN/v4pd
exA9Ad1DIIcj0aWvjJEt/+hf5jnh7b0EXvpMnow2aiQ347NsV7XjRdtOgLS9WevfcH/7xBgTUK6A
d0Hn69Dl8x7gFYdy8Qj8EP3MZeQBhYtU/yPtPwA3YtPSwS0xdG4ZCmqo2CyvU5havKTCA1lPcn6a
UJdKyK2V52fbYd5+A0MPRILe01oPZxRWhCWFJlKsTZ9bSXWpLuo/Ji8IPB57CKJhBAq4qD5yCliF
fnU3SZut652xmd96EjXzRNP8J2+NzDZyS1gWnABvqHhth66OuaBmlT0LMBRWtOBXV2JWKx55BsJ0
aCSjdr4FS/uPvFDR43zO/P/mI2ooEC/I4V1bF5Q0beBFPI4nQsJVs+1rUv4Ltc15R7QlU9yRmCQ8
FqZ7x/iVecf04XKlyO4i7JokzEWDwtLjPvu3Gb0T8Xnx2Bi8W8LRKWDFwwfn/cQGQ1kKDICOJVye
hCoOX/yHX/lR22+S4A+1oKvGYZf/t5JXIUqvLaLdmjKRaksNAT9OXVSdUoc7I3KImF6Uf/MFVO9g
isLVzSpWzjQ5jBAWiATn34qrd5MMDevj98NiGDl0i2et3hxF1ivSqxirGyq9dUiXiQi4kzE+16b1
JMKVtFdIth5gHdVN+WdfaVkM+SU8l0iBdhuzaY+hpoPh0aDJfY0EWlPj4OlMWjxMlp8Ou0fXReK2
0ojGAtbWgMZhqzPOjc2444CkXn2X4+wHtE9p8hGtuPXOWyLR/WFSXfS2TpcAclzHzG03LjPXIqzv
zDBNXoG7My+AMK/gLzgCOoHcMx2miH9BZiqeXc89CP+1fe9e4kU54Ayqaqvl/+4G17/aBDGvTmrk
4lE5KmT00dbhsLkQVvpnAKeDSfPmwDlzLmU8GYMurynxxQzFxyCtTHrJin/M7xFcVKxzt9nfYGuj
Q6cVv0N46TVg3Jzbbm50UO1YiDoDwNPL5fm10fUAK85PHKexXGrfqyijeuiGlrtOmrV8OTgCkytP
/OxYGKeu1GyvBslyxksDyXXk/mwLvlZNOkGlSdAR69GVIMcfOfFtIgCDeb7ByLe7rsh9711E98w/
LJzVhYekgDH7XR9jhB41nfOs0mm1JAts5LhPOmeZTyS8ha0UtBCnU2cw5XxtMQ+xWvYxh+r2JDIi
4hfSr/YwXQD2cDJXTXNAhO/7OePUOTVSnIRg20cKkndbyES92weOAbb1ZaAPUKIotpigrQxNmogK
LnHZ1EnohbyiIY1D+GYgJTDxjS2gHXUAccBLx7zfaw1k28EtUSliUO0vFgG8PDeKpv+i5NQCNPTl
kqMkYa8HKUzAlwxCBGv8k6uJE31jLFsuiQYze+tVwceTsaQ1vi0uobBJwyB1siK0fUBv2oYKaFSY
l0aSWLlo2uJbVm6BWKVOrbsGqAhj795vy594B2uw5jGCYMyZCcOAzZU5mDd0koD/Q02RJNbvXQ9J
9vz4dqoQ62E9esyQH1D+cEw4NOGOLyUWaenKt5Zj3LZqMV9tRNTV+p3tnKUvHkfEBDP6JuuCZB8Q
j2MY/mYdsk0/Fv9WovpqM931SdXeEcVloMJD49FmrubOBxFexxp8gWg2syT9+GuzMQYOHouuTBmk
zAGaa3PmcpObrOPzGe8Q4NfEpLydf279yRhoIJ/zYynlKnAHdAVkxJ+1zXfZZuAGXUE+8a2obz4h
j79VOENHaJyaYsDogdTY3vCBMlYQR8THJ6qoQLrV7wRQ6M1qxTk5NMT17dlnTxXZQiaDUN0UA3FZ
eLc5koseEs0ZVIWBPXln1/lc6ekWROU7jZ8c7Db5PCtQzA1Qvxct5YH0jXSS0h+zoHRyooaWMZMB
yRsXfh10cuRhHT+EW8ZD+lpfiXS+NSUkvS0gQYGyEyGm+YaRQJ+YbpnHR8jemxkYSTTjc1nWGd/x
lg9nLeyAyVuLItu0wyCPnSHY5KXUE4PAi00/zziGHq6yyUJKJ33Y0gzSA4sWyfXNd9FGoFTEK+2U
hHEspPEZqHsE482NNMLwYQJrjL7++lBIIJWSI2X91rEYkzoeQYI1pKQCraY3spBI1G7xwGZbXH5+
BYCNxnZbKrIkJPFQXxehAqgYRUelX8bAk32OY4t2HqcDZyu/7HI+vP9QTlGEdNXHhDyj4tmt7m/g
SwSnLnA5qGxCbKMInClwKc5PIrAbw7+YzeEBTKTgaeYghwgOfMbKo9hQR/lz5vZAEj9/GeWu6m4k
XvtHeDg0hiAtdjVaJYxwtiiUDXZh89cuN2A81P8iTuyKKLD5fqwpUQchVXK7wQ+VnKnmPDK16tuT
WPgxQr22y89kSHzV9ubnR3wWdFAXEwLgnMLkFrzEX2sp2jfeMoq09ie1aXLz5FF/palT6gpgfvLm
2gqjlaGqoBZVPM+eLlKCBduxHSKzQ61RF7orde5QWJMgD6mDbxVWSZOEFCVLxVtzzgwBf4LlZ/zU
hiG/XyDArVax12uSn0YQO5uICcnu3RAdJtkX3pww+9r1e7dxBmcfXhJc1h3iTbyhg8ZzKI41+POc
dWff/x6cfRPHGaPAhWZS4HVmMk6gtHvQ3EZF2SWFMFYYVgy6oa01G32Hj7TymCzMOIKwBEaXDDXm
I9mex9gNhmG3XI+iiX2MmtAubCs9ZWs20sryhytOYIczvdzgPvuXCeKC3nIc2VP+GEzBL+EysDRU
ih+ym4dCk/KKetlAZpRmREgnan8D3Nv5CqkrbpLS0vJevYrfbsVxeX47XjYw7fc3UOakbXyONSKv
P63P/ik799wgx61TeU9fgZ/rLe0B9jalVB95SMXQ/h4LBzd1jz3PFegKC0zYlcD+bh5sOkqqMz6x
U8fAVrKWX0kQ8sxRsVvJCmZyjbUFdp8tbdU+GI+nHtCXAjznP6SJ+knCyuW3GUnlVkjSNWUBLFmP
63yFfbzLg54hXFzDP0fVuBfYA6NigOjjK9FDeLtVMgooOGSTmlSzGNxk5lFU9BPVNCifSDDIB8sx
RAL6Ev+TirM75PRaJoA6dHlBmMO4xt2v1T09YKxFWAbJRh8dWGt9fv1lzvs+SiLvC1dOAbsiT4AA
/yRT8TgmJ6CGU8cpFUEm3/Vh6PYlU4ccBQkt+G1/i2KOFT52VBahhQoLQqwwD8puqxIx4rCuY6pP
Yqrl2WvOW4itTsdfFWaxK8R/Oo+iv1GcapT6kyirzFaVmX5Wuh44la6Frzm9BQi7dFsRTBSXO+0z
SZIheJ4hmFFIqtnH6IkGr4lH+hGv5wlJv2Yw8PvN8wErKJz7LHWgk/+O1oWq0jS0pK8rOXnL86CY
VoaucOwv6EAwpXsFfKwkhkHOrHzhKZRiyBbRAONXCG5XH0mmUqqzzpOAJ0bEQ5SUeO2ubDh4zUNt
AOGcRcrxJiCkNPzRNoCAAZVg9a3NJrfGg0k/3Eeeu3asYCI7IFmWY2Ais527yVh7ltxsf1LR73+U
B3kT7Abi/e1qojdWDCS5tMrQ5uHZiyJnsJINBiUFMzyBvXQHdjBwdpnPCYoOmdAlhNVxpSTRufO6
1wF90ajL41y5nVKnsq6FxV5l356X+11pjmhYMLQfIGSSNWLvFScq6KmDsb1TStH0Ndy1XjgCnML4
KhI61tFej5ILs15uDikpR7gUFXjdQCgMNx2dbZ7vKJQGVPgKpAt0xE9+njlHx9Wx8MRm2h30JhvO
iLuFFeStXuXggFBBRkZV3iekWQI24zOQ4GoX7QsaYraUHBW4GL6B0dpUBgvib+Kw6/Bmd7pKEgq/
awq00ANv1Bj6kXDe00AeQqUp+6NtEY8L3XDUaJ2yC4kR6ffFebWN/w037mSl9zgfH48gM03diPji
26CPRMvJ1gg+iFVFAS+xilzQHl4htkxmxczudDoEeFKXIIeYGrxPTdVN8+JqwdOd7gNAVmUktY19
k5Vllmkv90J9ZhfpQ7PMzR3aPKM3B5I6Wz43BhV7LXTYjNeXK3FAI/5D35chJSJ7H97afr5SQjiZ
T3BtiIJ4IMhV3C60N/p+njHCLB7/11bWhFvfHj/IPXVGSJMqtqIEsze7QYKP9us4k4QltssnOb/E
Hpj1d6bN4Csawh3/YaTMr+CK//vqRn9DttWCHCulgjqSdHHjxMQB2iS5ye58Rx7CZontk/VzaSdJ
MOzSTa1lWi0Cd+YqnEZ+OJqRsK6mUAhxVg05ybj3ABG5y2lnrlK8L31cPsGgAby0n/tE+X7RD4PB
JNNbGK3EM9s0FkVoX2qkNtks+MgirQoIlq3OAEeDCn2UFii8u2wwRz+jVmpSAiYqrOBk4vt9eWkT
xzDcYMxyHJAK1d7gxEq7c/IWJPfehkNe6hwsyePgxtgfaSB1nq18zlW/Rhfb0pEXoPO6Sv0Ye9sv
0RI8ls0RF8zccLcrCOKw7e4iQJNPhUjm+guRP4PDjkE9712lUoVQyrkVO4HjACqVan8LNQvgD1vm
5Kklm5qkxnZqxuNQAl+QqpWWGM3bhqbubpccN9cG+feEehRc+tIyhnOQd/bmtzNSVzz8gBl9eUcz
lO9HBZ/GuQy9QN0D6uYfrtpPi6f8ptleAypl1Qhx2h+G5z83ECjxzqgTI4kN3b8Ir2nBQ2BvWFad
oEsx5limFrtNxq6S2nE/hhY7n97udk81sn6byBU72UgrRr1iTWggQQcS6tBcZOrlDeZ3etzlwwCZ
8mXq8Jk99tHHNpXAAa6vBoJ/1WbkJI6oiNmfDfXqr+UabLeeEtiTnKGDUoWHemSoClmiKcAmbMhR
/eesP5a9Ahr33X8+bQWKIGA7ucrg0zxQxrEn56MvNvXokYsVpABHeY7+8TFehXHPIQ/ibBy8WUCb
wJdIm/KZctw+9LuSLeE9r0zJpG23QtZrutNqKbD+9XbYtxRE4EFj4uvJwRMPTeZAYHFwCUNTDxRV
pXVfLZx1xWo/N/Hs2tURCM2IO9f9/m/+8lxoVrUGn/AFDoH4YKNCMu/B/N629B8uhV/np35GIimC
R9LSJDoXdH2gkV2Cg1o6y+eEtnpyk3aUx1e7LQ5pNkpHqMhoanmB2chKPc/egSUdHWfHBIDU2B/G
AO9Bl+0LtJx31a9S5Ga92kqnM6cTzO7tMwrqC5Of02YuAxQ/ObY76qo3783Ochw/ExcVU+LOdF7q
IpPlQvXNUWKlLreuS+xFVHd4sxiew3or9ELCiAQNouH3uBoLIM01wKFgyCmg3aptfcKsfemhI8y/
ZjbfYrt963AZKI13nBiaQie67mTxxRQNTBWXqMncYKEHnsnf+bRmngA5uF5AcDFlGseUbMpNm/lz
E7X3q3+JbC5nN6l0m/lyOcFuSrBScjoZoevSw3QlOjImNIgBk0IfVhWXjDvAmwfLj5wAhM0ZajHR
0FuFEEha7nwO2S3hqmRZOwNOR8QRvEB87XG17cOo7KYsrZAwwxAyN9Ccg7d7wxK8XKvfF7xtuzYv
+ZW8WV+v+g6wQXNOfbAgPTZyXViwHgQCkcy2l/VwfhqNTn1eCir/0XK3+hh8VZSLIr2iTtaA5Y6f
+1LscIYfOor8A0TspwX7roDaQ7yl/j+Q/KN9dJU9Q6e4HXGC9e0pIXAoo192D9//OekIiTcR+gBI
gBAmU5KoaWixJ1f8zyy7hjz4akApbtt4zD42pIBv7OVeOvqYmZnmQQLN2Pr0AO6Ec+FwccK4uRRR
2VH7nJ/DjxXuLn3WspW/pCwsTHKfu2UavZvYE6dE/rOXH75pj4jApFIaJiV60pUBYvJ6saToU+QH
tTgV2Jg400ifC3EU+jzDukU6WDf96NMjCSyAxHg4yfMEyIYdDq2B+JKR9VzhmmqpvTgXR5ZW9buD
4ru789hSXhU1oA1WPeusSwuH6rfb1CYNapRrnQkhuRSVlJuyvfVwh7/dnY+7iiuO5zLxrlPghle2
EvCaYVgEv+bh3/qKVvgl3uwPhT7AFiDQYYHFyg5NakMBIzeSMhGmvedW5X7Q4xUfHF0FUqkJvY+1
0qzer9eS5Z6LltdIfrdS86j+9AnC/W0j/CQZMy0N81mj26j4YFh5GsE0mBGyA0nF8p47pVdQi+ip
kK+hwni1w2/1Zx82lkYM0Q/saqVK1pnYCiiPYGoHZJwRYYlppGBddJ7zevEJIdttlSMiDWKIEe59
cVJNqv4Cb1uiy4RklV7+WBThOqJG8+IhzyNw1MJ9ddCBygDesQ9lmqpzh1X34/c8EEN/IIyJR8H8
Os3B6e0iHPi72M+O3XHVAyClNC9hbHlD4AOZsEMRSRcpayo4e53PmqWgr63lEe+8dBzG2pjaYRqp
k6kTFaaaCBi9zAsAyeiq9m+cTd9DxAoGMLmpqgwrXMMX67+lfxxMpB992RzGh+djp1nIrwYswk1t
rU03VYxcPeVlp9NXWolZ/4LyZrkJ8t8r/OsubnMhbqbC21YS6J413HrKMxtoQFdgpNAYlpdNqaaw
9VGFw3tm+c6OM28tnHrcf0A49Lo13h7RMUjfCwTWlvWrtjwQ4tuZtT27PtAKaeiWziax8OHZtoiQ
wKAU5ndxNm7cKh/Kzjb48DLZIhEnEEjk/4xdavE4ztLq1RELn+Q60LJ4ii9MpSJ2JdvvbSAj0mn1
URfuBt5HHCU1jVVCN06qrMXvsiEwFZPMVpUw1T7jf9/eqjFzs0hktG3irErTrjDLS5V8/Dck+FCd
j+fHUt2A+aEscxGfYQZnPTgwSdRK3b31Hr2xZsfdhtSNqA6jOZlQg9TnROfS9J0OWIg1n1D9G/xx
7GBOHKnufcodIdTDVROz7IArfB+D4BlCs6xLoMjnyIRoqfMudcERlvhs6c80NKoTkvbV9Asn/3xh
GcawYoAUP8zxQ+y8igLwz72FJwR+cUd+c16S75oIWilTz/qRgOHs3IOFEENSJRe+DVKtkgSm3ygX
n9Z45qbw5PD0h6QauMWV142/M+Z33duw/yQC71XJLEVE4Rk4fZSw3E7+wQtX2w4gDzw+PDZhD3Xh
iess5GHYCU35HdCeo0auOGZXJbr8y/23IOPun5byNBAQu+3SW4qVWbMDxBlLXAvXm3oNVp/KZt4D
7MJIRbvmJWD+Rm2l+wnl2/iUT0oXpYKWasELu6bh7trSSn+o3LITpqaGfDUgKzpf8vR9vpRf4c8n
7CRt+oivdDOSICjqJaVBlJFpV7oKWM0a9vKj/0vxt3wr1IcOYS+j8OIqnClQyPYPnKmDZdC5TsKA
nhXHBS2+Sb20Tbw/QjirMNtN3DvWqlnEcyhPfvP4YudkFaWGiVTFUV7xRJFWQsEYNFwYlSN7DjuW
UMV9EykP5C1nyff9LWcxj5WNMAj3dVvRi3EGEAdez2vCEfYdKWp5pS6iK6+MnxQr3eHV9kAcCMzF
nzz9nmn6axWsP/6RM1arjDBrADV0b65QwpxKrie38XpQuDS93D0XZ6Q8R4aBokPPhfio5FHHIpWK
puJtO+yrF+wFe8XPLHbTUzLnqt5Srx0g71e/cm4e1OTKd64jZVPbEF8nw4T9P/PNlA3In9+jryds
0lrKDbOPWSLO0KSx0NVqvA2SppwnVcX7MEi5OaUEouqgl2a2dtmxHcx9exff+sa6Oj/YExflwkDd
lIo+7y9PknsSYq1Ajzp4UYzSpRD9k/lhmaM2C0DvY1T9JBujcptrKn9221ZgZtA0jX8Ua2cr547s
Cb9ir6c8CHIbxvi4LLmdmjGEbKAXQWsQ2ZoIoSs/Ahon7Ky8gFARgPFXCpJerLpoqvgaUPAm5w+W
fhEy5njQNpNkXkeCHXa8D/5orry+gThJxvaSiei1mPCADa28+zIVLzUI6M+tajV3t95ToXBpR0fX
xiQN8RxwoTZKj5faRP+CFIJGcp7RHeSJNng9ZFu/gIyUvhKRKbAvfbpVnMiv49aFIzWyShaVSaFF
kHe/lVb6cdjxI5rYo+O/blmIOgJ+GLNpSMLAB86aeciTAIAGvGmAhuO6aB0mPEhB4vNvyZ31NC7W
BZp2H/+3jWO96dAeqf6AP5qWBKGl3LYQztrMyqnlf3aeaf/xL49EtdoWzJj45e4Esj/ifHBJNK6o
izMyfOtMNVwfUD4Ta5sIYWMNw+D/j7WWW5V1AEPIM1TSGJIPyQOwcUP9XKRoP2fWRyB+9M6ldJxm
mKXYE8WFiJ3S0vwy69SKKFA27MPmBd6mehVa0+TYmoh7XS5i5m5f2Sas2I8Pxft9BXwPjfpABqUx
XOIFzyBpks10tCjiMlY2h3w8E9iFjV3sWIiR//c4yVFhyMGmufWaPyq6uM/ABVcal91sSuW7nrch
EAit3gIuXJHgmKA/gnF9aduWarf9BfiT3LQLVi+jB9nRDMvBTsjqC3u62pcaxo0xahIURMt/Ivba
wqCZ3f65WAdx1Ld7Z9HbtnQTv+RiS/WaG5ozQKFW509AAmaMUPnkAD0OBKpIpPpuYRiiYSP7fd2p
hjAgB9tseAs1/p+QiwtaCU4KImlBpLZea0H21iLgwxYGu/Bzv23Q+lqMAFkYaxRmE42ntx0ZIlPF
Akb0vhtHtaG/0jFpV4mk5+Qgv4op9nUVZGJUMeT6wD5ijN9UG2zzcFGvm2Iso9dbH06yn55V36PN
E1qPgNqXcRB1WpY/29YWMCeyYlmHBoe9aZu3zgLqnA6xFJMSC6e3m3MLacfyjuAOqsugrshWGEmK
4xt5tIAj0W944K5LvZV7E6rTdQjx6xq9TRebZXmxIdb+qJi5qCSYLW/l4RrGymdy3utSqoKvg5gC
STC6PAq2g7JEh8TddjyK83OBs/twQPJP3OThcvofdvgVv7FnvIgLCSYwrXtTHuqZYtvX3CcFufb2
dWMr4bT3ScJ3ZVEXVcLybS4vOEhDr1tLj9ix6LD8cI3DXsP12i5IgjgnO/NIhBUNVt+fugvcCYAQ
9SGqH0D1OrgAvKsKRCTTKtqiW8w8o/2onOys7cklikJLuPM0hwBNMH/xJScEIZcSFXDZycRpu0h0
1jg5L9jEgrBbMldDWXLxPScT1q3AVcCMuwg6XIWpw5Ox1jxjHMl7NLqCQvnoRreiiBEfvmccbo2C
AhJe7vLSniFDZfE2VLNuVjE+SevsVz8c+sr4DBZdqWsZhhas5KJQD6T0GXVc0Ev0Rww/ih7aMFmE
KMtHVJC6Au8b8qy0C9OJeEmjx4Z2aBssF1k43JZeYMNTYID2ekwiVzgJU1aesOnEOCGU1EKvlrP5
OutrbX8ERNZwLrl6sIxmgm1k5TclCTEpAITJHays1bUZic50G6LvBadLe3HtYRTp5TKZcwTjID22
Dn2q3U88A+8b+etVv8oAHfGy59FAFe9oLn4kbfRA+NLz46+a68XWov6Tn9d+UxODxqSg+8uJcqZy
7bK75YYbnDmY46lFe6O5IhXHGMPTqvNfrvjFB9AKUBCt843xxkHVHzFOs6QfAIn3cS+rPPdHiAzF
ftMxojvrxiedqLacWNcj64eD55ZMAAL7UMF0JYqKG0SELRShPiXtkLnhzI7A8IQ+N+h39IZ9dXkq
AXllQWgMLdnFtL0u1PX0pIpuvvlpG6mjL5VfY/njhiPewunH4Qcwj8V5AWQxsJWJ5NNkJngGmhRx
TKgZrtRt+WBkOPzwAJhqoxipiFW/GHFjSatAMMmNk/2SLScLqTwfmKGnGw1ZrytKyYdBwLNNq7zT
LbaxUrR22faP1i7SS6dcPVlPCwq9qd+VcTflKlQbH+LZBS2Hi1vTWgn6W5He49MkU2WfaTwldbE7
bzGFQDesUOLgqxst/fQNEP4mkK8VTA+xcAb6912+qK56giBQ6qIozlg88I9juSUOy8q+LQSlfGDS
MotH5/2hTgMeYcZSu/IFJAcz545+M/b6kl89iPlWFgkhI4PM4GH8s73LuiY2zbT+Z7lakY7iUT0a
aZyPEdOn7lHWbDzwEsPmMii9c1iZDhKTyhQRDOVhuB+aUU4ZF5pDv7nLNX2L8y4ENrdFM6KIofvp
ra7O7XKrEOaqsF8ToxdRUAl7VqUr1Lnd60BzR8r/8ssL3g0c0x180va53Cq3cTuzjuT5avH4VOPx
yyEjr0ivVW5mhrUf2C9LIZZyVx+dOj+rw2cPHVOFKk3D7jTtT+9AdTwRQHDhP1DmcCPOEE9hMUDO
h3pTAAu0AIhO+l6A26PcpHAhkXGSI3BQcV/fz13WkqFgXleLatgQZoXv/qZnOgThCQ3WCKR9iO38
5NsKYsz0weF6PB9O5xY9Mk3KwJp7j12FBWEYoUV7TH5Zc9xY7H27soJGpj+4jbCWYhWvH1a9HviO
k0GQO6vmZ6gPseYAh9RLFBb5YlKKoAZCoDm62rIWJjzorFZud/ejSK8ki6jn4qHK40I5V5EjcO+E
W13Xi/5S6f6CCw1gQJFr+89+fRQTY+EQMzY3wOmDZLxd5TQ92tE+swHKizSLjGsbJcRqN5WRCDbE
bpsOgDVA6TSyFJoHJbrq8J8jw4wtRSgwTXWPZE50Qqhk5PbydYuKfyZJV0Bs0PhY6y9BEaxtGquW
aM84stULhCRyTIEd9Utqqj+wKQ9b2PiPa+fu04mMRp3165NxnxWKif8OMYncAPW5DPAX4Phqtc0M
owi/VPfo4fsKWvc6+lUDHHsNdrqDZA2810AjFxNyIKt2csmdWFE424+2MNgcJJtpVVTURda3Q/Fo
7t0sSkba5FULnZzBj3oKPK0hUf5vyGVNMZdaIcXbexJgYu/0JEAw8gt0bOzd6cKLx4Zj1dc48h8M
wE+sgtPjQDwRZR66Lok5iGuVKFkMc1hrrqSiiVPcPS0ek2NzAfTCdhiRPcK8VzxMrLNLWQVhFPWn
Tux2WMpMIrBDCCZ9rzcYAh9pbzDJTIqP5LlisKL90yC54arXOzDrtTycwNufg6j5t0ZjWOITP5dV
SucHKRJHndoTlnTG+RZWhADglbdsgmVwL1ElLeVQfF2ImSPih0FXa/vJoQZXg5oi2Oyjgd8KFO5Q
um0KRXNyAdh7KBsxfyKzRf3ocmDz9YSWhGdEnoaU0xXH+ytAvbJR79IttjmUpR+9d5/KaYi60fse
IPtQS/4msN6wgFol1hLa4doXEhf8uwQAkIKdkOzNsVHMp5K/RbJfnu8BNBPSSnEICwAu3g5NAdqg
0rqPKSvtuBj7JvLCtAKlBbaTk3KKxYD/PiqUGXv00CD54J55lpyEt0ypDTht8+0QF08bfTwcz/HM
Uv4b8ukHF9EHp5RdsFU4AHJIGUzd7DuB3gcu0ccOyfxTzmdNUhNrjXoAy7GmpxmRZ/rtTuyfdUa9
5p05/wQ5tdch6fnLpZrmu1c8ACEI4i9xuNLc4XlcrvlWX5nF8OGrrR9ZPGdm5Cg/tcl+3PffD/Jw
lknB3mdz4emdMOYXqaVweqEfDyWQIXH4zfPbYkyLsZ/7lOoCpzfztLzDYghcBfhIxjZHMR6Yu1j9
f817XxgcSxOrtkVPP32plBBqnyaRe8L+c3MxSq+FjJ2F2k2ojYYgF6JrL7IDtAJ95+IGvwL9tzp3
pHZTsbQLoUQ8jKIHkK0Fq98GsKlMuWDqbxPeM62JluLeHyucHs0Cq7kw30GLsTwZypOO4QORGyF+
Buuzm4x31hpww/NRznIUbHsKGuENGRCfWCPMEjnfR/eDoU7w0pLSobCib5w6IqjQMoVjDBwngvvq
iuHpWGHVGf4ZEtuxJC9cigQz5Oc6f+fTX7CtWEbDboY2p4Carxz3vvtV1KzJkcw4ToQzLtepAQlq
QPN5ctemcm/x07nv80E87qB+G11F8pdheUC74+1oOlM8IjcvzwoCIrYClc+Ic9cjwo6FViCjctME
9H5eAnE3V5OvbJhncgmPj0QW+ldpO9QWreU3yTsk0ZEUxUO6GkAifwaY3DJtsd7NF/X4NUIJQBrz
tzdx7UOdauw8HcQ0XcMgeufRFdj6lcClWh7ofQcM0R7DImducuQsUSR1VvXU1ooecu/0fYtpcK5f
5FCzUe23Y+QtNJDdvnWOnbV+qQD3nDsRyykf+ssi13Ou0j6hvBbc+QysJt4PuzlIlfujz0kgskYB
tfDoNv2afeLdP3MWQuKcQ4bhpl46b5bbTFZHM5NfVe+g+0Fbj9+NREy/ysQXEE85kUHB3kkA0WH6
EYvmsViKrRM18Nh95GmNEq3xlH4K0zP1a0Cel0QEn4WOOBdfcqBG1ZsVWXAgLIChGA2+n9c8WnJR
sUmAlcxXdrycRLiwNe0hV44vr5xPGYrY3yzpUSKaNn0xFyoW4SAzPpLZknhuNLJqM8JWDTtNNifB
oieZEkmyA1dQ4GsN3JVeb6D0TZdxbS+kzo0GMOKtds0IwN7ixXtf1tqcS/VGtVouoNbhoD4jTrLC
4fAv82UG7SI1bJjZCrUieXr2EQ85n1qKYQSUbQoEHk/W1fOiEZeu/6J8oMLPUjhTIa2XBJ5Mjsm2
F1uN1QlwbOOQUEe/GaHSSqqjX4KIXx43FNA9Gk/1ok0/OJMkPYNGNmwP3sz9PbHFA3INrv5P2S36
50U3VWPR38juCpy6x9/Em6vodEzVa8Deh2qiW7qT6dsVGYCNEjBMkd79MJ2F/b37OECCZbISVXXu
bxWoBithACQm3vyg+9mJgD04375M4fR5TD4INQ/Tr90IXdiMxtrlwpWuHqnfW8NZTHbiOHYYBXGB
X6eEdxnY6HzBgoEVwPhYKFy4wLDRf2kuN70amSFjLJAmx1b5aCZgtYpYbOA37M8nAndkwDhfkgsK
bwbDXooa1dyQQnf0TfzorvKaMnzX1i823NpOL9kGvK98e3Q9SDtU2ugk1X2Znz12fuFG2vMMv2Mq
cXhjw/YY+pVr/rU2eNNCZf17x0BD57AVf1FYTDMNkbCF/yS+6Kdk14ZEzqi5gpf+5xqUwY6Tm+xL
4hyb/U2QNk3rN4ePCjtj0aDIo6E2kZq8SteVkwzpRrAYP5liN+KGOTy0/L9UrFPuBCvu/C6qAXaa
4Uv8A8YupPw81HyhJtsTnSoT49ekWuZa0gFtlhxfNJ5VolXWPyQuRXbkNPi1keGQDHyH5cSWrdeq
bdLMIkt0rz3wTBdbC18Hmbgn5sJ0areCXmDF9v/cGaSPxAx9QeonL2JqSCQ6YI1XQ+2pk7DYp8P1
jMYEKZu/uT2Yn+H4h9nSp5w2KrNoXQrsAmZ2iBAzRkCX4mr+QXvMwbIJPmYOa8IcCHmRJ6DI6kpU
SDJonVzNGf2Site9VXI6YynD4KwoFz2woskkI2as9B3WAUpJYaBvkBpTJY//j7RFt45zB2fF127P
I4LG7JCIE7cZOS7VHJRqLH3nKy5IP1qwsdRCu9m9wm+zwBZQEnUvvJLWYIR8Jqz7alY4wKUVXpiX
t483e9sDoPCUCGK4hfLMWU3i40FHvyhqD7i4i3KHwPF3S6ngwVw+cErBYyg6Sav1KOcdHM+cjnca
HZEmSF1xC+kmrB9L6c+MqX99zFsqloqmk3ixbFI1X5nZFVIofHhAdPeJE/C8c6RwuSFrnn1WRRRN
HHG9JYiktXKcsWmYBJPzMPRT7J6Mox5f3VZCICXpjsBwaRjiKfXTxObvVfmSzLHZYst29GEerh3g
Va6j5tU1CO1PxLTcEF8XTH0ptKMWOYz8wRSwD7EMeNIItWCBG8VRksW+MX3BN+tY2O8ORFPJeWVj
7LNFUjSrgJEwYLKbvp8LRuJ50HNAT8xceyO6kzmIComTsMOZ01jP8uo2BRkMky3HCl5jKT4O1Ev7
o3tjdpRaOeIj/GAGfZfxA+ZED2ZJLZJta6QUZmpAVD61zJHj4Y39NvalE+s1l+DyEa52drdq0N4Z
K/C+cbLc9hEA3u2NxpQKFoMgNfmt0n4RNhZNFmUzWyCSdSWFIW2US/mQB0viw8y4aY61vVK5Wnfl
BHBXfCft2Z/RR3KF4B6NONrhLz4qEHWVRhdFAGSNYDZqBx9B3qTfUFc4X+vO3nKmhw1etih1IhkF
NIgcLrK9Hx98t6yTZ+/QimkPNApIQ/Zi+78OZUWIm5FYde2/cbfLrQuNMndru92e3FIwvjdEAY6p
IPICye3BX3GOe+P9t0qZU0UM9K6fxAJfc/JVNMrZNLLwcXkisEPMVCN1QF9ZcThra2v3vao3U9NT
ceyyK1J1FrRkOFVa4BmLGyORsnIMuIxrGSHUgb4fP7JiRWAfOp02wP0wzNHKNTtf5Q8wC2z2DWc6
nGQWmEqOMdY5kgdqN6s8uLu9j58k5NWUVv2sc4EIFwfPXmYul+dgAcGVi+M+tAbADERERwGklYAP
9WOSdgWgSD3yDdsEuA5xSFzZ+he/+6XylVPyCfpvkP54jS067Do8FqCs1PJ5HYu22+J7sJgL4VJN
TO8KtddfhU7Oh1n7vUXZVa/q1wOw/PXEdjMkla4gr9UNSHifdpf8e9EVcqmMTzCTM8mWqXehNYE0
p5YO4sFF2E5PAdNxZ2eC5kHJ4PuPHjrdmaL6o+lvNyujHUwWlE/KJWR24yac2Rfk9/MZAJj2SzVA
K9YZZ742tAdYudKp9xbxhC8tRt3TbIHPjgRjObTpjB1IuZDITTx3IQqwqEdKQWY/4I9aLb8GTd9L
A2jgWYImAiNh+P7HV8QindaOBYLv7OUPTSXvjshjNPXevb4VUF8WtKRyRZ3DQjXoWj/hOHO716ub
6th3rJOYDEMF7a0rCs+1UvY8jgx1pcIKOYUku3pL2DruvssfBM2qK67VfFWEoM60STORWqeHqA8K
rxzwHOMPtnYfEHjqKYgtZJFBBX8RY8VTMt+GtKAmvKhKB4jN7/3BifpeoOjXPapHl0lhInKUnXIp
KdHp+82QLvUFG1GMAyJXnqjf1qQ7eDaLbxQtfdoCmdaQy9oYEbQjgxD5ueElsR+b2PhpgWDsG9qv
BjWfsENK+feXwJXH5G3yIrW3671vcqsKQBbCZpYrSARBlcrJhLwvll5ypxofEFhrFkAKgzegqNS7
PXGFnwPyUFMfaonP95aNR2PegASaRCbbd/IZomyxTQ2OaAjSPzuuOR06Vx7/OXacE1g7gQF4ZQVv
pwwODJcObh92c7TPU9lQqcHUoPrO4WkhlTR8NDaMQJidA4viFn2dyHNKVRo05JZYqrjaDKNTDtLu
L3rNAQZuhw/b27vyHCj3ZoaiF9l9tMDd5W2LnydDZFOVt0FTUuom5GF3k+QHx9/PdGY7yiu3QSiS
iWFl2qZ++eVYi+onmJ2FIPOcmc2sOk5SbE1wCpk5AN7AQNA4Ac9PtqoCshj+HcKN33oGQMX4F6Mh
6e5+jv7ygzFmVSgzU834kVu1X82x4XMwOu8/zq/x+p5+M6Yc6ciNGCSufY1wkDGKq8xW0C+rTHjn
FJU9iEw8SS+BqarJEO0e1nhh/oK+wMAQx39S8NoD7TyuRpVmPrBtLCzTcfXWAFlvlghu+jBkhP+1
acpz6mom2SnUbU1/hxmGBrBieqFqb3q7Ct8G4Pb8QhZFfAXtaurSbD1YDkZS/k7IDQwIIntjdsDL
NLzwwlMOEj5ps+K0qb09AUKo/5l7k7bW8i+PwFu7OH0JORfKe/wAil6oQrAuqzn4P2a59p0A4IQN
c+haCT9/ybAFcmSNHIMPzMvKzGpdOaQNoARXlOeYr4pffV92TFxpz3Y3NmS9JaphrFwuGFUqQcDF
jRV7NWu+GXZjxp8XXNwZOhfjZ56zJ6HNA2a0PA/Ol6O+La3jAXB+Z2bU3KiGYbD0acBiCxrDobGC
FgeT+X0B4Rvc0RBQyqCQUYbd+WmbRwocCbVyPS+qBhatTgNzo3T7/mN+mkzQPfkkr5N43l7Blpc0
rLRXckRkc32RaSv7uOCzxZv84LjREviOu3kPVdCEwAXB76F+Iqw4ovwuNQDpeZoLpkU+qNzN998E
jWJ77I00Kgmphl282YVsP6y/lueHn282B/IvoHEFUSD/oJLpNm9pog/T0KLbTkC76tH9PCQQeaut
wf+bBLITcmqfmDYtEd0XOqD99RjslWvklYUEyYhzBO7X6AZfd34pS29v1pUrBPaHRjl+KCUKDqPO
RwKHhTQXgCybgDPX2KiN+AV0RYVpvS06xcH9+biF3XKLK1dzad+0zChynWzSTb29PKQSrDD4MKOv
GfI90GC7jRUUQlQZKmigFd62eoyvxGPKyl5+6K9BawOLZPWxFlsaOUw1PyA8Z69m8zg6FU9WRZ9s
FoojXSKSyzuiDLnDQfuruOpmsPieFZtbBZxbj1FQJjfcCvSYBJ/p9hwr3Iw2avWo0OQqecBklmh0
E2/2oClHAesLs3LJwiyBuF31Z4u6KRa+Nv6lu5+7Mm3xUQFITgGHP+rsmkM1ArQMxJLIqfetmuay
N+h0oa8GIIVE6zE9FvBNoBitPMFkTd46CY4UKcGwzYYu3ntvBwukY9Du62n4p2XCE0mEgg876FnP
y7KAdAJKSSE5IV2brXEmBZq0MCw+QBn3koUNvYVXXl7pGCgDEf3udjqZMORm5TrlRdtg61Etytze
pCgGqmADpEJzbZW0bJzX6791OxgoBpqg5rZIiM0z80HLRZ2xpFY/5jv88TloHmhj929ZZSuyuVA5
N0+80724tR/K6dD+G8sHhi/kN1NLmgTTSUdAompB7A6IkBkXEa2FrnqAVEBndYUqXWXJxF7Hy7T7
cCWbZikxmc3BjdGaLyn/gWzHKANnnaowXqD+fkFIS3GZcBDx8b6PKAyS2WfTAyTiWRvXox954NCZ
Pk4/EOFinQ3BN28k4cTSon4FBmMkGvemlNA4x66BCew20KF+5cLDRnNOoeLpcDDJis1g2nYJ6nax
zaXwdn8E03KJzyfQ6sG0dIavujWnu/Ow0M4Qgu4UhRTXZ0blqs2D5nWVJhpZGra7N9oP8A7TFIop
X+MJfeTCTB5gpAC3bJWnVVxUOGk1ptXzStIsMIjZ1iCGos09ZEIu+Gw/NUUvU1eYG7uY4q8zMzaW
IUyNOCnngnWA3jjUDLrBNMO85/7774W9hzOXfxeGoJZTzXARzo7l+Z8VqpzR70NN32+DuxDkoZMZ
2S8N2PhQQsFcMXKBmQl8mmnl8xrEWSfJmFzrfVntq9fvnNXDVCduyTHoTYpBWnJUAgIoXtYdqXSY
y2tHmGPj8BQ4OIfmVqSbW2pXXzI1D0h/0HbfGxlEJSzj6J3fRDgNjA8Nyf8TbuVFrU/XiSDvcu9G
5m4FGYm4VJDN8bkRtWanGoE3TfWECXvO6bbNtrnq8Rebukbfa+7vKbefiV5JLCRNOnY0C2q8dAUx
fZG0UhrH0WotbGxmFpra1gqF8Zm3Ju01pIWRTvrTfRb1F60gvWkx9gpvFYY4ozdxUHc8pIRVkw63
+DxuInAa1X3+vkT4nVGqD4Fo+bJ9nWu5dP2msJvmx7UIF/E2jWigZjyuV/knnzjUjQBqPDMiAAFQ
2/g7YXO9MArlCaPeQLuviagN9zdSvF+Fve7nXuiKkE2nvNVAXnIhMuGpkwhcATTmMJch9zJ70hoK
fy+rCR4XZpRw1YabTR1PgKG2k6KWiqRpQ8SxN1yRg3ofOilUH9a+J7z+govQx4CyWNdI7UaFJWtH
4CfOCaytVbgFohdHsTehdcLqTNrzoSPsgZTugKVSw+tNzDCDvrvJNuXJ5x8VKhxUFMSgBixg3lsx
yMDVs5MzoOUE6GpftwN4tD0qdAYYacdzOfn1ZJ2WlegdoSEOdKTeHd0bG+v9iRZnWqRTkld/iVSe
pfyH5YomyTBQCU+z+PVUzhbLBOSOIfa6J89DDzVd9PQ+jsg49+/38x61gMuYweZMrTuD94NxFq2K
ULF/AVfGOv36zrWEfb9N2QrztijW5zStU3ojZfMQJxIqNLIntErVfyAk//G+IE/ifBZNRIfijXf6
4PZSUVO1jwwDWmXKqXx3rEfYNY4LbUHRbUzv0CDEhNczoS2D3DEPUCN+hNe6N7STg8C1DDT68Dbf
OpeT7PvztvnxKGHsVzWYa0ZTRzGkBuWjhuxCOdGSQfZwyhWVahF35vdrc7+EAopEG0/0fCvwQMDA
AeipDXXyK2hqDzNY/BhzBaEjcLk9wqNBjmrrvtD/ggWnoO6X5rgGSZhyiZPUPN4Pl1KF3yAQJQdY
OBT1KH2HmUlFseJDVyJHMlxnbWVxw+U8GMGQ7Iljc54xk0mir/x1Bkr0UYnveom+s2I2fNSXaP9R
Fsy8Z52W1eU3Eo0dvYi9tZkI/tYTVqwCDp49qbbob7Scfv4wWW33iEuZ7mbEBgomht22fzqTgoqn
f+oJLhp07sW7p9zwb7SDOnIAJ/EN2aST+5GlRDWxAXINoN5dc4WVnIK3kQSqIv9MHFy0PuSy6Tzc
wHfwK9QfK1B82xTODAU6Wx/vfJAdlxKSbiNJil/PCCKeiW+cDe9Nf7dKzi8hhrNEZh94gyC/vVWc
WLt8F664dn9AIIgkqw2FMXcXWxJZWVgiFjpBoTcNj3kx0uxwwFlgy6V7WbG78Sopa+H3NyVqkVA2
pFYYrTf73VATBRMKjuYUXRzE/Lg57ivoNtyz0JMVbBI8A8PPuK/LpByxKMKa2zb44QgYmYhz0uB6
fYgZLlfSd68FrfRBgjydcc41HMBdV6UYFCPcewaujItnPQ1wyE3AsLEp6ASCvDL20JWQLIsYU9CH
QYCKrkpmVcQeUSq7oLDhjJohwsz0Vq/6dZwsr8lLj7UmQfX47daKJIMRDb7xhdMydqNuTpvYLwsO
F9RDpwhWQ+MJBbLNlfR3r6fL46TqQwmxdFrYR/a8p657oV0NCMdvyW7Ua2UMTxYbLfjCluxusvQY
U7iSUBWrv8tPGv5a6zyqS1zBLcJ4UF2nNlVf8f+9hPMG8nVUeoAFPaTdwBHytoWGRIOs64Uxw/KO
m69xiQamLixMEPau6Tie9JaqN9DJ9JWMirSDQIf/nFF0SQ2IY217sDdTp75YLtFuzO22p4sbVh+a
2BMbh9QuLETkt8UHzhnaeme+YE9w0x1SBt1JsYW0oexD+pmLxDAz5/0rPvndVBDdetZj06wlLyMH
T0IvGyjWSESFIymrnc8nVoqHI9wkMTDGafdI+zTat2gYM7xqfygzHzopCjPHPckY1PhyU0VQNJsl
11YgIO32vyqKbrrmtQiCcfqt4cC+tw0Gmk+f6T/1/f93ozcVQyyw1l6PHJHNj3YeYEkkTdvZuYF0
ibIouSuT2sSCz5p3MjxFGZbid+6JlE3QOJ2/ZXTcJ/ylS1wwKbGUdvuRNif1Ft6h1bkVAMdYvXMg
X01ttlMtMqn01EtNuc1es5/3xnDGifa+JE9hp9i6gPBX1viNUbSLN3vwKKsySznNx5HdKQfOUzcf
vzfXl3eJgyOQ9ro85Rpk95czGcjXtDmd21mSToozSdapE2HX6WSxz4fPjySLAPMSftqAHbPnn7TD
KdDS2QblG4w+jI1SBToW8aj20VknsEsM6AAbCes267vyVUTM1FU3Em3CukGeUH+wb/1oQFsKy50f
q0deJXamp45bY8nSjfIF1tfyhNQ85brwEU+dMGHoIbily+3kva6I/5dtwufgIfAVRRePrEKEL+51
7DwoeYMpTei1ilX1DbvzpbmH/v8mnfuRN0Jy3QHHalN9TRCrUdCeTXAMBk0VSHM95mACmgCtKMG/
Xeb9viVncO2r8CYE6eiS07oTu78VU5i0JYBDkyuhDFm4ab2w2QZCLwyJMlNS64Ws1C7+PzZNenCs
PW+1FeyoQTHfO10eJjwnT6j9Dmr11HImkIME0f3sG5Ly4aPExqB18NJDpx/NGEikNZP+oqhMa3oa
ZLIyiEB9a4j7wpVeHuNAjhDmXx9U7hrahWcB5lrkuC92jmVJKOSDYenJ5jEraQDH7RYG1bZkE6gt
j7zHPV4grktO7WdkKsFRqgbm6ngC2Rlc+4Zi7h8q8PkzHhEwiwP70h7EhAn7mRtXsodTToRdo7Q+
MBVBLgNpRsTpI+7VoPZ24u0pX39JJ0WCMGpe5dPtP/EP2sxKxROEoLLluYLGh2Fou/Zx+7RFPX+Z
a5FhFcGlh1nodGKSN/QvaqLTCChnHnjrcsmCToykMR5AbylDJ8fcBEJt6/1R8Qr6UBIgCASy9hFa
5d1xqWFVpPYNADsTj1H8UPvuhBhfQ3J0+uroERZSvmSjQakqGRB+YEyQg1SA25+HL50264j54lbs
Lcev9f8qTAyx5XXG9NRkmSpBhvwzA0m6LosURQkpFlY/NfVW89ViQ2RIR9ZMUZZeW51Y+smo8l1p
h+f/WIEAOjnkVD/mveJh+Nc/uHfyifyUf+odIznz0C1GNnW9riEQafMuGXpGsGsvo1u8hhdsakZy
XiS+To5tU337ma5jaf1tSup1CCDnNhUHO+sSaf1EuoW/4KCYHNW+2r7dmtcCpdrSUxxkkZe+Y3C5
kl07lLhzazlfYjz6aBCcGroJDZbmMs9xL5GI36CnhbdHhT5apBWKXE+RP/wjh/3YSjC1kFc242N9
ueK/PlJuddN+z7wO0FpZa3vUM7gpcL077VWg5eqECtRbW7S/Mq+yIewS0OSLpG2GarpFySwAeM6r
wFhamv/koEUeTmUQWtg/UEaZPp7Vf28BEyLviSGNmESFpCBru2Z6heFOo5l0NBhdKoErdGJmhaUJ
koxq4avpjQSgSMpFaDK7JdaFWGOSsOSxqUcCvY0uMRz4OZ35BP1lqqvdHI01H+KMeYdQrZ2rshvJ
ya/5zHIrmyTKETTkA6nCUd6PhROX1rDkA4wagsScAReHiGzCYe+aIFN19fGXRLb9amGaX9iN8yX+
zPYMUTpV/pg8zw+OJegiNjaOdFPIEecoBZoIIwxAuG89zUpT8gG0ScY/Pd4actrzZ6QxJ1U6Z3F9
2is1aKqU1KxesiPFhaYvVQPwyI92+1pPmmXY/wlpLqiEQtu5s0/11n+EZmsOwkTX3oHV1kPlzGSf
BM3P34A2qRtuAbG8P/PImH1Rs2aJT1A3b+HWi200NavTsLKRKxOcWnGBjg98odhecuZa01VUdhrT
J9oJ+9I34m6BzGyeGfdjj+lFC41TUS3KZyOyP0OpDQy6zpUb0v1vnlt6vj0S+XD6nUu6DpOTj4rc
V++VcAp4PDzAneAz0A02hhOAclw48G/zZHpRG8KpWbIlO5vbLQR08k4OibgaTYgqRA7wPbM1SkRv
FPi/sCNXR3fjXM7GDwJeHSCmQxMcmc4IFjG12mjT6FIQnIsUqtRBaNO+pn+OFZRDdVEAgI0uVXu0
qM4y2Bu4soSIP6h1dh9xcihm25/FHIJuqack+9bZLS0NHYogJgLLmhurTKqUl7yQWsaYnxYqzOGD
oKvposeo20h7Qg6KzdqHqg/U4Axu8cC85aUVGi1r4wCbzk7EktOBWmfHAELQtgwAkXKnfOPYA8QE
X0VpGT59iqag4wZBzvYZHAB0hJ3VB5R1lsCbw6tf5IGbALeaiKm4Tottz87D5O1OVj7iwrhp0GZq
8u86I00+T0ukema755CZcWfcmDlshtcLWLy/p4VqYGOqGPzwk/8D8lZ26hV7yqvrAetYTCLp6dTc
uyYZ9eK5klcE4F+h1aeBPsMl0bfgKfv4HSte75WV/feTOeCQRkHF3lRkkDwdHgaaq+mamo3hSsu+
j4kYSU8NDsXmdyiXhiZUJzarnwkeJGcrUD7FN8D8bvKHXRltYBoCeA6bX98N63uWynPSt9dnIbnA
9oN3vgJHArpxPuthZk1rDnaZYgvZ8zqlEkYHPb0QHVkmF955c0YDbIrPqOvvnj5YOOj1vbCB00ze
j9LAC1hPdAEj+SqYnDPYvgyeeSo8NvcvMEA/udAMj2AQ8TwfOH30+ya7t/tk9u7HodZztelAyfv6
RBQre+lhobp1+40jKK/F3TvTpeWpYHXVwVHddyjzPuZThd8dRp2jVaOkqY3hT0LdAgGy/+gjUXvX
dpNtJ7gJ08qAAD2msXmqqGWriBvZImnC8IIskZPxK2faoQabzEvkV5+Lrrv3sOrYATYFBDJn7DaZ
j80UTeeIWgd8kMnYcywHaHs5k9jCanZtkwwx1INJeHHhqBY8MdHadQ7H5TaUA3kWtbcpjlpUoF6B
vJW84m1tZPBUUK2KHr67B2E180bnQlFfuIhlJYf7xD3MhZvInP1OVJH3iZnXSIU1CyvocBcmmWam
QnmOcgOKMz2rzECeFRQ521FEv+Wrvrvi5L6JX+5jeWJpobjlwG4/y3djLGpoDRQA3/C8/q/ERZ7a
QI7XYsTmWGIvZ0ijgTrAG6g92P3xoVGeQBJk63FxI638jRYpPbTadSS6H2EApTrJZfodR+I9grFH
XX3iKU6U8qiNRh7AHn3YMp+gWk5dHlT9UP03C744cuKLPXg9dz+1voQRqE6LTovTtNql9FfgH13v
1LdLNYDMHYq+O+ckSMqXWk1wG3i10NAYeAXDIMVLtRPsn3taw14S/IzSgLdwafmdPj9C9U595Q3K
wW7zk6hzkTyVMIq4KZj0IvIrifoHQHWtgXSP8132IkwdCeq2Th06N3J8U9JyHFwfGW4m9L+kkHID
fIpaOwfGqNPbt78iJ4zjGt+4YcqNR8EgnOMNU+RgqQ2xoVQtz6shsG6LiLOCUWzwtdtQPzN/6PMo
VziHyyhm7KefBGDm+suKDFJq81EYrdvDsEK+sHASnrHXTkuSMjMfteopjWX9owVlk4CdjCAMM8Qh
shYU/CAvnQQPfmQ4Tyaz18vP7mEsSx6aLIafxD1CV6w74l0P/QZLwThKEPuT+l/8yQ598TGMwZtL
Nfu19ntLs/50/ARKw8DuGDMKXIhQzmVfMRs0KY8tROPxE/od7sUIsNJgTEw99wU7E2HOeHkG3dGE
/HFe3IqNC7yyanFN3mycmOAGOilR4xKKOaROa1cv+Zrtn+UjA+o7NbBNspbHFOnI1fJyYZJti3mo
L/hL68KhoFTft2leOBY36B4BIQ/kr5qv0XVRDeF98yQBmTMiQvXtU2UPY1szTKqKXTQ9uDneLQQz
UDvpcspyt+XDwQ3ZFrTGRn/5q3Nwh66IAKlcEXqs+dloAdtIfzrbmE4DEeBCEqJSWdRKLRYInZeN
SHSn2LqaOVzMBGxEcCyEPscBP+JfdWi61kBO6HnDoc5NvpX1BE0RsH4n7SANYsco8ZYNLAs0UF/a
9DlskApf2nY91jIAgJJT7sCBAXVsFZwjf10fQ1dthYzJxV8QKcX3GILsyrc5gPDwKnMP4qD+VpYb
SRIxVs5JkTsJAMG79UPXmK9LUKhd/R/Ix9Zi0O56jzFYyWLBC74sHL4b3gdBbCpI8qQqL57NDtJq
nvNFIN94zTj/Y4ml0FJskf4bIcyA3flZPXRH/vBamwXBPPcUs85NxOSgLULyCXo7AaCxhsQvEB3B
S9ftDv33iCbjTaLo5sKs63vSxqrGjGvw5gbg57Lb+VKi50ILVGT2VIoYhu8mvLzaIROAVjd93SnL
OpYItClZ2p4j/xlthp8agt4iA/jlbc+mmhQGhj5tGFJ3k9NSIaIHXKhHDSExFuUhu3fmhxTm63ie
tdlDKComwOkwH0pI4PlX35uH/oDRNUCBa9yzHEn+8H5owAjIxmo8jUNn+L2PnMc+2byhQAyIwLOt
CBbaUCb5nyaIxeGFUfTwUIC425odil0vaBk2Ci7TAE1P8kYUAByEghJjNhrTZBOTBVVcMj6ueTmJ
Yjj7Ausqud0mFDZl+WM+9w6keKqFaxZVnFunjwlk18yu6V0G7VS6CkGDTiFLBAt++YkTjess0Y46
i7keLY2cDyUw1BT8BYP+8uRDc5sZU81aratE1WzGndKk37KDEP+GhEngLaRywtBKve4Tcr3oCjIf
dBEaU+I4ZURb/k8/OliDx2P4Svl6qgrJAQPPhV8RchXRDKcTv5HaD2IxdhhcOoZCDlCjPT56p5rb
hp4rKvw2oaQrQt6cssMCXPVok1VDGf+fPRMbS1/BIiJA+LTqOPjFKrzzxdC8NTY4DSclvApWrjj7
gmAYl9TaFfIOg5PlSJFSlNqiZtCaPtLC/3pMCIVLxmSkw6EfEDMe9sBoYwV8x+dRfk6Osaaksbih
sINafdVVwVbsWKcdoIY0azU2hgGjpTZ4hOvqZu40mGMkxQSIYIbDMjKe5oJD/NM/M1ep0h6N7aQ1
YLRn+xabY5DPSlF7uMcLrsgjp1t6mCMkYPY/ncHFoM92fuCfs+V5l+x4ZuTt/zw04hZJgSEB+7+c
poBMicvzs6EBB7EEG+1zDmiDduM95NrLN9y8iKB80NUhCsVHIQjzpxCy53FpAhXyiojNZG4qm9Vi
FQmcLdJLGHrYZhTT2c5SaifU/OHltxGX9tmHsqUl2iJHlU6iO+2lrIvgu0zR0iNBLr/JDPxERvQw
85LBbtmdCS3PGkGm382Q25RcpEDOIlx19OLEcz/ggtSzPXjKkXDRZvwFDTPNbMT/xoUbxtodsYJQ
y9eSTXQ9BTzeul/dLVxQdgAp9Q3S9EZfJHjbMdKVTK4hNRBsUSV4OK2StZwEI8ArllZI2m1U7Tef
KknWbPFimlfYIgP6mha/wQNwA3CVxMwMJfAjsbRHqZ6/IN3ZMLKjz+Xkqs02FreXiiPNvhcdbAEU
bFtzGl9LSmZtYA8OpZnqlXYeKI2mW4AkPw5EIVj7VCkk/DPG89doms7XQ6MQN3IGwNACmOS3OazF
AqiEKQj7rbBjL/wPUcjU8rTx9gTII0CXgLs+Tk91gvnLXwZEiaaGbf7uQsF6H0D475KJYqXkP2yJ
DlWzLJiGMDkc+tMODx19gkp7fDbKh7QuKkHdKDtpF3Y5DtiglXBHu2pR2qzq/fbxgp8M4+jUDRu4
X3WZRxxhq2ulFaYRUkUZH+5QZyrLLpBmGrZyOMzR+fDKNGDB4RuxrCtEi8kcTdDUNgTzIYFdHbHe
rLsa45+RvbjWNlcFmdflvJa90Vq/qu/zj8D/7iWOUbMlwPY6jgIaUKV70856toUMFsA09Xk9oDqw
esqyYX3mwwyoF2UkIQd91QNp8OL61LqjmEdrpqBW3DSwrzAN6FP8oFChEvEJ6jVQ+om60Oq5+LIO
2gszaoTLso8t3XdPNtYGMgxfcMFXTUUHF5uqoveHDVF5dD7GLh6eKF1d06U3/I0bvm9a19IqbW4T
EkhYYaMOZ7MJOCvFhaixnA+4avodRs2OcjvhvurHdt6A2EyQ1lvM1olGlW2f08UXJeSDy2I3uIgj
djlyl9qY1cd1QeCKBwQkfZ9xOhESsVVWZFp3n2FFXqdLJV3tc059xjsS2n1ySTCSvSIHJUHMilbh
jtwH5xviBy1PFNhQaSK9S6eDedYaNBqNvXmnV61KvcctUET6Wbfm62GIewSw2Q3natAjDvRevR7N
ZPGwcM+SbghzXJ/9dTuHDNvzUEMTg0mai9jUujCy4Xnv9DlLfh+xqaHiKstL8q1hNWY719E7inqD
9o3xsTxdUPJ6lC4A+DDgTiDHOUudPGMqdU6NCJXOeGOSMEfxwmUJ8TmDHOvhw2ePBMsUWTeNY6i8
uDzg9KKm4GdzNYp9HA9bthdVNxvfF0rCFKm79DI4TKJpYycAVFZN7VsAU2TRX3PBs/rZ+q1kEimA
d0OjfHKq8yp76SPexaFOyV+KTeeqVvEh8BWuoB4LX3m2XzujmNN8gKR8uPWhnEK9IiFrgS9Gfvzm
wt05gahsVq47AABY0aOqE6+5n4xkcRJRPeT/ITIwfn2s0JBfgEHQPW3yZlIzwIBJiVsXQvYpPDIl
i1gANHk0zzovVn65up+aTzcxCLSz6CTs1LHMI5rHc/SonSSenMFtu/IfM+cmjSgJTkDxyJrcHPXe
xPdWWm2MXsgFwA4jSVwBnlSeuFsybzejcMdVvQQznZP++gBQSYZrQ6pgjaB4S/WHj3972ZbT3Xrh
FSx+E3x7S1bFdpzw7wLukZcRlwGJE/B/NmvZbX/J2EgAsgTrGwLf3IsGbodDWqPuw+h+w+c/EItQ
LU0UfvzsW1dE3/iE3IvuwY0BmzBx2aF9J04cPpEZHuMpiJn0qbQnn5k1Aqnc1Afac97+DV4SJn7G
mX+gYMyvISv9gZtuEUZHYHiF3d8xVQf17L2CrUVMTfQV2st0YPj1U2+oltGRDc2G2KBQOp2YLF8K
iobxSXqBvCPp7hcw0YKrQm/voARSL7zr1wmnnuXHu1zRODXjA0iu1/C+8Q7BSuwZ17oE9H5rTtcN
ujY0oPwNjA03dHSJ0rVSeibxJSz1zbRjRgTtJuEuU2y7A+PKcbeuMbgo2+g1/KBJOfS9wD7nZIBj
Kda5WY9MZMlmhSIl4DnDUvqAYUaxebFUU5qVMHi2JLdrtV/R7pNyhdCWEVkkc8EdogkeWyzPiSpc
1CzoBdP/XXVdGUMTvnm6ZlPRRc57QFVWjCZbFWYtm2QbYh5CI+jvssI9HUXVkDnQGCHJ2Jjx+6sC
GBZ3c7VXx7CCEUPm8Zf59TNrcaBejgovAet3Xbi7JLXXOSp6oumlDovvpr8kmW+442OxQolkvzPD
r2YD+t+Frncjo6PUaR5Tw5czXfmXi5OnRDCYG0fRtm2iX6BJ8SlFtT8AN0jrTUyIuNkJQVwL7cB5
BtIoQX2t4i5LSoyc8EAt1vKal9xTHrwDQNG+21LLxOwuFUxfanlNWa026jFPKd2FttZxJqCG9+aB
sWAzGKkyJukhFywDjyCIDVB1r4SeHTVSnoj7Mm/jcu+GA9M9Uta8yVpt7Q95iGjgB3uyDzfQOyrK
oySbCERF2WA4VEzlvRSbwYqxvucQ4uVW3lpr0Q3h6/8HdUJl0KqWFWqNjZvN130+CHzfN/YTeaBQ
THyPR+T3wd19+Or6ZCRB3Y+dd+4NkQ8e7xF/bwou7YU6dEpi/HuUGXAO78PXrgaQXec9wY3NXZC7
e6d78GXO2vGqfcYREEYX+s/eBlq0GrShYKHSDFHukVtl6skCcWaQpTn1vD+g6Vond+ze7N0Qxble
RM9X8pn0XHOLUTvYy7SqEXR+z1DA0xGCnYJnSvIYXBwnlv9dTgtYpuBBBktauWmD6iVGOB57pRwQ
gTfeHq2e7wXkrAUIh+LMxbROWgfptGOZbdgYM6Wa3W+ndymJssXJ/Y6cbihAThvayQ4Zgx0VX5CX
dpka45AzdgKW874b7uo07eWzJWKMroR/mo1oZxPckN3aNhPaOJp5E95TvGVmxl4nVUYB6x0KOxZg
2OYwyDrDXblPnTv7j5N/mGQxIeFf2chyVk1YFvEJ9mCiUk8wdA6SA58cd9bhi8lCSfuNfxX4Ckwk
iOlfCUlTcGS1xToUQwWsvJGLN6+w3t5v8bNW+d+psxnNgw1E2r9PKL0n9PuQmgxcPtrzlppoFLEi
G+4X6R7Hh8LRnM8GVBJ5YkVhynEiWWuIjyPStRqUyrpuwktyLrZtT8E3ytBy+42tsZ7Se2l2id6p
lMQOXntSGpBN4gyx7W79fWMftNKBoDS0H4eQ2pUOjS7LQcmxeLJ9WTX+CTO6GptyjPRp6YpdKklB
vO5+mu+Yv4zKt08fF6F2itTDEmadPHKCQ2eBTIYSVf7+AgKSZIcKePgkLarf2/EBpUShbKsnAWnA
u9LaaxE26fJfAd62PXPboAL83rMGHAdZer/EUg1gBCz978e9X7uhcyCzTtWY1sHzKCtrjHr79RHr
qGp2gz4jmfwjj4XYjLkrJx/IQta/n0pfLM4236HnrCD/J51HP9HcuCAn3yWg5goFIhS6gFUun1ja
54STrHcSnObYe/R3cytWfBhRiJVhpU1SwXfxbg+vHGKpnJTPnMcZziy36F5ZZAZ08btj88cDwGTb
K2Yg5q4dd7+Xsax8+n6aITiva2KcE9QbrBqh+fwMwa7mGXaXq+/iRm4dtMTBvCGDTeYokMblW6A9
qqVO38bu5fce+Kmr9mAcbK4YKmYOjK1bZqHmpWWDnMjrfLDdPCc1Zyf1liSbwtd6mX0sOWoeFUYF
pMiLyRWsBqjzKUcTcKVM5LmZUGtGY1qpMiOWWM+gNQ77vI/za3VbCvgCRAe77b+F8lxC0kTUNlfg
3xnJteutQa8XryTF6hb3+mduotHHuicJY/kiubfJLUuPIkXfKHiuckfKcy8ZcbTsPoCcfR1tx8+n
LXvN4lExHU7tnFaQa9vT2GY2cK2Vcqfporfuf1HXi5KbAgD5yCfbb5gh2IIl5+RlhcOUTJiWYOSq
LaMyJ24jIcAdAteZh1EavZJGuBzGahdHa0+ew2Boi/QKyGmju35q4UeT7cRIGiHHpmBcagysCWF3
5cEmicWxuQ4dUgLITdJzZE9ZhTBgp8KceejM+CuDx+ylF3pbisllsyibunOGYc0Jsao9XdmKaEUs
hWRpU0u933wsiQPuGK9XnYubRSslKi9kQNCn/me6SVcZJUicZ1DKBgOUocKY3wJ61x+Oi0MV4kum
LQRGy1IjjvOz8+ql2wpD44yMs2KVT3Xl4dRiyfyGfcRJVGsgUh10sa/oAoohg+ryFSHh9Om6/Y9G
lHdAPSzvkVWANmaKZW/7+XoEW4dEmXGO5MffDX6XLr74Nk7jFpvKq5Z/bbG3L7JNqXIUQ5N28254
6TggIU7xB4AlPjhjH+SKg4mo0g2VPR5gA3yEfICWx+UWmEX3ppxxUv/1XGVR/J3D6YEVCy2g9fBz
niKIr9bfxwQVuh9vbde09VGNEVx6D2Av+0bZWYD+4im8BISp88nOOiTzYzb3gzzzJK6/Af5McYDj
v2p8SWLEFSroVndY/0Vst8ANBJfhPZ7V0yDyRV5r+DzOKXqqCcWmtq/lnBhk099ssogGo6aOokgV
LNxRtaWcn3coAOmyDh4Dcw3HFfFZCkd0DPvmg0IT2qhFIvl63k/rBhr8gNc2QjgMIWgaRM90xSGs
dbRAJFutY7yhFwlpVS3ybuNwyTsnOYOy2qFTfphO0Maw9hh/U/VmwvwOONA0Lzvwtszs72o8NxYn
fqwHTFmgBPa+xzRe+n1p5UvjVaPiqvp5V+mv7Qyetzr9VnDwEHLL8LebWFnlcqqvEBFGVLEcIFiM
/LHiZ+myt1pfOdCcv0dNsq18Tpx6zsUVA/bL/QW9uaU5PFdPEDGi5U8LVweiGyKGS+vWsrEQTMML
ss5bLejIR8fQ/ZVZZ/jbr56vvwaLbLrBtvwLDOFKk9jswRFJTJYAmcn97uyTRElILSyav7COd6jw
BbYfQHCmaYnOmwBmCnWSMkoN92XnjyVQ0/7qzdaGhqBM9/B5AeXIJwxqmQLI1pofkTdiiDcyfK86
XRiU+odtLpHn7V9ESMSD7dZHWRYAmzQXk+OyBzGWECvPBMvgB7vRSekQPacgaxTll2r+EG3OVieL
4hVRk2xrmtz1XXwLJ5cVMviRvI5HpV9AXOgby1cwKKO6vlIiualJc1hpES3MtX2jVA7V3j+80eez
sEkqrOL31To1stdwnAoj+En/hKl9JfdC4hnf925el3Q8Mwwx3PDXek57s+zvYxkSsejvt68GwZ51
KEwznjTmZp77k9b0pUZCLIyFOlGjklQa2AfRCEL0XG01W3VCFBcrlatBm2kIwuOyT0c9HEYwScdg
wARvJMu/qv4VqoWCxFrCScxSNaNJY0rAfzslxKpBXMitRsUjrsuLbXBxakzyPXsdg0joRaByWeqz
xxuS0TnkuBlDumGj2ucOsPJz5pj5x0Tu4mFLBIwKr35zQsNjran+9Fhzlx5pHqxXbTFACL02DdUA
/t3TI/yYs8gWqr0vaOiQwKDcTAX4k0yl5H3lB62//6QtkNAa0f9iSGIdu8gNyvGsDt4TLC5H9XbO
/gf/pkn7Uob6EEtfgyGbC78idPeuWPolLGfjCtruT9PYShxc6cIyMuzjsllWFE0sllZ+6C9E/v+B
idKKZbs5WEO5PHP/1DJFAtobLaRvVnj3fSCuz4IxAgA4pwP6ibRhU1kvG5yoomSJ8741QItLi43V
uLEN5h8u3qy/SmV7qu1TjVCxX4dDozdobkXEdCZ1cZwiuIYKGYhMXwd9lWG6x0KpnOQXRGBpCYbU
VFDkeIcssTLG+rC4K3kkriQX+3jnqquImQtF3+iLUL2+3VUgywAxKbnAp34jm7by4ZpY+jMS4bTA
XiwGETTqsZt3oL/2tiQhqWMVLlIP/Tq8x/dpeW4Lh7tkFxGcch9jxfmTuKwoR9x26NcfuMzeuCX+
EDGfGKcwEW51SExRq7yJT382X6/kUjIg2E1oQrYOZEU/A94XHlSu8eNjWbPxZ42260N8ENXbmwQd
F7zasGzvc4C1+ZV7KCJu+dm8jaCP2cylt3KGE4voVsexH2abJxvXlpOebzDpvqxWl1sVkBq3I4U+
OBV74/VjYTbALJnaO415UCBZlQL70ZfWVcdijraQlbv+1UGbs6zxQTdCDyGd3mKxKAfJfJ3xJFUk
JdYNUrvfH1lhDve0k1PGddZznqou5L9lJ6LXupbEOBtR1OpE2wAPi5aLiHDBW6xm+s7rTz2N8Jcw
kf/wNwMWVU6wcDFBD/+atR1KzgPfCGSnx5bwJLti3G0p9uifoN+hmXzl08L0IZiFaLAjBnWqn98j
16BYn9Q6MJJ1Q2P5eNaf9e8JAVtstFc/Wd6eF0TE14CNQc/c5JbpSr8TjUUBCtTx511X2262lu/O
B+XjIozwO7v83mYGic3sklURKiRKPJ0RYszspxYDKedrxFbei5Tex99yp6Z2K1rx8+dYFVOKYJEt
Q8Q741/I/VQXL7rV03TeBk++z7bYCz5SdFtkGzBrHMkOsoNDaQX4rNk6WyqZ3i97R9C/6HR65nhz
Tffjih88yfsQZ+w5OzFJVgxTpyMPCi8NtECrfhKuqB0/SSca+KoyW18AUeY7D+WueiFhQo6bewx8
fThl0YzwSILdNF2Bi4iRZ0KSoJmDWA5mrW8seiWnEysSYyku/xOcqhQY8fwg0WvSuuiq8dyswW9S
3JHMkZf2dKNOX41up+M4rn6C3ITs2ywC/QM06g3zVShXQNBRTELx3gdJuDyjW4C7LZki2M7cyt1s
RJdwb4m9jw1/OChZLyK1nVqp0PBJwFF0+Ryplzd5xLJ8EK4zfWpDTdFa7RvQKkty7tVKw46EtJJ5
+Coh4fzz3E7cwofvLK6slwGienBBjvrB+/ZZ+KmN7xaBm4Jjb6Mq/Su1BZiOGLw3DwPFmjXz7NYx
iqQXZ+8yg0gtRacFkG8+ISyfVFrecLLsTSOU6Fa0hIsdN6BRe64GXWUI9IJasZFRSPtfzihN7Vgt
/Og3hG47aafNTWItWXfNiAJ9V2ZqPX9I13IWIipU6ZMiHeHUYkAT1bjWKPfU9GPk0CR6+7UcYREO
FXy+78I2MhnC12qbi/ZcMrF1Ly9CCIapPajmTQowYqTRfrKb3uNrkctrUtMo89YLRTb6SPhrPREM
Avai0GT13l4ieBZ39Ll0NPtJ9t91EfUKVdGK/PIa9w4EPbqUgzRAUmpnv5j8gwh18YIZQcWPwAy6
YspFmK9jP8oOtSub8CkI6K4o+Dt+IZzOQu2/AKHDKY5k8DV3ddZVvRJEz/DHeiQxlvx+sRPyi5FZ
6Y/EmOssM3UnkpImROF9bNZztmNVHq4yhAeNDTI/uD6xd3f1YCLQh0q7xKNGIjdaeKKDsmmzVoGn
E/qGWhXqMJ/Mt3DWpbVIV6au/FxNdlP1VtETvekos0M5FoqPi0OSUdYIL0047P06T14Xi1r8OxBn
Qhp7rtWMCVgQh6Ysi1QEjRTod2p6PP6jm0L2IJul9WoG9mtSF5RFidEAaqCp8NYW17sJGL6UEkrR
VanLz6WEknDQPbsI6SdsliH2eK8LyeTxSl4Gcf+py1JIy6vEJZmcrZYS4woREnshidyyYr48LqN6
YlkegiJFgjVIz2lTyVRcwcDt6yYkuATrOnRUZfnkaRf5UyUFyViGm1KiwV6k7rpriGPbt4bi6Q9o
YjRNzpJxKYnJhCAxCLATSi6c5K0szIuIZLLl3a3VMf5Bm3slyMQyfwsnu4gNmFip2dgQDnxEwmSt
S/pSE0SrRK/Z1Jdoudy03vkbRYuVjaUZZ0iJFmPgh9Uya6tp+Q/z0sSOIYbT1O5cOL6dsJ9/1TX9
NC7J9hdrnE5fSrTwWjHWblyd2suokcF21RDXuTVmSWK+qCjQ2ENuLv364z7e9IqZZuzc3k2yu7pk
rHk+TgRDvy8XMQ0opiqPDVFSqLHapinkPTFkRht8dUFRA77Da0zIvs/WIdMnCbbFQjSrUMS14xYt
6Kf5tvxO6DVHymXxcGMGDDfJCx7l90CmZpdxDLAqBhvbkx6MuqFYSwMkWylqbfRF9mGQ3o+UuSwC
TOPeQTf3DtjvXeIjwPI8BSHhX9EnkSp5WHt12vvGKRtTPx57g/i2VgAeP7P25BUHKpQUsRbqyE9q
+0HfDrU/8RMbqdD0BK77KNW+F1Vr5fPoHIFvfvkCI3RSqhxr9rTP/P3x/C1qTeEn5O3ZgozomzVO
6VeM+TR0MCucTu2VRK/nNXXaf2dzI7PT8b6awka+DdQWlQHgobVS5imq4bXeoEVMu0cs+de4dFGo
OmtGIynaPTKNuWpbOgpg7tiGbcDdjBR7pv6SitJscj4PKjo984m4Tbu7T2epVegrioX66E1R1X2F
1Z1WBBLSUsav7g+N5XCV3WTbMiG/QMV6tBe77JVddvsR3dwvMGtrwM2fhx7uE3v7BzAHkhCkh+rH
jQSoweDcdKxZgJ2vLH807Q6Da0HjuYiHIZSl++MpyvQ1zOqg/dRPmUXf7k83hpzJEBI2SpptZe7a
a8KtCHaaH0mLtIdL7Wy1AZ5gakAxePvhMBdZqrzbHjwVkp8XjM4Zqe+7yvSQegydEEi7UpXQ+53X
shjl1fCeg2zTkhxj3cUecXBFQ5W1EdD+4kG8De2dJluGVBrT93mzLFUNbk3BS1zTUGM/8yKu02Oj
PvBwMaySLBSJan0NN4tKKj1fFpzqH8ve5/rTPg92kEeS5Srbe/H2/PHrXntjLVIM5T45Wf8Lail6
5OTJOlYRsBKRP/0HqMQx9XBK1p7JYTPnvXCxHPRsfx4FdRHj2M6gHb7Ag8ptSVnRQabma+tKG+kI
O3cI67y1bHWtk+Vh78m7cT7u8zNUNUtAirWQFJdGUXi8W89c8CnV5mGfGOtUMLm5JnD0GHzLB8IQ
UPTeJBpBvBn3zYN96ehrTPp5pIe32GpUXiiafk7rgJ2iUXZGVVsyHz9lRQbjHLoxJ9DcbpQQS7To
KHkUuk/R9bBxqcMaALxFdKgRTFM4hFvKDPMN42PlCj7wl0fslqy+7Ga+XiaTqrg6UJ57nHvbL88a
nkrk9yk7lcTaTEf70EW4j93riaAGm73p6glwLRMaknLt5Aduyii4mbrAjkj2PzkxAQzZAkPCbPo7
pEAfv19GcDF1RalRFsFd9TJ4DNFh9KnjlE4Wp/iCLoPkyfhpOGX3SYU87qLoGlb27RXFh8OCmR0G
xaIGtNwGZnf0RLlXeatGvHB/WSOTvisHKhLPEo93NjxkJq/3K65i3Z0bJ/7uJfu5grsiAxTEksqO
921XNycI2FYqTa3rUdmm7bOCvOFvqGtPIj59Ljz03bVe/1jJciXZVB1uwRQLAE3nNG4pueIobT4S
Y9xcDby/+h4rvesRxnMrn4OlhJtz6FthE/ksUiXHND8b8EG51pfs4CBQ5lzWAqOQGxXT9RBLGTCq
2aajZ8NhMt9iWstWVRZ+cD9E6gqERq7U3blnWurtT8ojUmoqWMFvJAAl+TCsysQjwT4qrJKBCZ2H
kGnxCeMA0Yb2LLBjSAgFLerqkdtmywqiVVV+IHLsV1XaKUUbGppNtc5xvkRpY47kyi/TkiT8rLoL
tTu587z9FVfwJKXb0jp0uve/+IwJHe1h4ZoJFxTRFChRRaZCESFWYsJXRJe/u6vjJBr3iPnTX3zR
IyRNIhoVxcTjCIoB9umjm4IcjoM3QoBS2IH7Csggo1ohGGRAN2FtCqZAyOSiHLWrtd9Uj7whYBVN
u2sEAOnshzn6oKa2HcrSEp5VrnQfpeucw5RdgImkHiSvwecHWIkOp4E9c55qoQWo4ilCpAIDEL9x
XK0KBnmv7rfnkO154jKdph7j0BZR7whBdR2Kh+WNYIl0vbapwTryU568WuIgfXHtLXnEjmJG8HU5
/qFmm/PUaAAXMkoynb2RXwhi0qSlapw5H6jgkErESPFkk7FBjila71H1B5y3ndruLg453sm5ISqx
uYI3/o4qFYpw/O5m02nZpTrffKWEjgfN+jsDtDHeln+kImX3T7naBKUFARusV/FbxqApan7+BU+q
d5uTxGOhmSRv+kEEQST7cVVgbCgtp0dE/+W7gYk6JIPzr8I2TYGitjbSUbQXhQEU3+pZrhWzCwwg
FttzE3mK1JyG8w9GfN/69KwS4yqQp2PuzDRXSmDEvwS8gyO1jiSdDGXOp2iX1DHCNMgSje5mhsm3
r0/IRKIGpSyxm0+6atSxstosYP6XSAeQ65DuDF3z0+BMfm8Docsjc8AVYqlrLdkPYswcXcGSFL/r
Zu8s2XQ/sFrW2pP342bI+zODyeO/enqnkd4/yv17/O4o2+17AoyV/PiRZnXG+oMRFHyzU15Q6PuM
yRwLz1Rc+KHBp7QaOqzpG4w948gBngetPMdhuET0US1szLnNFpzCNVzs+gIwXcTnKtj2WDvqHj64
jDRQwmnKGQt2NUmee9ptwyw/S3UXnoqP3XEltRWqHs05xTZ6RBB6WUP/lqmqfBhmFCMdgIAofHc3
G0ckRM2CfzPK6jPqJ/YxtCpnYb1PLx4yl8XFyAaiDggctarDD3KvyaOFdtWN6Br91/ADy34YqKI9
ESXaYBubV9nzQf2HgRWxLdjYKb50m+kHsjqBAenlqkcj5Wlyk6ipG7Y5xhqH75wWMMY+8rG7xixL
ienrh3ukE5g8AFQUeGWKGHHN+S3Mx2rwgh+fPrF29gORNICp5bozpM84RVdBMWIqaEugIF1udn27
JGokQdavw6DnTJ4H7v3KPPZ7JArotWxN0fXkkKrdW/6RiKn4lxIxp0DWiRKJ2R/iZTI3EmtsLyBk
jnVq9jhFUDw5Y+zI6mU5sjEx8BeQ84jVvzh7dqJAZrKdPsqzRbfZaxWkO2zOue8iUfajn4/e2Q3y
6TWAZhmic1cAvb3bULZpc7gAODEwMxH76uIj8+ChaVEOwBu13dt1+vNdreIs0ewL190s5ZL8FY5N
FNhSoIAZ/4eG2XO2VU2VkhMcEbfB2itNWxj28gZ5tgTJYYuvSfMmZHa6z+KxWN3TOFxRqFxSD8fs
QYtIvrIlxNL4ao9A0KxoBbzoH0FmDajMkRoeV8+kIwsQQJr1ZNeih9VLyj3fZz7DlUpI++GKu/2H
J4K0udHa5kWokqPhyfVGtAkJyDRy6Za3uBXYyWQAcvte9ONBkw8yq6pguhFInIwkJelGPvFgrhRC
YItwAdfDzUYmvG5Kq9lPfm1FOxiZIoNMumDq/0B8Eu+0TcuiHCN5g8JK7ddmtq6xKVeqdT0j0RCw
JSgjUIKLxo4axvWMt4vKsL1OcOCaJ6CAkSI1eY+Da0WWr4CqRXUHPCfR7H1TC539xP1aj2D7SCSC
keGLYrvZE1CZhjZ2rZ7ExuwFLFpdTlKXEdaigDwnHa8WiXJvMXfdASyK1qywl/Kwpc171DTrmFkz
pPsiE6ervB8zOA9r52Du3rWvxo5z+RX5JDNz+LYCFDvcPtVLYt0SjPGn88HvLD5Ussh77fjZ0IlO
VwOesu0c4qRtJXxxYd7THHp6nK4R5qHaLzq2dyqW85dIS+zcpZRz/s9Qf9MbZ1PzgDYAJMbjrTBg
y4KPftNq6TliuKvl8ObHIV3bKz8E/WCgWMZFX4BwI4XFQ7O2n9o5x/eWaSlddppSsL5ONwOvomdK
9o69S0GbKl3wPEbwaY7fZutXlSsrJQ5b4e35Mt6HT+/YldmC1A0vgOcHqv5h7T/cxBx5fgsG4OIH
y1BRPOS26Jxz/Oa5g2HKkwU95lpmeCd/MxPJd3buFwckbKomXlxtHOGkGT8Td80I/klg8Csb3IvH
pWvrwKI9+37tv3QW2f3PRw3SBr+WdXOynEAdAwiJqmRBphUiMLcTSca4Fja5jt9Tjh9n5ns4FE4y
dYIyauiv13/bkwSvniRaJFmp6eTbo1sP2/C5QxUcuSiLxJAnTNIT6dvlgg8/q/LUdnJSHNUmgQW7
nbSHjNvxkwmKm3HygKZ6iYUSwKH327zgqpozg007XcRrwxGpebE3BgVwLNgC9t+/eXkH+n0xrqz5
3kyJ8eqNaRPG1ph8yYestev+sEj19g+s5HUq/M5pTUpaM+bYMA2OBsfdHbLmFhnC7nYhqT7niIY1
ZAetRYoIfeF/ohtNSdgX6Why5LETt9VMde7PZzmhz1oRNLgZ5+y5hD9haIR9ZpHJGVrcnIRyySvb
rETe9m4EnHH9fV32TEjbwCb+ue6gvUg2JnzlL74gQ3nRZel6s0ijhdCzqrmE22E8KzH6ErJhpKaG
9usfcAEs078YrgUJ79cA8CcVdV6ao6vY7OVe0iM7puW48GChP4kBWC1GzqD73BqEQW+dqHr6dzY9
wjRzJUrtvJVMMsuhrfO48ZxyEMgQMlLz7NcsD2OdcdiI2XKvlCdP41L6wBmvKuujM7H9I3OLiv/F
Ds+y5mZjP4h8UFmGCeKI5SDyUXQB7BYL2Nl+3pr/oiV92R4Cj8/WU0ggY0NuFE+96Jb7f9h5Eu3/
yrMQp5s75zBu7voohstvp7aUEB+08qvJHTiwX99QVTGx2i8aG3DkVXubhUmN018Uh4oD7/45Q+VL
JTQzPXj5fDm9o2rdO+b3m4hYNufwmrKtAARCHKWhyAfUa7bmQSm4tEqTxVFnyc5cqxwo8GTnK7QP
aaXMwbJAxBLbU6iBSIk0OckzUpB12rlQ7QPaH5f0Vn/Ntt0XB9+PYZOUlMp871jWafTcWaiGGB2p
2X1dypA2vH0Q9MNy8fofolGXJSrdmLdNRMifUph8cxRjDSxuE0Z6RmKfWQ0Er9oFOUo2c6clax2s
I6AEjBj2Ctli4jUd0h92JnSnTe4+5qwgHQ5uBx4BJMRsHQgx9vDUDKzZjPAsPtYCv78+Kb6oOCYJ
g5s0C1UgK7e1a3Y6yLFJmp3A0skMo2nkZKL5TfKO3bHWPy9R+1W9d58fhIDKuCio3r8ZPIXLqfNa
Z48iwCPd/NJtoOkOaKlFqtmSgTkkneads5aRN8xpErIpjyFOoEuHavBH3zXi2zh5yGoTYX6kB2EH
7EX5iIKEiNaryfKmcQyTUwBtQZ7/IL1JF4PoiQexPZaWJwwKjysCa5dCxteLSuZt8JZmSrgMVXTy
qmw4NoBKQC/SofJ5KbCRM5PyZFOaFnzv6Yr2Axc7+IIzelsTWNx6+sgFI5+Fr0IM9aMTD7h9Y/pe
pgqfdY8asY9pavzKe/AqPb4HFR3ar5ZGjU33xNocFW6PEPYuIp6+B3YfhX3YSYBXYYvW4URxXm8V
TdEWJF7VFFP8REDWRnelSNo+rk9BgFKYBt3UyXl7e0t7HDLcN1PlUhQOyetc/DmJbDtSnSteC11f
5JXfEy18YnyyOu6mYWVg35g6N9G7VPLSphFjkHpK/DS51bnkmgO5EEro79oTq3TA6iNdbxADRp9z
GFHfEnSh+B3DChHFdN03t7jNlAERcXqQo/Qvk1fdgV8d+WSiVlXJQj4G7F8+8wGiKDuKsC/qVyVr
+0Zdx6mWCNI7/HZNyZRWlI6tv/QlGtfc477om5HKaQ+XzbXmoSIE2oQ0dqt05h1wzPXzk2DHBF01
jVjB8UTJAyjwnRfTTDYOAXY80kWY52BngvLUqkDfsH8kbdqodn4UmeeOEgKHd0tdcJIiA+32iNzd
LtViTOGpKh3mAGBwSajnGMjYD+NhwCTVy34/urvSY5wFud19RYf8I1fKbIsC5ARbIcu9oMZL0HEY
C3QZZ/xi9JJZpjaU0KRWA9u38J7MIhUJEYGgI9Lvee3yQxIhVoUvUxCJRO1br02sxA5YvPwNdziC
m8XQt1LkEd0/r+lijomOtl93+3ozHF/iAVwhzfD/6XWgynsQBgYOFMGGDfuuhG8dqHvJYVwdYzbx
1r0puozAc1dI/5+dDt5//Ku3iO7GNS22i3KOfYvs4UTQNJBsLSHdnEANY/cMF+KmBiYpsUdmIbn/
Ci5ha9rsQyDRuhJIvN/pa66CZxr8nFbJ6JfwS2wy8LaLrbIlQkT753B80bjulBmd2WJ41ULFaWzv
JNe5aFVwNj6FDU/ZAKxophJUNL8IfsBBskcOVvq4nA/ptCifGy/7KCZLviAmoW/VtDYBPVizyAGi
BEKLVfxyUi3s8NbakkjCuTjDaIAkvhIBP0jt3znNtWmOOrHTvp0jB2No0qSAlPMPCt4ssd9MkFrl
yCyHpZq93czBhT+EBHizP3ZVIe6pBm0T3WZ6BkPD3OU+1qv06dQbnQs8VMWexILKGSiPbRqYTcmq
qj8bXFYTIwgWNiibRUkmvlVfpx9i0IYWtZLT15hkv6jieANTotQvrQi3HKvbBjZ7wIwGHO96R4wT
uqzqDwN+lobaXe2PJgmROAuGB8h9kRF+B9WlviyxlImPucs/UvO780A05+HUwp+weYXVNmlXj+Mz
zRwSr1Yw7K4dhWSm5xiXH6uQ9wDLLP2kZjsPxjco66F0ZrMW/CGi7OBcMyB2ORb/QBUVUJjekRfX
zIZJdCIgdc62Pdy4h1kS15gvxdjgDVAOLBNVoV8P2WHI1fqh8CdCJMdn5gd6syL9seW1yYXOxFEn
B+qIy1KvOzUjlFIjADKQvc1/azO8kp19JUzeMcJqe7+NgGkPWpOgWtGYxpMXId0ih3/ip6U8gSeZ
HWX171oo5r7vRCKZKh6IDOMDDefxE3z53NyhfdOBU2WWP6mzez+wgOrJv4jCGN7FGfxypvgV8YGa
7sCFf/cdVkDoanvvHySZG8+QEqKZKUGDTwsgz0d5HdlrsTza53k+jm3RJMps5hOSPo1oGwj0V6iu
48nl4h9c0KfwDoiPoLkNFImaa2dTFqqTExl/qgBNZMQogV2MuoatG2gAZ56XXbUAj+xe7A+a5ZkZ
EXgqCtpjbRFvK5tuwLpk4K/uGvei3sSjjmWkdFLI1xn+34Yk1SxjfKnQLoOPk06lmPX9c7Mpb8W2
Brjv8uymvDUce4hnmckfZLlLdn2gAtODW+z1yrgFR8nbGUguDGrf+fki7cvCCes5aGoMKidA710Q
ekTVwNeooUmI5NuDk9+55MydLQ+CVIEwivTSoLD4EH6AUY+aIunFE+mfVFSizHHyNclOcvKGmJoC
WNlfiIp3vBfkkCzn1pTzkhYV1C/ZuzCoVxt2U2SydoPjmtJaikUbt87iNLffW0yJdP+jz9x2wrhE
wN4XGgbxvbVJW7N5iny9TKL3winizgBjY9fA746dZn0N6/crkv8PzXIYrzoI3wl6+LlxscZqD/fL
NcGxcEWu1dn9OkLvV0sUKj07EDEhydT9Sqk/5bHUHmY/5JQOq9ba788VNgXf7WbKyHC61gdVd7QK
/V5gZ48KCaRFMAyT0G+FUAoItiPCGdcJFCL5h/KCo7obhI1M5V7aWhnC5gIitO0+fl27mz1h4QuY
OTYhT9KCKkFmnT+S/1AcjljE7fkW9U/A+Ef7Zzw7PZFTxMFoNQoxPem+KzjQspwnneBpAP8htY2o
9e9qdYW0g0cYDNzznvdRvvSXYjdLWJdGRUouhhyUJblukypsoJ37ptfoblYzF0Rytb7bs4SQBGr4
N+HqElDsetq4j2rbfH2UEPOzxBuVp+Y7/NXE6zkCwPY+nPRGXEEGJcftvOYKUhJqX4XGWlAHnB9J
vazhAPgnD6oETNe6x5s8lTYclpPlRPM5hD8zgD0N94dUEwx/PeF4w8Oo10OEtEWUd8a8Mk0TOx+Y
E4HAOR8L+ivdIxYiAtL4cZE9PZf3foADRi6p41ymPMk94KLrhZ6q2gfDKqob0T70ojOJbnqrpnu+
Uz7mxEzjqgI1aDfPJ5UIE8wwJhO3HAr1ymiL+TOcksOapOFPfLVNly4IfRiAhvoPjjj8kMzxg9KS
sZ2adUQRTVOg4foTPFEPEawlzPj/xnmKz17lD2LDKxjN9RmGnRGTfNVOyfYwV94KPed6hPceS28W
4ZGIcSLAwOdhqjRYfFsPPjSofxwwRLiw8VD+2iMRazoaoEoeC2poWKhw0ssdGtXenWWaaRXmDX/B
PI5NLDEuUsv5eRul92VyM/cjCUqaXhATqwtJ7Qwz6NwvgsGHtqjMtp9WNxc2PYM2jFKBi9Fl0qMA
XNSHfynrlYodS1TSkIM2w5om1muFlD/aPiFlgJhWCHHNxiIhyqZGQXH2n8lPbDbJEFK88jDxc1u0
dpJutA/aCC1YjjGWzUFMdpDrZbDsWy0keqtuM6oXXJmaj0kpdHAT6WY1QLBkJ8Agfc8qpBEH6k2h
yO2NLs+qCpxfePG+7/OYT/7E1aikKviP+UvC+4q0cYv9/XoowR6g4btVZ1U4lNB8kHFoq9ALF0ju
aWGd1XTGK7RNWrWhjQR0kA8do+dp6g5DtdqWV6koZwe/eykEyd4UT172dpzFbsfYkLjViDfWV+hH
1IzbRWLjle0H8F4xsnPkeD2P7CcyPK1DT2zAMvGFXkmKnXiHTVcvdVXWmDI0QEIy6tWL7CvqkXZA
0saOJJ1GK9w1oHaGMN+rTsMMNEBztXcafi1rvzrRYkXLMhgfKmtYWuxTY/UOe9Zsz0kkuOfKmRDO
N1CxMvgf3SeZeOyCj3KrQdFHlDzYsXS41A0RvUTjtHNfUFMB0IS1siRsDCprXKTOTdFs/c7qI2Eh
8pYdCDSSF3uHo4qKmRSO9vBPIb9/L8vK5Kk3qsSHmtJZTVs76OTFhDlayAtvAcFspssGPRKoL0be
OpViafXAlNN4HOnxEbClfsGoD0f7LpkQoHTmYZq3f4U3Ze+TF04Ec+uE0x5nm+alXT9JV0Y/cW7l
OnWbO2OuJBHYRTzbtx0a25yybSC9Kvh+T9NiUZj9Xco34Zv890ZGD3EA1tU2K2hfmBIeKp3qFzg8
9xL6J2t+2pR00SwgJYWlQri62mrUkHgkw3QgbpP02cQTHZWCzbgHxBeDCUmK33Xah6jZ2bxNbL1a
m7NWFOGkxyde+nrTxKFgfR1OplhiRfys/bkgTT8L+ob6INXccoM+cWZxf+ntVQmXf9g5HG+RTvd/
QTLJxoSQLd+fEDoC1gzs+5b5EB4s6YjprpZHuzXXm0a2ef9VY1haBOIocYgRD5LGPH5yfjfQSUK2
SdK9jvYWDyAr3Ksz/pZtaLQoEIg2CFiaP0Wh1DrmczhR6VGpd+y45QYHJ2SgVH2v2w3p8hMPirJY
jtKiC8vbkFtC3rLdU3TTt5rHNrOyURZ56eVivqCialfo4lu4vNyOQhplLPgKI5KppptfCs6rDFmN
C2kynpV/n6iquV36GH9cZXIrKOhhnzX/rfYAdxSK2uAZypa60iLqLqncMPNaT69GRfBtMWLMUiKU
taolhs+Jqybs2AxLxJlmHHJD/kc3PYy+XI9LfZCH4Z94nuW8l4flBeL8sAOpZKu2RVOooCzj9RWk
/F9nZAqJ1gQ/f1u6UGoIutFoAskfyw92nrwqAZoJkigCpz5YEemNpOZvkqYe9sAunJ6dadd+9CgC
QOb12s+E1ju8dK8jPLslvwC/UpxzJVQzsxijBkxjZ67i3Kgjib++KWbOh1XRRkbYfvY14E3ISiUi
SCypkXDFuwHb54DwHGA4OChFacQmoAIxD62FnaNlanUolhMl6nHTz4aynyrr7TXgBj6/K9jS27f9
7Cuxid2LtBPtFYwkZX/TGXP1viPoUYuy95At1WmtwNA1Zh+1g5J3S6uvIUi8bCSQWJGejtugrIHy
5CpzLOQ2ZzuRjpfAkfAG4PXNvYQTlmGohIG5uriBByIqAcf7ETPsOgDqGJz9krEN9KTc5x6g9ceq
lKRWCjXJ/IPPXNYwcxcg9KMbfXAtOJJxvUGrBIfQgE/rYDLACF7Yze0YApJSkiCqc5cKJ7rZYExR
6IOVgkFQjr/YUA5cpGkTn0JPfjWygtPOHz3eSqbZqFGA59bwt3bjxbTh0dT2s/nJMvMphVCMmnac
IpnT7ilRJICnemSw98ghqLez3a5xm+MjK3CVP2UH0Q9M2knUg/ZD1fgE3y4fwXek6CvFs2qmav8c
NleZTPLy5gqhO6Bc2cgUwoFhMYfIT2wbe+rtdbrvV0/se3KVJ8GT/NOVKRVC4+cxgbSqAakd/4K/
o0knh79Czei1MQpmmNH5Kf6za50A4YVQSKiakRZONjGD6EMLQr7gnsMs1EEQ6WyWfZQbx7/gUma0
4ly4Z8ipVgCd11NBnYUCXs8kct7xoh2mGXCv/xh1wfe+wvjGxDqRtx3Q8XfpWMhUFaiEXfRHZrup
I/YrlkIYSW2yXDlBrFnN7CiP8Od2Ow83B8hMTaQAGoFgna410qBMJ+iDVu7tgnPNI5kSuw+pgFSh
ZkACHgXJD2V6e0kXe5ob81QY4lqJYhBR5GlHUNm/pTFtu0EHH5wpTF1d7eRfRQRuFxv+bIDnPavx
qQqipwMWVJwiOE15S45497a1y3Biaak/GnwIf49hEw3aR0U6MUNWk6xAlDM7SgPfkAEDUk7EIrD6
kYQQaiT4VjfCVgjWdFjzAz5liuFmONUTY2SLbLUAiAsNfES0NAhauvK7LbAuXtQ92Q+01CEzgvKb
14gR4ERP/Iw32+bTfkFH3B8X04VuI/5zunny9I9K2CMDnqjM1nnaikGukQsphZMcPV8GXkBHzs7D
+tp1YJ1AEZkiSm7mTB93m9tmuKvdZ6UYtZqmwnOqE8TGShgdMK4Vap1qa38CEUMmgS/IFnZRXOxX
FlTSZsrn9Dqm9uhh+SKGWqnHV+ZyucPoY23VZRqBl7+k1nj6rH5TBBHzZ0RCKoguU31jWHRQOmfZ
UeSCj/+d/R2tyIBg3nj3VRHuon47uAs/pYLuJeU8nb21XmoRQ95PAT/PMDNoqdpciNLI3otw7kDL
O0R3jA+JJBA9R/XCzzVlnwTmYpj+nW6PP4YJOoOw5x3nFilBO4ME1XUSMgHZTveGbQ5VeFCa5K2D
mcygq19Syg2hSzJ241xYkkdHu/D5mlKxHLUB+d2kybaw6CcUouEndXuLAD68jtGtf8Tr5c6aQN3U
3xnHnBMm9xBwqydQY8JdaKBZVetsuo9dzdVRoIqEfS1/I1RWDuL+4vP1G0y3vqLnEgjQ5gIkHCgP
BRSQEgV2Gw5iDYK1jA/8HuelM0cb+vY76hfZcBK0y9CKsyWLShn3YfQoxsMpKyG1XLmQBtIKzALy
su++vBGk+fOIt73aeDBN8OzL6GisQA0QBh5mRLVwn3FHrxUxwXU2D49j1RILhzfsc/UBKBSMuOVM
4w1y+nPhDtFYHna23pMtWbGwwT3mAXA7JfBdFpIxZfD2Nnbo4+XnGE9kysapgOow4iHeDs9PHV62
n//J6qHON2RWi9Sjq2L2BxOdZB2mQgNlpE+oroldIzifSKbw4C2NhP4uN35H5LY6abmdXJSOCars
5lDG94mtOjMins0guXEprr8CzYSF8W33tXJkKaMo9tqtdO/u5J86xkeOCUutyVDEEumH3XA/2mL2
jr+2104Ufm8MH1Nk1w4TCheQnt8Zv2ODmCbgydhV8mQFMQUOjh5oGf01Vy87eYeNIX7cc7nIVnCo
fUqoqNUZdihM1V43d7nmPn1bXKAK0O66J6wdXojH1EXdrTBnp948Ld35R7cYoWe5QA7PMiAznB+x
pb6vd72AhIWz4MguhcI5zR6uvPTb50tJbpg1CXmfG4sr6FJ23QqQzAXEICwlzjSTo4LplZ4tq4mE
5fX+qdi+FaBxIVZ6YGe3tElfuCNSSOYxhKCekssHLQFFmNSpF5L6s3yNDpIDdelJcE2A4PC3mGKe
jsGHlgKNVFAIr6Ece1GGLeOCOPfgpGwld9H78C9Ws1PhvyDtwhUrCfS6Iln9WFILpQDYfpT+Mpxw
ysq6JZLZvfhY7Vg1ERXPnuk8C/4sBt7plzLUN0qYYySdR+iFhQ/RkgFZG9H9oANkCnCILBVF52fv
xGXkAoPRZfMCnpW66I2NPuBF64EPrL+aXDzOiBRFaBpjocp6t72lARiDqIS4fT6Z5fYXITb9niAe
4z1jhLvBo5SxSOiTQ8VlV5zZwK/02uOhdJzzk6BzRemhDxJ/zpyHkyRy3rG/KE3LOTtPEBIdxBL/
ngrjqcZFq7XL9yTINfJlYOHW8ZfLJjIJRC9sf9mCWbyqx0N4aX1yvaj8Yusid+ZxH1MMQYuQHirT
Ak0bmo2sH12EqQf24Khe7bx5bdm0He3l9b8I7ILiGdjx+YWd2ieHtfDrtTBEP8JltKybrgWRPJ5r
bUdvRSWCLuNbLLZa0BRiGB44rdR6q5VvbXUif8fYCFsPGPKWSNgANabBohIKZcjy5+2W625b7E2g
XmHva4ZvhpPdxpJ6JMp5LW4rzFuNLcYqRmd4x6LT9RMso9d9ImDLHWoxhYN0R7uz4Xd8KQ850DGW
WyF8aEgWD/2IXWbzEe4fpbdzGI0ksuV1+EgeSbfCzK+jebzus/MyYHVBYPh7bgKmy0IDkDp9vUds
D2umk7EaQhmbfHi4BzIkVIP0jlgN1BSJFiLR0oHnuy5WhNtmtjYlYHH7jKfW5fJgrmXwTwdFGmCa
TVsa7jCzkplzSxBl9zAgXhc2WRBvbi6tOG9yW3La8m3oZVrK1MxvoQHvxLHSrOpuogdaOkhhNRRm
VdGJe9/A3oU442lt9rMsruHgt0z6vqF/ioyZYLee32QjSmjj/23UMArrC9TggkMWvAAHg5vOhcxL
BSMtpgmQnPn+CMD1eSUeaEZlLaq6au9SqYv5asTfhUY0Tq0JVlP+ZN7rEWyyLfIYVyjKmV9vsxHr
ASfu+zOCCYybY2QQfxfqf/bxzLXXn6VHpiZppioP3ZjOmlQwG5L366C6hSGa66JO+ovq1KfxhW/N
ItD/69NzKNnCXN+H3zskqVz/Dp+T8wigNjaic+b57IMQgUkmhZnUGesGbAqiUMtEPG+lgJTyc1AV
HwkGVtqAF646JBNlg7CjbgYy4dopRPsP1PVxxoaM3t/wg1sUcCchk85NRFDs6t5zEz8WxYC1fhXe
sAwUAuQXOTWF6fvY3spbj/hDV+Ql3bvJRHsaZzBVvYGs/YnZ3RjYt511BIW0vbCLm92QoaKXoBBl
ETTJowvggzgFyTZQxjVm0wI8q36bLbQImZ61OZNG7dSZYjCvWDXxZ2sPnXXhqLTlBcMwIANNjH1B
zeve+OaiHhhS24h9cp3YCzC1OXfGrCmOiCDFEW9S7s1J7aMXxikSh3scvxqtnIJgj7yJz+U1LLrY
kJ68jHpfBgXQ2WPvATXegm1Qaqq7DAm/mRnkDAql6d4U7LXRWaOrc5PLZrX63VH1NGms7CMZgriW
8i5fTHgthBiOkc3nOZPL6BMapy4jMN3IWz2owGlnlENagDlm3o/JLCIwoKOaECtUe2TnAlmSsFWo
EYoTIA2+CMup4gQSGV13sFR3cGKExLe7ySuUoL5OMReuCgtpeQ/Kg5HxRIKmKO7RwchDVikdrIn2
LjaAoPgPlMbcVGajgmYXH1YERD3QlBIQpPejmmT/kNICWQTYHpSDfX/7jAqOcJ5IvwYfNj/R6hyx
r66TrwS1mvxIDwAnOH+/Pmo9AkW83ixnlCN0QoEcLD05nPzm1W+dzY5mAZVdCtXtrnd32hjlZ8jz
lQNq+gALhNqcLxtPQs9b1hQuSZS7bI1wnZySoZ1ZFEJzeGgUtGxzguwIFg50SE+BXyTgtK0163ad
vXayzuOYEqXUgJttaeHb1VZA9Aq3dthAdFNAs10wpsX3qUFdmpTedbBfl/sCwz5z367XYI1DtcmV
Rlmh3pJpjUv5sfDmgpKX3Ho6aYCdt9FJ3V4roRz2fGKEI0BiQW+WF6m26HaCLXRug/Xveb56WY7M
LDb3UNl0rCPsQXTeP4ZX9YEX4DV8mfhpgqTNrUQAKwkr1dvNKkKAM0rgdYa/Mg1uZR/Y8dAN4zaw
kisiXwVoklsPzoFndEyIoFaRQPrZzvhRiqFJcDzggryxQc/hPmzhDp+D/UGrYQKdvudjhSjrNKx9
zxBOWfbz+nu5ojpheDQChDUBbOFSMObeEEAwgJf0KYWL8J6LrB/qquStkz0oNG2q9mjn+fweeo2N
qSjXd4QlTkVFpDYG01k4JUcn6vrqKQ2iAMxy4lh5uljQJ+j8/oeoj67/B1GJNUGEGRhFYKBdSH/E
jAR43hqI9WWs8ph25G7QyUnFO48ufWOdJlSGpJudmc8fbdziLlcZKo6RY5wSrrYyr8WuRzFtiitI
oyCfvqDg04/0MvMPHk0+dknDCSTTRuRHEKyCr1I8JHZPJLRFfgLF3rAvVw+pBI5QNeYZIR5meSQr
zeKRiJODbE/DyE4IPW71xgqPclUwjIf4yg7Usiu47cnxUrJwLtAONvZPI4XkkC13I9ZPH3EaaiC4
5SREk07F4z3QHqGjY5Y5bAICMUdUvfDL3X6lBV83dZ3CA7+XYfXnNCFR+8n8e4KNhxUGivE8rg9I
fituP+GOe2BHc0V5aDQ1i3/y4h2jKxQ0hwMo8Zk7u7AWo4BvQtvokOxGVD0uoBkwmATvi1HXt/3Y
X9TocuyfDwZZFhk//n5lZcyWlaDKYYjsKZM+2oh0oQPn8CwxnToYukQj4ZqknXHdeAZt/PwoTEih
3EooRsqKOfB2NJbVaqtEbr2fBq5eHJe9TICbkAyj5iLsomJrbe1vVUafwCWVStTbtbjfWRAMy0W0
vwqgwz0y4kR/C2IZJW+YLhYoZvZDYevHIqz33NqaookUg0O/dPPYNK9IXaUFLb6bFh4kCUm3fI9j
j6YMYBGtqlyk+YQ0c9y4t3KE9J2d4n43KK+tV9tj4xEfTsvY3yjNWjh+Yv0kL2e0mDavby7rUbbd
4Qw+s0xLTDsgLOEOCi051sw2ebxGWDltvKeaLEv65kap76VZVULSuCZaeXU+e4mLduwGuuG4BmDo
KB0AXK1aNmAR9N3DwHn3KXeAkQRuyYpKWV680mVbwyG6rEWdSMXwF5RrcLTBAgnpJUolT9Lfi/ON
7GkuTuBa4Fe5MjhyfZ/nfB7IM+5cU6umrv/YmLhr5+jkJt4VW/PfDNRLMdHQWPHODdpYYKUZHVUG
A5lBCT8tZObWLBkP94c9C9LHxnsL4YPAwvVY9Rzx+BHy9TZNTAUfFxBOOCGMki5yeXbB8Iphc6Rc
eqQSPUsJ0RnDwEYgEAlX7G4n9e7aN9S/ToTI9eBjFPsgwKdVm58sGLxD9g8va2MIkfp1+7nzzH+3
PAzyyxEO5117dr9X0l1cB1UoSsdVetd1CkxsY5Fq+Nhii2aptA7w+hRBHdsyWcLnFMVt+9cHjTAP
EwvvdTmIBgsoebikESlHh8rsOFp73vFVVzRV5opdXGiqcmKGPMyUULhlaK104k6VwY9f8n+Yd5ZP
Zt9A8TaGEd2nMWtMgK+sZDmAGgKEUtdze3xNk7ngrSBEHnILPEVJ5BN1Bbw6ddDa4/KYiCGhruxj
mV9QQLbJMAviO773P6qyqdFp3zpY5rstWlbfr5V8kIN/e2RmCHg4q46/FFL9LZbitN/F2AmFVWd9
eWld7/fbMsoc5CzkGfNLHGgPlXJHFzoa4+w+9/c8ft6yEY34Cpx6rXiSu9mbV/UPSNyNuur72+P4
J9pTA5djuGE2bjd8UWvWKPUp5zdR6i7e5OjLKBgdiejjqz+HBiZM10prugBVHPCYVTPG5A6EGt49
ge2mswuAsn7f9ojgRCRqw93oiHI+hr0IOfRS+7iQzgRJYxQMRSn4+ehQYoN788FyjqCxXOMAtwJY
XZajWjl9+szzFWHnTIv6QKUIM+sQ45DH/yXG74ECiLzKzjQ82O9z14hGrhxzx3nhh8Lbb91TDas0
RZSjAKXV9dLJLEnd3kbyhGuB3+4GOTefQHhT0u9M3tKCHAzK9M+712VtPdnCTy0N1Bl0q4ROpaEM
2vPV6EYLzEtZxBcQ11JYC7+Tyz0lQpxDYdt8MH++1KneyZGrGG8Gj++5CUmGoev73IWKXzWYKKuJ
MQzXAc7lnPmUOz22y7+vNRKVa4RawBhadyvup2hWUDTOcOTkZnsB4rymZYMgv5uEh23YO8UnlwR6
YCj6rxtwK5tfFmv8NW05hoURSRV1HC7gSfFSuCoOQ1f7pwzexuOaAqAZftPrbCrR+avP+Jb+2u6W
oq7zpesV09yAD1PNqNcvn1l+Kq0BxqTFzHRgWVS7HhkOMt1S0WHqXGW7YY9c57A0rEtjydedHvfU
nEJUP4MD+LkEtXlMbK6wvuCg1YQv0Y6AfB45xMRAAzJraKjzvKGqdwW5kw4vjXp+Vjae/xg2/QT1
zjQLqAGYTABwViNp8lXdLczOwFMre9YGChq6mYIf8VCIFKYr2jztDQZTy1Uc+1BvBBmPmW1uMEaW
82DGDedagz+slzg94ZU68NAEl4M1UVFthoCTdPMYj6nG4AOiudpkCB7n+XQQ+d+Anz7vQ05RznIF
VRh+ogP/MYZnPT/rfrAZ5qdakUp2sKdMbdRkzor0uvznw7lrT6ivTCTZmQVmqk9gq8vcSgBrBEKp
KRugdmAF/CTeAhZnd0daSExqKnC3Ko9RY0MoIPliFjcewBLpDK0h2YZ+NgAnwqzgcaFgGrixEuhL
G+tlxABHUTVxFebaaP6pHr6Oe5jJOcXRhQ3g0mCq5JjJpHfWaBrPvY9iWCRjWLQF+9gu8FJQPuaL
oMDfQsNOcLT1x66QIxJf+3wM1uIVnJ2Qmzs3SfkmA5HOIyY7/IwKYK4PeufQDOmfDCwULF0Dm/Xa
p3ggAwBNxDt78gpVHDVP0F86h0c5j/yQ8kNC+qJIaonQ1TUi9FQ6hOxAlDFtQVWq/Ho7FeT/t0xN
kvHg/wcMljVz34aQiql2z7YaaMB35AWOEQJc6oi15VF8J8J6F73rDUV9P1dejoVf9JJWIV2sm9lp
ICKh29ql01PIDP/V06mewVlQMcd/g4WVm+YDLsn0MaPGheFrSuJJOoM84FFAi68N7hZ4uLhyysiE
XTtQCGkGZe2rg8tn3cGy+dHsO6zxtlvRIxNINeuzdRzY5HM2rthIaush6xmLF+R30OSxWdEhLXY3
ZdcMcKPtf/AbEWvkZyIMUR6tpP99h16IRM9Xb1mVX9oOE4K6+noAqDjM3YxdNOUL6EgdEgCfepjq
sibNKv4UtESvTHFiap6hO04hJdjKCmdjvKREa30p7dBRbG+H+2IC9NlTsiZwXlRZvPtdK/lTNzoa
c5kxMSvM5pCKmEAsWFmbQ2SYIYLy0dUcdDmO1Og4VPGzVW96zjErcqJ8LjEurdNnfdePdYvEbPF3
nJT0p9x78znPlClnlPuheoQ5AWEEaiHkKYZRIuV5hmbJghOd0DRovS9KnVFSdRztIC4UWlT7qbBq
E4LSW8anzu76QD6SWj5G3Pp67hTXAjvQ0CvgOoTjKeeYAjSqQcV1ONxY1XzvbFYE+7edeEKuzmTf
1fxkZxGv80TdCnldPoi/cZeuZ5xZQLEHG51nhIQMdBrmaM8jE1B3X/p6ZkXVQzDoSU8/dVFITCXD
LDPY4gECPX7cErauEH+RZeBREv4cFx87epHsaMjjwAz/PpGeFraCUXQMDoh0gRHjFlt2F+3jdu9P
DrTbRxPfHpPvQDAyMSEPJRG9DJwam0kP/1CYPWFcoZVFxauRaQR5JXEbX1Ougip7M7dMf1ti9B/5
5lvePXkAa1tLLgwBrfTRTj90r9nKdNZFIyiqjNfMssAsEmUFuO1wIqy3bhbKNmG9SGVhm491Nqeu
jQg6qiH2E8uD/At3HsDI7gryXzKxfOWbZDyfTR24JQvcCdogotJw2ZOEOyHTGHk77P/UW568INe6
NdKhKMVAQveyo5m/9z6qDnBo5Oetizreg3Qdx/yodXFz9vkmifEqZowDZ0QXSOe1rculQBgE+3O3
qlQYG++ACCki+3Rnsc7p5AFsZcS2dH2KxiULMm5LwFeBxftFEWUMR/sa+7xQ1Iaza7l6N+eE7/NT
SytMub6s1lK/Sr0FQgQtKtqN//T69CSZt4ScsIACnzkJfHf1v3jZUqtLCwbvNFY87VvTmDVukuPM
/edk0zKFtnoPwmCptwP3jG1xoagosJEDysC6AaLNJsQIaIyLPkXOSAOKWnxdyDyPYK2j3LMIOvB1
7cyEEux7kiT/r2IuUdu/wLUUl50stXFBv4Cj6N+ARxn5oU0RxpKZOseccDeNKrkjgqn3m4QNcYFg
NcoDl7vnoYmB/HauLyPZKWawWfViS/JIpPlzSlOGEWeGcXqB/vbpPP89n701deSLgvhKpcVrEqCa
NsYKwJkxvLyr27T0nYiBxO3QWylGyCbgQKXVC8LMumPnkEZPRwkxIR4L7wWellsQ7xHDqkV4Gw+n
U7vHIIHwsw53jn0crV4AnirLbu8rZbicbQDXZrV2mo54lhtCA3c0mcoZkpK0xYh18dWepyqkhVwo
P5WxrzBDWjHOILezFNE8amYAKJpySh5L5sMr0gxtgBj8UXU90m5ar3Nez3YaupFt4ZRp2snX69x0
jFb2OtBZbiDpYL3F1ML63ln4qgMzFBEhI8KTkL3JSXKR/p6Yh1HxtmzRBcjxIGGE53kMril7wu0f
uLc8urLPyvwvWiINmrqTvf2J8VsXSIfhMiwonWbApyNTesFHrX0lXmABdTn7H329AO6Qt8nCs4oT
yfNUiI8XSOxrCpIsQXnmxkPgXGIz2WpGtrqrg4uMbcD4Np9bMon9DVhb+Dd5bG6l0Kkdnbgkr9AM
/6gfRK9xYQENmDM6oVFVy3lStW9hLpL9Cm7hiyVfp98L5H3ZOGcToQ+KkoH34CsoCDGxz3AF9NbB
YZ2J9vb29PXzohv7hOqg29PVtlzEKXV2caw30F7C21szcJ/oYV6RS08dAN658OPonEJcKOd49GGU
6w+KLuPtVtARmNAyum+Ncs8PW2Ir0lhdWTM0kZCAJFSXn9Q/F02vtEGA7NH5ueLdTtkKIpg2dlaD
LONKEsCcDVOzvL4Rt5lTE+5y4bdsDdng2Z55spzkM0p0tJneOkCdqoywirCc+PuNnpjJBX5n8vAb
VBTzMeh2iFvt/PZ3zNWL2SRPJVk0fssq2oWZRMXfr4EepCUSAiwpiH11dz2w6FRlS6WkNQQfOrJp
3DI6zgvfLYCiHvdCe4n2l/zWicClBnDkpVTkoWpOWTYMznaSnRkRULfAgxKqOFocbqrpqJB/oN0k
wX4b2J6JsVPB0EE7YfewgERaFIlc00QovMPCi0Wx8028HHRom+sWZwoqgSWB6F2+3Go4bXVZXPm9
JDtWRX1f3lsHFRtoyhB+1QM1W5IlnhOAWTVTE1nBXWMrnWJE+UwK/W5oIfWJ8lt1BixNS0SRNERO
Qba0TzeQRbKTeTE5M5A7H9wmXVCkcCVv55Gy3mgTfV1PkqrWXYKe40GYVbwG90kX9ZzwWZWLojf+
1KATxFDb9KbPoTEJ9gXBcHULu/0ynnOFOCpHcaUXZ0mLsgtcBtP9mpqnuVfRpiw31xgnOul/1HU8
Q26cJATSOqg4lAquyBRWBZzz78363tb5b3gWFea0DiagV6Ji+aCTglrMoaDY/m2x+IQMx/M4aZh6
mzY7T3yYUf1/F8ceBI+KpM8shUWt/Nuxn+OvqO68EOni1rABFGETvpELOXeKuLB6ZuKmbOubb3rR
BZlZanH6AnRXYtA3Ba4YTz7BaMQ1k87Ra1yoX2skrmZMj7wYkD0XrAfbK7xrpmHxqJOAz+uLCidz
5sQiOciGqHTUzkTvU4X5yxd8mO7Wu5tcoSdW9A7ygZ52QBbR/fVMs0mp18W7hG6a+olh4DSWRSs8
Kbg9pxnpDzm0unqdtm70tY4PzcsD9O54Qjq78fQ7Z1sNDNnzUiTyb2Polctp5LE6ummrZhZxpH/g
2pLZU42SqhloQpXLx8IQreQ8Vzk8SIG4pQ5CbOwyZAiOr1dTETC5/7ASVFI89CuFqbDe5xKOEVvL
tvaPcMYfj7ILEy/t7/ZdEpkG8YwMQEBg8fmqx3SkGDVoE8unn0//C3eazoIsMPzqRtx9P/APfdQi
8ZkliyClwTi9A/V9CMDLIbrxRVDWCJEe1DyWcOzUZP6MFqjpl8dXIqdnnY4kf4Bv1Ijjt8JTiIKW
10+fTtpRM4i+Nw5EhTGCe0ANEKvCA+LV607/JbTjtu1z5251Y9D2AuS3mXjs8SH2fFD8Im7W4Khs
gOx9Nx+Y7gmxyEh0tS9Culd2QHbw+xrcmuF2ZSvBF5veU2rzBbSeLu0UjRNVvUMmxYQ8Fr62SPDA
BeDmnofAC6pZfxPy0Q3/q+PcjM4cEJZrPn9Qyc+8HQKMz5g/APdyYxO/YYPAc2q+azl4r1/WVcIe
ivxbeLkL6XT06foAGKDEmX2E5AzkxKRzyWP1CVn7eHKjAUE4lT5+pKhEqkZzwxBuvQgh337KxltF
oEPdAr1FeP7GiedqFGy2vMxSjCyx9GnwyAsaiXO7Fbuoztft1A2i9LrzYZ1nqrS6eorAD1eNOr+u
oeEwkQK+/HHY4MbazLvgAFd3m4bNR4Uvu6hkK89XrEJnx8pXeU3JjQeNCc4hdtBSJgRSlCq8MXyK
3UZ6zVbWQkGg798EwvP4j77L1jsGSjs8Db7Fojm+E5K6tdNPELosDRmEWX6OwW5CGdTZh4Egp+UT
fHpdCLJ4C5LgNXa9bNs9QOgFkdvh8Yu5MXanKzO+i/9hU2KHW9AGn0OzRCPgXg+GlzDcaGX9MFCY
LMYokzChprJqtDmqqf+PK+2UoEvz9YJI9tOHiqS+ljraexuwSzUDvXqGiUz3xty+AmkDBmN50l4l
4C3lngIFX9NojF4mWlJvknzdRlYKwznUIY6RvrEPB7EOeqXr10LR/SeV/2A+j74MffMmy0cgWPTh
84qUjWqLLmde6VAej/kVvg8F1koYYsw37/NrgPRtD3ppwoeFN7/GyhfYkfQcyYiNYpwXAmrv+b+o
waWNPR4c8it/SN/KAyQUylXC9vh5IQN9AX55HvnWksZf6LV8sRaAdGnRGRPwS0e2Fl10gQOtZvgX
a899RoELq4+LdFCn2kwQvk8vovM1W+RpbnC6MlISB2PjkejowkXPOeq9mHGO7W21vbUykjoW7YZx
xjHEjQ4F/W+ykQp+Af4DCHtNi3VdrnPwsqXjTq1yytyvJkfh05hc+t9ih9p+veD8cQFPCMfU1Epc
HUTznlCKHVbZcOk4lxm6wjHKdEnXl8TCkmGuTw7b7fxBZo40w1R1aK3l5vXkQ5mBffnToHZpZdoI
B1FkSabwdsJ5fjE9+J988xik1juJIqhlUyzvMzXllnMNkdZjjwWwLZa++m0Df1+aXu5/wsS46rLn
3TDO5aj0Yhth3RhAgttN9kYyxCp4KBMrT8TNJX0cO2Kj0GlyMsQr5y0mUPDZHA38kK2Yk5ZiP6dW
3wmfG7ka9fnfHkMbRsc7A5PVfYMF+qaFSlM77JRWift/jPZmqxohxrpOykTbyTIeB1JoHg3JhCpR
+JENn2kL2nKS6uCH8xv1FHY+miJ5hj3OiwsWuVbccawh5mVWtroj1JYb4iwTBbgwGOaL8bhIhcx+
UJ8W8FD4fY7EY+kWn9LMUe6Z3gDf9kBBBG+dYveDVlH8c7bkVpHxaBjLcEjzYGCtIR2KytjcUaCc
9w4jpNwETtAE1DiU452E9wZ6yWEX6H6qiZ2sRLsWQb1XYD6/zXD2uedCUOVZjrBJ8Wwt96VJV2wf
5UiG772b+TmGAuPMz8a3yUAIeuLg7AoTQqgaJKfQ/aCAXNEO0DEYFRuUbm+dK5I6cvIafUl6tPSc
5UU2TGBbzI48YIx9s3YWlzp3ojiMAkoK3mhP/5yNSWCgm2Iii5XjCZWguOGv0B6KZxPG9KBqL08m
YDciFSqTgQmAgkPc72XHGQjkcWgiWqFrHbfDMGPMwSuWsQV1k1L+tWT2FZllG6CbR81wHIYbCqYk
ztApAcJ8LlHazFzeRWStMmseIaVnq+xtr8I4vnghvTvjDl0Jdvwz64/EmjraQEoG5ouxtTePOcFd
J0mG8gAt2lZ5Rf6FolKcp309Vop1hfMEWXfIWFntZMVhLDQJNxTJfCrHNH8by6VJ8741MOcjg7MB
VzkgAnT5OnCvNU231AYi9oD6zPBLw6aq931mDVeK66opZahhLcgdVEnNA7QU/KZE8pdQO1sYSIKX
EOSX2in2bUYbYmubZ50iXpWlpFNowxOVHztwXbuBoSQjyiePBNMgp7sW8JHjXPiRPztewaVY+t9N
XG3hbd0f9lGhQoysQpNR06FjtehjhnEG0mvAHr6bS4uHTz1gWsooTVuPsBa+5fwEKdaR/+Rf+Yd5
2IHYp61KQi8v8CzKR0CS5s22qxOUxrF2elf1hQcY2CXZV/D2p+h5YyBRebbo7Z82FnhAici1WiQd
fRYS7flthkh7R7ZqO58+FomIP/o7m6oJtFBfrY1zQzNuACZZsCLJ1AQpa1Sg4NbleyJwDD7MKJub
RCr9SpSqLlcsLbZrJj8vbRIGxlbZPZrFAAdEdlDHSqpYG0qMZdY/eh8a3pUp6ZOCI4a+NehpLDjD
N+EhSx7JoXDcIlM6YkUA9aZElu0J46lnOGO32VIxL2hX/hEjeOzHCfmh+X7/mnoyo1LmkPJjCxIS
6WL70LwNxmzge+IR+VgPlHaAKfKafz+6OCp68XfuV7eDhb+t280UJym/AdEchTtdUqWeCAv9EEG1
wcsxMQP5za2GytmazmdsYY/STTBxURy9/rad/jGO4YvLTxl3Hv0qFdi6cvUzMn70NDaRFTezZP9I
mP0Xzgc7orr3y1lFuJoB11z/I2uoW6OrlXcNQ12TXrqZmN4YDPmBQBtHUfsXLQucd6eu3dNhdVmj
urytQfrUNZCTFl39GLpDBOekcVeWgyj2U448Hp9NKhK2iACGrZtPgR+F44CWCG9q192BeRsJDWME
trD/zn9/r4H5S3lQZ7QYl121cbtJX606AhvovgIVdGFZoikRd63b8ufZKNlGIEDq4mwKx8GL2jlw
/ovi2jVHyBN4diYFbwZxMxPEAfEyakITWjC8oRMYgboKV4jM6doFR6Ui43M4WLcjqW6bBb/DHv+m
HiVRQdKDWRoDV1McMSZMGyvBigXbB4R53NmZfONoyCaVWCoTXEAKKAx+Sy9yVHhwkr3vZXDVkCK4
T3557UOcWoEm8aHkIk+F4rywA0NxKEJByTtKGOLJZMeYzowx10vA0i2RC8RJ4MkYxXCF/BEiUAyk
oDDtjNSVHRSeEcL7dtmBCHYmsPmxf05tnvDPnomolpnBfF/yzPiyANqveoL2vwkepr8IvTpj/xsF
/VW3UPERecZJB3lcW5ppzUGlHcxo4t4X7iQ1UW0DCSleyhUBkcm78dhbGM88IZwG1PzLPy7pPBEF
1Rxe6eWxh66cv4p6ZXWPJblZUYVd8gl3fegmS5DX40VKH2P3ImFErQjhOzUmZU/kasQ/tQsUDePp
GF8/FUOo7wTHnmIL2oijMaYxgGmG5Ksrfaaml9xjmhMF6fH013++UmbDmSimn1ZLlr4d+Syzvyqr
p1d6MMkBNEfIKbSsQLp/IEkm0sYwHeBhNGMg1IeYb7nK0mfo/o83r7lJ05KLqoVYfoZlaF4WBog1
rzZD6H827OxeQSOvLASA/Mo7JqxJII/sE+gfasSw5RnOHleA36S+mS2V4QOGaUceUerCtRD5hrNV
U497W9WX6AZtNmIdyTDMmxwr4dhgkKjOMEczPl0QjTv9VQCbjo6OrzIV71+dv4KJOC1xAPkaXhk8
7kcu2TC4Qf6aXfIaDz6S9zsD/dwa3xqi1z9T2ll2swWWfzqgd7LVqAO/Ay1O7KEmSX8i2yNCwF3r
vYnPx7yX5NFQiB/6H566vyimP4maBDMLwu28yEw6W3SrrLtU7ndDYZu7u6LQ/ThJNctyZ7CQyDxa
yZ47d2PwLi/zJCRKYa6vDmY9I2VSYovgdNcQO8CHHllYW6m99TfyI5fxWxCZuJz+JvsgXJxLQ/1L
boWLAj1TVNWcXM1pGOlMbBSVMoCb/+RXviCRlWa80OWX45TGMhWBVHbFw4Uc1WJa68AUbu8oXjOK
x/AuUWXvxjTb27wRmIhaoNPHz8qRW2AXb83zUFM8cJygK+f+XQ5TgddbgkDPgyna9UL1d+1Bapl4
9fZ4xl7Q6KMYPAYqADCxT/OyQ9UZZ+M/1h0PjiPaSuESt+ARWc4k2J8+933OjBQmoeAluSgvISAg
AJdD8RryJIwH1hTr0i6QN4+PADYor0nZlSKpjOz8RCfB9P8Oon1xc0qsXU0rWdGtM8VTjv4klWKH
O9veaGIeF0jACC9rinIIryxUhehglu/g9lB967N8TdnVzQ4ykBMY57EnhZj+L42gnT2kDKgrzCX5
bxoOGHA/nRP+riO3Z/SR5fIvCzyBmKWLdsFi09qI6irby8mA+6XSfO5vjDuWLQhgqO9UKexH++k6
0KYDY6zf+/tcsWkjrUfHZ5FL8oFuJOYXMFAuNiBEKnC/1rEItf8/lSE7OZ/vKcr4wKyMCmZXm5KP
eWgTMSRxr9YTA81pkbs1EktFfRBg+AzS5BHrxJz9BYQXRPoyCqpA/X7WwZ8bXhaRLNzcxfd1nOeM
K/NWYf6D8TPU0mubLumSDcRvarGADy99GmOAcG1bmNXt6isg5M4l7lLDZcxHkAu2/Diyb0AJkxdj
Pgt0bNO1vwACFyoxzXtJFb+YasSArmBlqUSaJlde98ArJOQNrPPLWbrjLPHOqiqko1c5+hIR1zn0
pWTOQXKkPbOQYu8F3km8geFNAFz7Y/HoqtkRl527y0g9Hr8oLBwc8HILIdH2qykhVrywWNw+bQSj
zeLI+/Z9fGeu88Z8mb8xEF8cOUWqbZL4/K879JydWVdaarkwqmLBQWOyoveocKM2NQaJJH9wZTvR
59nxeMbq+SQR5ckrSQqQouf9S+ObG+w9q6ixmoefdzttfYJMLWF1DLMRwHgVTBkX8Uiv3B3WFqU2
YfwbJkFfhWzU77kafoPCw67i7dVy6wAG1rf9gzZKiz9oGhrX9qjIeHmhfWrM/cw0PR6F3NLhCbiQ
LD0flrA5560K9TkkzneQwyZn03decPb88RC2jHoUHlKyNSkOo/dJrs++n04GarPaKbaXyVG5ikq1
TCgY8qZhOHqAsLgRiAj6TuZJ9RTmCWYtQyMsfsFsXjVCbq2AwaBaJ4i0kN7I62hjoaPc5xyaXw5O
aXK64qSsqx6HbU5wvVv0tNpl5trPv0MgVGXWMOQzyiSAwm0ghURofMuUbKzR9GzDgDqTm9p13vQF
eqXSxy3W6qkReYMP657Q1t4CFE2a3/SOCzeSpZFlXy57G/6CpOqBy/qagf8VlX+Ogx6hAc7i053/
Ymz/CryxRmAlrJZSMyQ/brRpjqR7NM3o7ohxkHWp0XeHLeRA5GCufvCN9T/5qYz9AamCCkzY7Tev
xql+/phg9GcUTacfFDdN37xmv3ZjnMS+zRI7eazGstRnqPZb+B4Dw7rS2OB11a0Lz/tayjaIAGNM
cbtBtM0/Oih/b1Gz/v6qQ+6rxKSkpUwIYZrEQqIwB3pl519m/sgMapeWLoV1fXTUOhao/TJ01uQ5
Dq4KBjDQLMwF3R4cZtVUwG5p489TqQM18bc85UfhVrrdFh7TjmusTgmWip5GTiSQYx9RmN+a0PU6
IrzKjpaM8ncjsi9c8VNSIHQKUyRXpc+1d1QGxlEJt74r9TLcrgiyBzKd/3m3D8DuLaeZV0FxTDy6
NB1nZ7O8hRgDFkuWmS9qse0Gcmbau7CRRodp++FMjGHtSVf7nEah6y60pxNWfKBg72cX28aMooKD
8YlQqs5Yl6+DO/7xBJRKr/78kB+za8iSWSf5GIyIcDi5lDPPxdD3qof0DJGde/7UPmiWyOmO4+YN
8v1y95Ua0pU6yLg49+CYfKAh9xrix325aV6nbO0IrD91/lJDPIjkcdAHhIk34oYRZwX6CliH3lHR
ryKZZS1zQV/4TU9qffjA17pGOTU1dcB2lMGFX0mZ8Us2pIdcPO4SFkrqdz6IptQx1nqPIqcEXN2E
wXPtI3ECEM7qBe2b10dXH/iRnDa16Xx+ScSHspHY8hMG0kiOTeKZt76x1xTM5nVnA0GyDjQB1B8f
YC/UYmR1WlUFlQDDwlEXu8GaTTwpKIGGGe90yZwy8IlJGWEuqivcDvUJ1XJbRVByYCcvSvJbl9Wq
ltAlrxqDLOcblkXYCnPdZXB9BUi0xSgRGrY2nMX/u1mLMZMImio7NUOBYc/TRQ86hnlHfi2tovZf
F8NoI1AmN3OlIGYY9cC0NaFDgeJz4e4mNU8XqSnKnwPeJfp7sKZMnkS7nzOQ1wYBg+zTMOo9KZ5j
vAIZ7A2C4bXo6c/dLW3pv+UYptNQWIPbggkcW+rkF0rqymweLjM4le4jMKqkUulgh7eXlbt/aWro
7XCers5xFbcw4N+rz/LEsfjgwPdya9l0nN8DEDhBb14SYvj4bnYZFEFeIG3vYyfoc8u4OXadQuH4
Gph4hD+dsnh9V7lU6vhgdYVHUJPxEl/fUg2FnNoNQlsiqpwUz9wCQB/T5uE4X5Zo+N7rH9sVCl8f
qNL9K2khhLAfYoXYFcdKw5fSnJ149NXlVmYLenk8O6U3sFmk8RZcaAudvPEQPt8bw4CR3yuVsS22
ziBaTHNJA1orS2gaGaj73tuE2MTP+lqDdPG5fvQQzfyWVvjqKoMIZpTC2/NYL7uecwqg/9GGIoCr
XNCNdaIgpqFFhHSlxEokQygA3bZ8wb8nt4soHt52Fga/JMZ+7ojw5wO5LJAsRVFc7i4SVKPrgY3k
Y73MTlUY7PB8mvQ80QVXqxImKFICQACua/KNcwt6DS1tkzorZXVZ061HoiRSWteLwZrnOlCKPad2
cSN4bV+LJn8NgAtO0VUoTZU1uE4vKaHJOlZTfqr52pOl6TD7SkeoWOLLQdkFnazmU7oNs+ungUeU
1TWGZksHFhTXOBzfaBgFuJSk/W75o66AmmHv41FI5nvg1FQKUDVlGad3PHaQ9z4tzunDpy1NqiK/
8Zsa8IKHkhF8w2cEViP5GDbcFDXOSoI60l6f70MbEIEAPwMAEAZ2SGCeZoHnLSamptLNFA9GU3BC
qdPYZn/Xan7opYv04J2z391+etTHYHyGepjVqa37Qz0lMXIxjIiTUCSOfD/HYBiNiHtUqg/ZS6D8
8uEY/V4XVeF99p+G8SWJtXyj1Cr+sEsQz/52VAEgWqpltbpmzY77j7nC3kaXfYZkPoYsNt598mr0
tZd/bSrbW7xxoT3HLuPnIh5XMQUlOLMvlvPOwCw3+Jy+2NK2BlfBYkVFeLZp/C1hhKS2UDMitmLY
8jszGbBIMGN9QqZokvZvwp/Ukb3QW+oYB7fk2bxMDbQGm2ByqTrLr0c6+ZSlX9KZYQ1ol4E3EoML
JT91M5cYSXRlyqJ3Ist46i8Ar9mb5e45GR0/IUpGJMh0Mn7Wua4YFvZfq/cEt/99Qk4+c5JD/Ur9
XWTK13DZXtIzaHy1V7ANkNd/nb+vVVA46mEKjqszIj79to59tHIcpAt2xEZ/hS8LoFmDRdAMccNE
J1zkHWSpz4iS+axFA18y/1rl9L9LOnTUDknldBIYUPNzaRfYyDNBZY/p1J9ukow7QIytFmb5jxQd
UP9WqfVhHVAqQYtnj5nqiO2Dk+yoQf4GULzsiP3vU9tT5BxnXmGw4Jdvsz0627V95OwDy9ZvLmVn
W+BeLckt2UBv6GKggWOE5XfrKSUFDjfsHpmV4q13fiLJfISUlYIIVT2GAOh6cg9eaGPrc7JwseGy
Y0+DpIKD2BtbROVSeA+MmyJcZ1b+E9Gw0bXMETmFoQ7UdMWoL5eMJ8OSA2EXuOZHRysQoS1GREto
Bd/s3nPNwDDm5M+DnJ8RNrb2taKq5w3OGgmRYUlqM7gG3lVVAXjiYZUCjuqdp8VtXMTGlmzSSvMY
PNDcUUufPWqtSESOe26YlhcVEhOmJpTPv+A2Xf8lo1P4l2/pYb6T5KM04EKwajC8iPo6H1ciBUFg
+5X53T+VpDF7EqeUTKPmI425DsPUvWpxggXq0ddYM4VBiOLRcO/UwKyeLnrhdw98HB7Go8SWn8XT
m3uZvrj1uPf359El3RlcFXQq16HR29amIq3bWROYT/2JXqXhgOh9h+p6uD2lrJ4PLzSnycgx0rwQ
NB4W1nYok4nRDgCjHfKuiBCjKxnaE5Xp6Fog15FJsj1XVeYluiQcFngfJ3M1PCb8tvZyqadI7wmX
gjXe1HN8oduZvzECSvDNama5HAv2hZDw6ijO/Q7LcnEC1BK+O2QsMTAAKRaulJpGmcTJ04Y15/du
FNMQNpFWrzVv7gScHyhb4VLFyncj805Pswv/UQnAFz990G7g9R8tXsy+/EEekjun+daeanHiNHh/
JokieaVsGHjf9PbAbdVm4jW+Z61RG7Ll41Pymrqlv7JSgeW6ZAhYoIxWlPNPMbdD3PpWGf1zB/sb
HNNYpXhw2evvdRHp65I53oZqOHM7KFzTp64q5Vxe73j+dYPX2vjZDr0yHaGJhfGkCUVVuBd15F0p
XBCXONnfo/bTfKKb24ZVpwwFGrCJLmMqFDW2nf7xWFvwtwormW8mEHcFAdGKpTDFLmTidZMrnSBY
XFgNZ/h6f0DrXSQUVRRSUoFJ+TpbGE1aqEv621ToLEdfip954cO8AQZ18yh5HjDYikOErQOjEY2D
sSWBtzzqhZldgoJTiWDfxPx6QTtTabm0+zoa03cRT9Mh+GS7K1RmF2yXqHo+m/ZY9oi7f23mbW+0
5+B5eMmrLuPfIaEOwm7AhCi3W2ls0LC5lca3TzDAOzr6Lldai0TW68ALJM1Q08DtaTh9A8t2ijKv
6YKP4EkAz3YKKcT3KssOfcdFC0Y+lfTVWJM+8CBJe2OmC/PvCqKf7PDAWmPvIfUCqrGgucIwwizZ
V+ibmQyuLxmSPxfyQCXGxXwcIuTHlf2eWeeLkpkPAD8ITfZsSAGoyfGVQkyApG451Nx5Krh4qAWf
gghY2rCy705WQFT9MCrEZeUbci2J0jmEaLGJwSzWG9WpV7m/vy+inZarq99aIqTsRxKuPcEOMsfi
gxtwAEm7hPQGHc2/6n+Rb3WRZOkbOt3YpeIuT4DJfpf8xLjH4xe/WXr1eO1oeV+XBoTLFrpw/m6M
aGT7pKQ0YLXY/sPPx4eAsFqEdMUSli3g5CCHLhpuaOqwLA986cRlkqSjW/Gr5n/qPTUi2cWdPvN1
mLiv7+DO/1A0H6UlbfHJRgJjLPzXOrkt3btoSwFefZMaYPTadBNzfB9mt3ka9jfgAQYy/cSCpzEk
dvW5IFFVSuQyMUwsd4yzPeff8Fp5sbrLdZZQtmn7KVv4+cGoAN13E/5KGh6/jERSVzKdgfiqQ4+G
yRU0Ragd38j6joq3B/IYVlG67GAQLETlgr0RbvbkHk6bXtdjveqtjfO821krxbjM+nWmsyNi/OkQ
CgMiR72KuFtafif8Abcrodhq/WrG7tHFFGyH9kF38FkwF8Om8bKA3rbAuDpAIKi5gKHFmIspmLam
2jRJZjccEhdYo49luK+TYmHUiWKgOUJyG/VAhFFsX+NF2mP7oenlxhk9Tg2pUbEk4a6n+vBIpM7n
PIuDi8fB1S1M7JgaAGpyHBiYwuUOFs/GbwjFz1Qm0Nm9eTYVXIxh/gA6yGfZlVONWwsEgraREfDG
7Bp7SE7Y3k1sPU0bYaUWyrKFyKZD/eJI7TF2qNrhWZfkH4nkqehZkWQ+41CD/8WmgYc2QQr1DXgS
LwguDqlCy9LuLZn2l8JKM7I2gz4ZLd1VVoWrU0yw4SOGre2iQ8Hqs/mW/cT8zif9LHEYtJGCIHM8
5g456ihHoibJ46s2zROJCXJGeDWBJ5a5q/QohMzUC2B4/roj0rZ9gnGFO+yvdhjz+FeXyyNzmP7D
cre4mvbM3GpNHLrEBuwFQ8Cw6iCAnVluIKJRYVjI+QDVpnvoOeqwn445oRPzFu5FtruFTcj2w6RK
ik79ReZ6BuaMMEfiQDDR/WpQOAgU18anUSZrUTAdVtjD7ToGMgOHF6Yp9CJA0k5Evvx5+HRggZDA
XJb6Om1gZNk3AUw5EexSJPm0Dgig0irU/piLDKDC4HOq5PrY66y0WOUJT9bnX1WZe3jZ06To+16S
Ntqkb+F7Kdmnk0r28NoGWwtl4y9ks5I0SkeC0dPOMkWB0k/fPRR0Gp3QUsksBmFr+4pjT8w9JFcn
zSa0hEgT9yH3PtpaobQqfhD6ZtQiDJXM4TWmBZ5GHyzZPBh9pDvnGFjzPTXIaz1iB8PrzY4BLeIe
IJ8Vsr7o+T31cJVAFTJBjrUAZaf3vSSABFUn5o6UKkxpSGPs3upIcq0sIBjVQObZTTVLCXU2dJIY
Km0auzdi9LDiMbi1FqaAtU66fwM3EZkenq/yLQxte+ZKnFVO0S4cJZAFQsKBf4wp6cKZJj9Or0Pe
7xsyYXpEA5vJIKfvKr8sSiaCIDeUw2NoEWuWoz8aFWM7FQgcrA4Mo1RyN8CoTHeweDBF6+REI34z
0uPBt0qVsb1VUKWyWZfxsDyx4zSH9iPtvFcUYYHgVRyjXbjBHw/aYyE2Y6xaPEWkOHYyZ+1UYwtv
4Rwwklwr5M0GcUC+LFu5yqr6iL1a5x3NBOHju6ZtorrIDuYBZGH3nts+MF6PUmZqD74A6lHgvBtw
FCUgh9fNtCEISHp9c7/H92kA7SsA3Q2Juf0ia/OF0SJP5+3QE0fy74PZyVgKBDVVc4cIPkBE9bru
4RQRMZbgXl/dms5hVa0HSomY1OxecgbV39yjKirdbp2N8f2Sk6VFot08Wjn3xuQHrpEAnhSP6WIv
olnel8oTRt+l7nCgJxSfikSQ1MLie01rjX2+3e6J3b+AGs1c25aqj9EuBxdAeSeaM06i8pTlKdqO
fu5j1BE4yTdEUvjyIG4ZiCW+s5NnczqOdp89xHbVxXQwYHFAOJOjvhnGQgvYwZFnt5ms1ydlGHs7
MNxCF8uu7FKJOxJHKv6TAOu5/Y6H9/5yakveTQ5hzFdsnw8ETDpesDsRXSlwLEDqaxpGo7K7455Y
XKdxUVqqiBCEN5AWWE9Y8rwjtEpJ+jJ8htUXU2wajgi2M3JGMr7RPJnYP7aK+7rThf9ClLhSPL9s
D8/UbHmqyaoALpLdtg2yVORQjD0S40e7VtHM5B8045MxHw3f6UlRRDrNXhiGtzoAAgRaeF6qZayw
eArTOmirWKB4yMPnXAF9+NJ9eskd+2h+Ha3+m/KeajvYYdKx+KG/tzAoQNckGaGOkUr/to243kze
ooeez62IvNZodd+yD0ckOCxicG0oghuRiccCA/HvWwX8LkL6RvJvYtQNFQIwxy90UIUcFbOsx4K4
+rO6i3HeBEJn0IVuczhA0IcqzLs7QHZ0nsXzheDhshTlAsFU3WUV/E1omovp+Y/I+Kd3Nw6sJDHL
Zo7eD6gnA1z1CB6cRKEafOSupsOXGL+Qa7UaEXoKK6wwTrU559LhpfyYBNHv3aKky9C9WeKNL8v+
cVYbPBH0NK3AuCJ5Vq59F06CLQ5KBaE611AF+4nWF2WfflDDq2I5YCXO9C1nxWJ9mDdrqpazTjyG
R3va7WmZYOj/8tAtbarl/k3Vx88CAI14Sx/dtXqiHYfhXikOtJ/d3cy7ot0IW9J4OltxeVgB2EvO
2bZLIbLr8FAZf6BfBpB6YqyI/5o90c54cJ/ZcD6DiilUP67s1GZciRMKB+BFba6pgge4/NLcs9pk
lDbI6elA0FgO+qn/q/hetpLC0GVU6vkVM4aJYn4vGjDJ2enThlgOOpEcyQnIvoKM1jc8UDz34cyw
CzV6ZRYGyG9b+M0O7G58LXmQ/ka8lTeKzgcCAkCkk5KXNEPy5N7Nvx0pPCew0nCRe8kTJ1AZNmWq
MqDALE05wUfOs1geldk8qtBKgg6/lMM3YVfdGB8OeHAUi5LDPSXBHZOudaZjI66mYAOGLnC7qkv2
TO88qsb2NiXP0fTRBpK8v8wPawkMAbMM2UYLUTKtOKSDlHO9wgDlS7sZhdV2f9qhnIvYu7zfvYtd
TE/NxTAHq/MuL03L7JwSaEh8My5E8NcvMNffW0rMpiDrK9gNNXsDmCANTDjhO32FOdOZN5pIlD+U
RdetT+PDVSWVDZ8zRd3f5AYIWya4qWxVwf3N7l+ZoNyxNereNt8yYcjtxWaXmJzWZhVf6hgdnH92
QtMcj/yYQL1ct1RysB6Yp2oH0AqOPVPnK9dlMhpcmVfC3olrSupTDoJJp7cbu4wlFMd/VDB9O0KM
beA+fi4MQnXROUSZHMGlxrLXubOOo0WwJiaULgpzIHqHAsfLCm96HNiNm5fVBRUpAardMeQHHcG2
Yi/gwKRRqPcNx5kB25ZPEirSAbMsvehTGTprP553y64WAyLa/1hEpYExefMkUaZh06Imr8H/kATf
8kMXUJDTYAlqvDJSYZVwfeYPoqJRkaLTwN9lgK8R0psjqX8N0Sfee+2LKqvi3xT8ZKOEynbUuUig
K3iyEydNs/lJHcYosIdcVG2usYwKFVrwEVBJAUmTU9I/q+iNKpJZmxZt0T9IphXP6ck7CCvGGLru
gljiDN1oBoo0YJjqGPydQj2N/3Fwp0ZDkWSTh21OdRra19WrzDW4//qz9iyNzThHMMzumzLhRe6i
ltgnjixgX/Qmkks4IxUwYYi6/TFJ77f1zDdJi+2RLxTCPRQKoGSAKYJry1S3D2B/z2kneWfdxYIP
fsmUY4qLfUBZbh8f+ITgA1ykG64TDZ6gAI/aAUTqV943EVb+nMhNOwclAfnfMlkixLPbqaandZ8r
fs+GHbWscMrZEFaLazmzUwiw1dmXemoCoPwVgvn+k3wGANSLtxyISTH8Yexfjhjdwf0f2K/SzPFM
o/k84SFr7e13jQ+X+FZ0ZBJRoAcpqW96P4wwkXNAmMNFknrar2jy51SuOAeOwINrJ/UdCVD+Hk9N
pp1LOKBFn270an5kQDqV4sycdx4Kb1OqidlDnCp4z2GTCuYfJEItgbSgbiPdfuCuNZT9cbrc600Q
XvW/J+HqTj5oCRrrB6rgy9xf1vUso9cpxXhnOVx6JC+voJWQgIVLTQaM0LVt4F1S4cyJmOxfJF9G
tgQjkjhSQsanGUoIKEaQyhxjxoXs6VwrKnY/H2BFaXnswNmGl5/vK+Z8/4NXN1HFGA2EUnEdMJNm
K4hFFopB39zDAop49dutE0DmuQmBUD9MJ9sUw4OFJeNoVvRHCuze0dHNqqfI2gQrcA0m/R5LtZCt
dgsLoHUTCqWQ0liyOa5RMhKIqTubw4ILQizRVCF3GsYJMp8M7QoHzHTtOSzUsLSEaLNbz7srtgwn
Ut/qencwIbTkay0qKOwdP8kBD60qI4rCwHTunfw8JQhj00vC3DZBjoOAZPF6FR+sA0tBqUy8Ffx5
VgOB1WFuMD5iY2oqIVcKSri/36AfkF28Ek6cZAGCbX0JeFxhSm+P0t3XrUOSPO8rIVHqHsEcpdRR
TG5ON+UcBclUJNmrrbYQWwCVkOowYH6beAMdKAlX8t1W31Wjo8mS8eRjRhqszn2fj6TIzkOgzrWk
uH4SWL7aLoc9QWGSVdlzEy5gIWYY+v0GzPcSj3HAWOvWgQHZ2/5FO8XF/QRLbtrivyOXZp2La0ie
xVHvLV9mE5GG+fAFBs4YOwwyFzpw9NSH044PckvalSUb5F/ghTa+IcWAMhzdXn5E4KZBrlZ6Uba6
RSIpszEnuy1WlcN17kXwGw7fN3KskmNqQUPDXBhaSXs4lOojaV8W9SmljZpGVGGDCiPt1wWrMe3P
YZ3xr+FN8H7hsoF4wjo35z07v25FjbdQJVS6TTGZR19BbBkuMZ/aQ7a7qYs9/u7M6x8wog9HLDa8
P1is5mWla18ETSSFe+yHy4ykUKt80lyt6y0OXfXHSMqxy1CnjQd3Wcg0sQjAS2wIrvj12+wq+XZ4
ReEnGzE2aB5HGE275VmRWdo6zlMGJbaMOYCoGGV709r2VoaYZyTr1hKZgvOD9KZ73qbm7eL4R763
gbuMPgHtYvVlgQeYkMvHtWlFqUu5W+bZvsbRpcudpyAmqNHB2N7X+sZ9MJ+HDozEOVUPNEJRS5gM
/ThrH2/RHPzSb5yedpoAPu3Iwfy0/nvYJffmJNUERVkuU9KJL/9rmcdc4ritvbF4Sq9fmVkY4zSW
5hr4R7DxkGK/w5Nx1FbecouCep0n/xriaN78gHRyhON2b8Z3cc+oF2Lq7Bgt2FE1XgfSvSyCMIaM
9Oqh85GyTlwDBrPKJPJ8QYwRygwP4JRff12LMQfiKGtVML1KWFKOZNhq9ZwlHK1AzRGExqTEhxUU
wUQD6BR7fwOJcR62DE3sKoUji8cXG9Ta6FyOhcytdmuZ34PER9oPJKlV+svbdcFekwYBzFZHnVcc
T1eYmnSUkvGQLBg+VHjX7aeY+rf1m/tlPC19UQKjHxANUlqhvDkOGd9COFVdt7S82fc42KW2YmsT
6Z66pPDa8D4ZpJNdfw2LqlvoP+itq7cgJ+4H0e65UjrQKMzTnC4pH2u6PIZxY13LrH9W6Xbt9Sjk
K7XMPvAYCW5u6pjl38Ji6qvCauDlL9hiW2Mb2Eeb6ZCrG+g+mXwXoICYwLFB9VRhy4gPPViDIlnq
1CCKxdcGHUakU2EJhf2MEUiYfO7dAnsbODvOrajZeqAk0NradW0OemxaqP/i0U/PMVArcyBeNyCT
sadCpx36jJ8P+heTjTTVfgmXZqvXjRxWgrIt+x3NL+lQtWKgbRi6BtsPqTZTLw68HuT438uifzCo
rH8nkmPPrI/WhZM0JoJK1nVu/35lmnFgQQrEE3MTOwSW+s80j+606mf2m2yhQRw6z6/VSRCWBoc5
Z73T84LiJDmBkWaUvlH9b/x+G+jdJNFTTFLKPL5CopNjJt68G1BOZRGFCqBVIQpigo6jNpWXaMvF
rzAlLvjDhOrTx0Webg0QeN8vxxs28+tFQBLKu5F/eZiFSK3d5LNsp2efhXKMThl9YfBh0Ll1kfqD
oCO1f3us7b4jvogWqFmiP5wlp4dNBuoAVWRwHO2bwdTqkbzxt7fGFYSCPhVT4hKwlhy7IOqfEDSO
k2yqwJHiRnrtvI7aHqUQYBGHP8S/T3ArTin7A/7i0zPiutIX/fhEa0VqqwKIuJLP97HVwDEI76UP
pS9GwNpIswkln055Kqj5sQVw4HslfNDi6bMjt/DZq9mwAenX7emQNwED96qG0k9FxF9oNOfuoVde
UKZ2X0iJtrICStn5BkF0S3iv2/2kt8h3hHxhhmjsfz7Lp4dgyNHjbb3eY+S6MhAd2V8oq1Q38Ky9
aGPYK+IJEzNvZkbXWMk8U3pDcgXaSy/Zu0qhhG4B97lAhtr1A7RQKCh9sh1cW041oM3zljAN47WS
965B1qCutDHS/tvhmRc3fa8IyaMShn0jU1DJMAby+H+eSXE1mhtHugvQJOQxFIRmrvlItIRhWCuL
dPxykaWa6lpVsZ7KVwC/faCoirEtIVKJpHoYR/J/qUo1WQoSJCptCBwT0VrG7uQtKS/g3hZ/ex6+
sVOvutlePvn9tCcR7i1UALJR43pDqj5Trw92fY1yzgqYcoShShQl8tXnJ9J4plhtniaCcGiWoLtg
yfdcPA5UP6f7YCtyFP6jwjc3XYEa0ORclVIneI9IRJsjrpIsZp4GD4aYdLxIudFEmo2vbHO+mG7j
t6cluFRdia4CG0LRsiEQnaAT3f7fFryAMbPPFlU7dP5zvLj9VsC4WUFWqdfqJvq92xmDEikpZuNA
S7XSz9JcDLor0M1LLeJnVomFUTTpy2jZKuRWIA4TDBrUflLVAemla4FWvrvE4uhEIELKau+CVnnG
6aNy8X17hGn9jgG9Mzp8x9qBCXkeV28XziZqPQ/wCuNUyoiW5nFJpIVo7FHM7gddv7rQvPrBVlvD
lEDOxCN9cnduNf1SyKOO8D6VNbrPToEcb8Qa9finbYhTgQvWj5dEuG3SvxDiLpZDMynVfUKitK2i
ss7CRvC8i1leI8JElD8R4wtA6IHmlIXkUCJv/Nccj+ex34MPwnqdj72rriQQAX4vwbWOGc0yPvwg
nDEh6zPNQ+olNbG1KKxfp6JFmVw5oceZeiqM/Z06KcJNITHJuDKP28qtbJrjeF9qgQRmGJZN9UjZ
CbuZFuf4ODo/wuHK3oDhHpCm7shocwYMxYz5wDFhSeJ54+FOgoQB19+ecwfX5L36DLF3IhS3mU7M
1LWLXMyhKLII+Qjow8bW01XHVMwH13NAec/jolxXB4pHkRJd3fpwcTFlYEdgtGxRDpK8ZC+angfX
etN/WwGAi1wlSWvherU59qfKGMZb3QpyVMQUO3C/l9bwgxWoCEndpYlk2MBgB/QMBNK9qxLMpkOk
yzcB42X3B5xhwCksw0woSMN/IeATQajwmWadFm2vGLovZIHTI2Z8qwu6stX6RtVAG74YKhJdl5WF
CvlxqNmbGplMKVpeEsxDzp9SB/OAhDOGcemWGaNxHneddaDOnrQNv8VNZk/kMFMf49gT4ShIk4Ym
xZoXLwoyUT3ChxFH/LR/xxlJoRZpM8cEe4U86nSN4VM4f/vaMAunLoatLBTIIad99C2MEfsEwKbc
qCWwPwy2MTPbPLwvtUJTso2N+wtVhWbtb9HY8sPsVaLkdU6Sliny98cwiW+NVyxxDjtjnAcURDQu
mfOD/u9GPCb7aWDi0OqGRN3yrMVIqHnPZXe2mKmRHraXWxFB44HVhaIdQLeHd3BQ+se/dfJhyat6
TqC2OF2auqr7BIg+dXd+NNPCLmlEKe2fOgqOnDU61ogcvRTtxeqFrb2NECEx3+zJRPTlurpDj5iB
zBzcGTSPIJoTlrY4kRJ3FAqNstQtB0x4cJ0TdQwMwbOCQmlYS2rYWb7pGXmcTYjwVKUj21xGuUcX
mJXY9gSIEVAUIQs089a7Mm9AD0C9pzFHjxPMFKpzSQ3+E7oOzWF/LJvMSJLaCqFOYPNUzZLlhWZ1
nFtC3WLXxyf0NyLat3BXAjAy0z9F49/VfXFbWOKAnOGiAC7NuRRgZrWchE7m1u2pFRtF4kxdVfnW
XKobwEN1rksDrj9FrS/DF+U1yrh+I4rvFZRZyRwIf8+5SqTFPxax3CgHeaMsplZ65vQ4Pl2lKHZG
YIuZhr2f6DyKW/SidiKY75nkiFbG/InmoTjVDoznnu8EurGg96FleRWvdtLtnUm2ghKPKfZyo2VT
Y+k9Ag3kMT1+gUHzHLmYCtNygBwJ4eYq91X/NZhG3kMFTsN3nTSRaRXTlFNMfOFbZBz/kp2kupOc
It2pTsCxy/InDxeJauoHGWrJTx0Ta6OAwPDevBQUlToIUq4O7U+YJC85SBqH1/5WTOx25edSN86R
ln8RbcQx18qWlrUwMMOcELjDJ6nLIZ3R2j8BuLOsJ7emTy6ccVD7udGTH5Twmc/bXFgrXznkCiJY
yklJeaSuG9sHxQS9nbNpyN5ZNR10Jnbjlrmwh5m0bfkfnFGpvD6Ou2dHpL2mSHS+u2hcUfqAgT6I
vTG6zwE7PtHfh8TPfo0soAj0/HoBQDVWiUlSQWRJk+Djv2ZP/DYEcIao+/zeu8wcFEbjodiyU5uo
zPPFDrcWdzBavVF8m9R/duUtrJC3CBPFblKEnreWIbl3hMVGyozhYy0uDa2bhnJWyzLsiDMTdex9
AVL9yrrUKZn/Ot00my1cK0SnwgDpyTFa77TkmRIusPpjU8eX1M67HiOQVgQqL+x2hqcI6IrUwT8Z
MBI7FQlrND2XQTNfM07vL6qTgEXNr5mHCdOdvJcscTdexHNfFXGoZeZSfe08d2dQTQR0j6oEF/oK
xZ0OpljAUubBuV+PRd377XPD+ptTL35uHJCCBVaE3624eE+vvDPQnM9KTakv8my50WL9CNDP+nay
++BuHRxUs8L9MD/7e5Y7gOkFf/ogEeAKNX6sYRUBRmDiu8HDtH5Hvd88EdTd46TCONs87FRew2HS
JTzYBega1qdUmwm9RLwW+KKSYCis0PQ2BjQkBbrGqdeYWlgfFqOs9NjKlEpJuGTNUaeq+Qv7uGmV
+Bl9STTqv7HCRNRG2ct8EB8efTdcJf1x+rpieWFbCYR/t+KpcErTmMT6E7Uvg4rrIX55LRdmg5aO
J4HX4UrezzKugMKcUJVEsAqpJ/YKqcbqntCQm3XhFO/nxDRFWZeIXgFhGYo5e7/o1kXESk0FZipC
ub3n8pEpWzepdNkNZnQ8ZspKfJXaxgkbX+Er85TmJH0dW02dNAYA3lRNY221jF0ZJ5Zz5cYqKnbQ
vh4I5sgL7FKYJ8NEKz9pEh45apXTTX+QjpyrE3mNFTaILJRr74a6Suq4lQiUEPffdl4iDAX6kq+u
dHT8p3mrDonGdxQ4bxMRPXGr08aZf4o8QYFR4deRX+zcRENS88CBeMx3s8Ayu/AEiUU3XrPRZ/QL
W5X6EWGQomV5BFjNIiq/B163USlYteylLk2t5faGSyBY3ZOKr3OQkdUwYMI75MEJUte9fc+Jpg6G
Kwrwn9/UC/BbdeISAW8lydI9f5HIR2J1AoB6Edi2Mt2vHr3Xj2i5sSeuwngfHasL0wFJ/1kEejIq
3FA0LhWAttUU7Ap9HVnY0GbvgqOjM3xyYo3wauOwGjS3QARCu8yL6OJhaU1ofKlkpjyV9TwWz0XQ
n8VpcrA05j2zreI7+9X57sKr3HZMmkcpVPI/lRRnx6Aye14M1WihZ4Uf0qTWPVifldmlqNlFWQm0
h+C2ECz3obh2d/louzUyGgdTq6o8ZipLD+pPX7sV2yVMBXDrMBQZK7b9PqSfE480ZbNdOBiC3VrX
Cq9RvzLu/Vz4R2IEKVafU54odCqSBa9ArpHHlvaF/0oiz0rjWIv+FOR9xtjyMcHMp18nkVAFju6J
tiboftkMqJYK3abARjjZSy6WlETBBLtSUhlrJo3CAZ9058y7XlwypZ64Dr6P0nK5fFRINpQHgBKn
q+sb41NWzZHjsgiP1aOOAsVruj2sVdioPeO/3WHnZn4McYAkv9H6Mo6YxMb1Ax0xhC390/H9zUb+
NGhzsW+HURcqlgRMPLCORwnuvwHQviFmz6dUT6ULeOgccwkys6H8BnoxpzaAGZPa89EcH28YKm9Y
H7DNoYc0GP/ATGkxjUni8C6yQXWce5LJjsa3DT/ZNvJLhk8OJGtv0R2GB2N1dkgbpS0cD2YMcjA3
ezqKOxG98GRvo1janNCWsdoJOyZmQEpKagqPhdz1BLiDu8rbLVUt7G7wBQGax0cO/bt1+AuFPesA
7X/VAkELbFZlmx+S76gc2tvTYoahg0xiw5STk0Jf/u7bcqIrdbWUlXBFnPDq2w0Jc3C26U3s+PwS
OmqQTjhri8q/njAmsEtMApf/6TvgfrC97/fIhI1RR0tn7HXbhSd7j/l4K8qbtXA800PQpfBvLq9z
zr4gW0/zcy6CohdeK850OB44GF7adXEIN8NhTffJZcmaBBCWGTadyb+XCNHXWnq5mu3OxZcrAw8a
ZI4xxNnMKYsyFVkqWWfo6Dxf+WnNv8ArI33UkOxrXQhbQ9ME2hjP1jdeTcD46iE2g8QBOok7wR4h
WwdLsJ1H098HnPAWD2j/NWLylhQfK4jn2pA/g7LnSnxQODBvf0RPy77g3JjDeTYJ0LCV1BOKrD39
ptAKjwcXCrJQaA6nffu6BxAKakPGdpMMNle0tDgfOFO7eugDdmzqI/4K4kdzejkNztpbDmtbMUpI
sGqu2WfkB6zlIXqoyyaKFiuAzmDBFvQQQM7FZ+Q6XD6N5P092C124wbolCCkqgPJ82dGBn3NLynp
2HLQunamyxNNJS9CvTQh3XFa0nd+moPqK/WDthn5i4Zq0qmxAuRcgBoQlCRZTLu2jLut38Ey6rNJ
HSNgDDHGlbWOwcnoGfo+ISud6Dn0KG2M4mRSIlmikeln1map94h1+akqXC40bhMv6oLC0upTe3k7
ozces0bSb5rmfkOzoI8oWeAoVSpHT3ImwroLkUosWw6XLh1LhWqovbR3+dbM6EqXaaFZP5mWtP1B
aNTZlsej9JKLKd6hfvbZju+DYQP9fnHSAECyJxahrBFa/wp/9JPfdfFQmPmj8fmvyb2Tyx/q38Hm
M2Mbwkj8jZKdDVRuVBaG4qPfRQvDcDZXFf0pn0v4G+JMquLYb/vqPj+xE6Jb4eA4+AwVJ7eo0YYF
4BvrRtnXNwNulUJBBkG6TX1IzPKoUqOy3hV3GizzdPaBntbUB1fAri3x20R+62zRNK6ll79yZB9o
KpWgntnS+O1QadR3Q5WSP4eIdJnGwXozEI7GBHvCRK+ybRQGkIkGf3toKPS8ZA6p77tj4GYLygmj
oUTKYCPfd84p+DfcfXD9nWhxUPq7V74aB7Ptp9gCG2C7dpI+uAhwX19n9OrXIPa+Pp+qh5KJUeHH
95GMp3BKSbg+lXW63rQT8M2Vh+A946PanFvx+YM8OmNvjUghRGZLHAscQwPw/LjeQlxRJ50siL1U
TZeySupR6C1GyHmqqJ1lmnkZPjyW9m1bvnvkvFpQDVdEX5EUzrjQfhprYxKOAkwnlh4A12NmJ7hu
sXc8LQhcCoolFAzuYr3WqgIzvgj/xJ48KmlOgufAMxb6ur62jv7wr1ip+s76OdR2eUJl2/LHbKZb
1qrEBrGOgEIAH62SWmCnbjiwg7Hv+gFPbQ9mVOY7qrDi1+xldw/cVBp52ATS9RSYc0pX901cgoLr
6nArFI5nmoJO3QxmbXbLenckBMOHBpyEx1FrdgK9eoF0I17CqzwXn2dfPv2Sjl76CWY8Z3LIL85E
xYXZnAPHTYdJg7mnLDLWo1xwy8JvrOrOW/E2TD9QMV6zTdmQJK8TqfW2CDf5xwv9sHPwqwq1YFlM
VK3mgGSMYwdx13OgjRsLwTaGQfnsnqQz4qZcCVNAYnkqpIUC+aLdUj+aejjnlmxH2URuX1ez+Q2g
kbXcmkZTlUoET9vbai38DEfGbkLsYoD9uWm/jMTglKIE9Gr0az4kihBU0AAuqfQTJEVD/DRaq3IK
iuq4+vUTCyGmb7W7HRbOGTrnqBiOyYENSazDgN4n1eC8EKgsFXUxjnRnYzhNFWY5uZ+Jyr8OPVop
zSbvPrDd5m/vH3oVBSQesfdg6014oyo43wTMXrLMgxcLpgMcY8XME8hYqMi8gC8sfSJ+WIAobbIg
Vkz6E54xMi1/gM+HxqXYHgLTGmSl0gIq4Eostx4A0BV67LdL4UmE89O7RMka2eCJXcmKh4nsyPaS
0aBbpAk922vN4I3Anqu7DODYYnq3TnlmLgs1nf7Pt2D7Sntu8uzg1WnObzy24x+W3o9X3fgmoTY5
4JGoR8LHUEwrqVZSc0qMIFIWue2QB8xZu+KnUNB3H+P31qeTk4OoSeUOfngJNxDybEswV4zHcXYd
mtDJeI4xvdznOdrY9gr37n2mSR+8AidCkvCxAuuTqnXX39i5LlLMfUFVCXYl+WXxqOSFOkZzcZ78
x6/ZgR+70iL/8yQUD4zXFRDMDlJZdOeaS+m7k00r/gIaiteOrx61O3cmqRUxbjTGKHuGpZlEugRc
h0dVvdxnHEWyllgPcy7LfCtJGCqa9tX5aLMSQY3V673m/7yEB83egbKT6V7hRzSya2oeHn4y7+z6
xTO1GMBowNcp4rZtg5es497aBTD6rSwx9iFJEX/g1MxOmxRKB8O0pwP9DYUiPuao2uNHo4m5KHWw
dQQDtS/XtTbTxyi+SWiQS4DNFJ/9/xoZ3EiMGRq7d4Kj4kz6ULK7kW3zM3xhk2sXx8tZjzscvp9x
JwLzE/mVCnBEcwRl6+x5WDC9YwTqhuKdobZpHMjzO71luwURmwdQ+YrNFD7qEEhHag/vOH5pCmfR
zS5utpQ6mGa6IzKl9drNx0I46bhnwzOTKO2GsqHdTeeX0e8guF/Tz+gsWemRIskct7dV7zdr8FiJ
ISKs131rdKDkY1g5aDnYAf/+mKJQNV/FMs4z5gzAMy4o/2ei0OPS50DmG9ZwCEOIEpNFunHIrysO
jKgllHW/m457nUcV93P9O4P8gHPhjaU37q5rTsKF6biIihS3qnzWHfJYrayYgWYTuyalj1aGCTPN
846+1GEvzZwk2qKAcs4A4aFxiC4obOo8TE+OcQjSIB8f7nmQMjOz0qrPBfkuQldDV2ZGoz7oQToE
P84EzJJmkQOZRFOhrge2FFBKi8WajQbtEh4f8ZviRKoQJ7MBLfdI0WLH9b9q2gWGPgRlUwQcb9TE
fQtgazAY9TFMwglzyCw0yPiS0Fxgi3o3/vgyAJ+uVxslJJOZDabW/FtQBIKvvKBB5k4Sxu7U8zzi
SefUe3wTyT2ZO7O+iBgkgRzUZPeqIm7bNcgdBMZNKnfGfyx/GBH5DXddduqw95p1Zpb5cFtkkYYI
0B8JmrVP+OpDVhLO7kLj2Fxa8dwGqmVY/gU5dEBy31DplAWaH6YS8XOIM6YPrFrTZEfHFH+P0hcZ
zUBn6YGurc5StxvqBoXCwaSUBExZSp9/esgsUVhakhpcTmeCocOQ+5bRj71MX1zaIjllqjOm7Q5/
wRu83N/2vwfOLkTSUOMdCct5d3h5ZSivUkjNSFMIouk3dmPzZ5ddRhUgMAWkiXhdDJKIgpZbmPwy
IHehxlKc82NcoBMfPDiwwalCCfCErk0TuVthqPXfPm8L+YxKbJYxWXsxCpKKzTBUFGbkrnKutPBb
xMSQSEU/vjxYLNFEfUqcvKZp7bE0DUKHzKVtibBiDYN4QmMD/jTOZwN3TNYnDy1zpTXUr4OZZdF7
tSAT4WjIuLvVEUG6PkrBxRsU9B9IogEG3F1+hChOkp04BumIy8b7/EIDzNDRX/2dFlUX5ie8TNs5
gxIEXIcqID24fIi0dr4T7mmHEBOGH46Vq+HOdcZlWy6xUho2ZB7hq5GbkMwlSkzP5KoY/klCr35Y
IeKGSC79X/jg2/Xdjy96J6d+3LHj9uVGtwWq9LQ7SiwQzq3qAqVYn2bHVshUc8/P7/oOd855q6kS
fNvhwJHr/gbpTgFjnik5jvvAYf/maUZxzalj4/M4JvtpioY3c31YOJ4WgsEA4BmeDg+htLDBmlpG
5eXe6LgijkKxB8Di4JY0gBKlOF0Hces92y22hJ/QsjUbrE5HKpVtEG/Ao/q4Y8vNaVkC/L1b4pSK
N7k+QPtX5YFPbRrYTAC/6AHdPg2dh41l9iZZp4sReFbMPDLgtCB/AA0QW+h2YvE22u61yKzzZNaA
gDCaOGXTuyyHSWWmKNWuzfnv+uA2ZHZbYMg1wEisd/hfLcoz3roWh6h1agx0/bcjNhJLyQEiu2Os
gLymzkD4xgEPHs5y+DuGd6ZqLU+BwJxW0ewAiTOFbnuuPh+cqWsRpgNJ2jycj4p9ZzTaBfAqVUS1
/opRpFhNrexjvo2DO0IGIMWpuVrhxbT0t6XhRHjCjpA4ULtaVCcxHg7LDqf+5LA6iWrko/caVZvQ
4mh4fu4UfkbUlhCLFClp8D6xabvYqcUfsYa9ccs7/Ljmjk7v0hhR23xZhmXqQy90MduuI+pXIGPs
oLLmHs5yb50wQCRvLWShdrYULzknIzTDp/TTiBC2neaSAevEZdEmPUaG/g+lxhhdw8WkroX5/Jlo
9S7QpZhg1Qjr63n+9s178NYFoNFdAqLEw5GmqkT+Xl4uTjHNIOh1d2uZjaU/4yuR+iGMlcukk1em
emIbPVVk0AV0c4PQRjR9kKz8SDUL2xt4XlJhLMXlNDr/rZb4cONoHeINsOqkL88Dsqmnv2+dp+Ak
H53awAPteTl1G0MJqthf+cO5V3eewspBF0EluwuApCWiTcu8wka7M0TuarTgCfcaxvsnWsL9aPKV
HgYVMNAhxgDQp/VpZgnk2ihRPvMWnLZUguB9LvKi3q94aLgcVZxN8L0649ayG7bvlDiYsgBBIFzY
mR//uZYl+EIQ9rfraj5VZHd7KmcN2p/4gkmgXWL8gwYf4Vz5Sut/ejAqyC++snDhE2DtWGFBf5wc
DFZgJ5vvyqBCvkXZ8f849CKoDAN/EsKDc1yQR6b9xS22qquH6mtn9hhWp0AcdDtdFzC7yYDKTQKZ
vPOjVroIOsWyuGN5AxAF8wuRscQcpwB4dyjgWHe6cldlMvyLAJmAtYVslEqiR5Pb0EIIAUV45Rfy
v68bOFmeBvlEIH2KWA9Q/zH1+weKKrclSZUpPkeJzXRB/R6ABt9mnY0XD8onhaZCn2k+zWIh6DRt
xe4RUedQlpy0X/PMKVRq6EXUH6dqMtZMdVNwNedhQvlve3NqWBnFQPHTqSuORsBj7GPAjEp8EWni
vBxLPcGbBH1L+U0nbTmwLuW+G9BcN8hOh1PbPm92MOE+mpJgjofxk3lJR4nrTpZeZKxxv3yX+ek5
wWd32kxXhgjLU1bFQAgdYJOup2UK5tTAFb73cx5ASuT3VzBanl0DtP/KQnDH1EhHIYMUg2bWwGci
AQLG3t9ZvBawpq6vCNerOL/HrgBeK9WAJ1H3lmEJZ2aG+3Hw5J5ZxLjHGpCJssCmGgm6Y5oGs8eW
h+44ltY0U0q9C95oYB+Q0NSTGvyWviRC2at/47aGvNiIWsn2jAr2MoYO/zM6zA07hpoJCSdBjig6
ClbAoqG4y5E/24b0OBQ9WJf9d4a6Q13Jtv+FJpYDUQ8JUFtWRVeQ65+v+ayAAAE1iYdPTCMv7H+J
JNYGiYMsNwPnQxdCZk+x58Mye6OfJnZQ66T4c8XV1MmMCidB4G9dXYUXC0y0iml3nD4Mi9xOHmNX
W4nf2Xu/0nw+0oFcmnCM/seK66Hi3GLpNxQFIYdmZWTM2tKs3hAkMXXQN2o2vs7jVRp+WW9l0Xd+
x2E8A21X5AhOQtAwDqsNCT4iuXOp21DXtVOPHJ3dIO8m3R+eUn432/CVbCEiyp5S+DOzassjz3f/
smphrGv1jEsItQ3PdGGXifT3EX0mBmZIJR3uet36oDeFqVq4qyOrHvN4R1lk8XfVHNO9GZeUjNIc
IK3SjqXKkGasPRlLZSPFtgFtBjRgAnGRlgFpQhmdDTVxXJ6TojFzkAgMIk/h6EazEBNvEnAZClGt
uIML9DGPdAO2csWr9V5929ALRKR1Jf1CD8aVLqcjAPAt3Ac65HyqzRznKQzcBPtBCK5RbR/CP9zR
GwRR5XGHoBh3PM4IR+1JjTAKX6pJAWWRl9ZOD5vchkCkxzcVOaMtGO4m4OWwaO6kqGV5q1Fxs6Ji
LY6kK/EEIyoJL+Ax+tyTpjKhd0o7l1PnWW/Tl+wXCNRAb6y1xekntDyhzH0OVAUzXb+z/gwwcNOU
mPPuUUUZiyWa1yt0gueJ55XLOes3KbF0ISQaMQQ4ZxNiAIUCD8CfzkkEAUnn/SVtwK14KUX41erR
KvcTNPhHFpIabjEDl9fMtX8aPX6mWRgT2imnGPlMMtiVzox/2xJ8Mm9aV47tZ8VnF/T55xvwOVH3
awfOrlv+MN0xrZ4i+2RH3Y1lwH0J5mHDwSq5/ds1BGQU1IIIW0B7kuDBNqoLBjiCBnwirl/NzFUu
2uM61g+4Z5CnznvIW5ClzX13SfU/sUAD2I3eoorKpod1O7rWz1jJbCiK33wJQj8+s/5q7y/CeB76
U+fjwq9pvrCGX+KN6mfYiMrByJRqn06OEc73W+rTj4OGnWoJKHrDlaU3RRDcOUWl2Whn00SNMvFs
LKIr6wrwRt+xhI+ACcZo/vQwKtJoBIA42uWr9hEr/s/Jo2HT9k328IdMALLACRlnonsMqHJrdplG
xumqSGup3fssXNl1qyzW0tE/qtaTSKcwKq+EJVYJAfDgd86R8i5bveN+7aPXXfZwkEOwopiwszFV
DWPMbBXmiCb7NpLPkjh6aXl1O10G3Eae4PkM/OsSrDeRLSb22Ym1PjNjVj1kR6dyrmRAfXU588mr
b98/cFjjOAxqci4FpQ22QmtZFmvG7/84JmaD9D1pJRMJ6aVAOcmSFQOJmEqcWcJFPvaiFgTJhwdC
K1ys7mkwtAJduutV6YC6g29YQXPAPg9QhpJSRSaUeRnGDL5fLDtVN5ISUcVV9zqT8mZYfNO5mpU8
Yx7NDniV6asiJMzUxX0eXP1oWYsQnEl/R1s9griHBbAN4F1wtSJUjf3Phx4aWrpqJ+6Zv+K8pMrL
hgoesedX3z1UWOodc6pwBtLSRXMex01kYGHfPvDbrZeh5RH75S56zhbbzXY+IPzkIQYKveA6nxDZ
JHHhf1etLsKtTHrqIopMKGS+G6rK9KcIBBq3qMQGyU5Fc+JR8wd5TgI7GtNuWRZbhm7/bjf9lRNm
/UYpG31bFTNW0jJIyywrp1rxv2s29TY2wg33DwpQfXzfuPvCJGbdvX6X7BoTSEtMHzZOQOJCAcBz
5PQh8y3jTMMtAvrC8U5AOytS2xJ4taPvUDF+E11FAXxpEVcRrYYORrXUwgA3HajnLC4k/6sd/TM7
hqH0K/D3v6xRbYlcX+frAsmtaoo3GLbSsCTQ+WH88mpQVsl9Gejk80BsGrEQy288XM0XhMnTe2XA
7h34dZEoIGBTOmq7qC4pxnzFGKyO2neWc3sxGTato38GkqFXWeF6kLbXQtjjEnVFvhaXzEkxRveb
m6ewhinN0G5I5prJL18ZOdgZlVa95dOvrQyM48KdyIEnMsbICh/nEu3rumJuXUOea5UPBirn15x7
TLuhS4SG+tXEdKMwDrhfYTfp4b1KlF1dGAujQJ7IAbf1egjq/Ha839cuRieB21etyVTMBRu1YcZH
cE/7/IoXwzjL9oGhFbPsrWR4bSm2w4D2XFvUgHzKyrbqr00VkHFJCgPWjbT4jyrdOyueG77xacm2
YrWO1T3+gvS5U/PHq9rIlDoPSi3sdvvUDN4TKtnZIS1Tq+y5i9q39N1OfmxCmOjh6guRVsIayK9z
PKY3Ba5StdWD/BoLCo8iLys3Q5VZdV/Cd+UIsei+iuQ9aFcHlO3UNiS+VXD7+3Fj3xkBH3i6HdDo
dtJhK5ZpjBNGsG7+PW5fw5519nE8Pzmue6smtPLYtQl6OHEpVp8kGUca0L0NUpFRGiN/X35HRNpk
79CKp5kC8Ve3GRuoLi1VSK4C2Wqw+GwzOt+U1jCUAz7F3RPV0HP8xMZSKfAluBurp/4tVcC4mbLX
3R9jIpvXQibfmDBwcMBjfJNvHwM1f3mXgTi/YLdlKiOWgaXY4uukifI02Rv07xdtBcW/j4skz3P8
Y/g/YaKLyGkXp1iSryH3H1FykOOimAhmfMQeqVEB4O2/PLgNTXyqpr5JdywC2VRY9WyIcXJfCLvW
HVVQ2krGB7jw+e7EP2E33l8I8bPncz+GlkTIWctPLeMjnOImm2MTfpgGdhcuapsMmpT6L7+ffOlH
fhG97/MfIem2ROMLa/YgkSsPORCryjVAe8+iR4hsoNS1jo2+oEzU1SzjJOK0ZMstU+RuWq5RIh74
h5veHnGIWe/8jyLEC6nRGCvLo2QWi2F2kn6ZbBEx1Gpzq2FHINJgGXcIJIPOY1Pbi453ajJh8B6F
YSieY9My+p5AcOrfM+C9rM/UaP+QuiWBNj9UtYU3tuZoZWUBz2aKiToSzdyRNENcFauHVc8iJ3dd
7iKo+J40XjrZuCQKpDx8fymo6jLQke5DAc7rFHUQQF4+VadMQy5J0Bo11q+965zxkBlqZj7p8BQx
gUsW7O+ylS2lMXiLSpiQ/SCyrfPkCAtAYGnUDWT4TGDjgVJ+fgsf5fdpAk4AJIgtDiq1IxR1T5T2
oUIWamUUKEYu0pYr5gsT2nrK03frRF282zMt0Xy/zWspE9Pnbg70x+igp7+dusjppPfg9yakZlSD
F5vR2u7VMLN7/33UXYaHw1iYJohhfvfvE7im/Jz4ngZJYvmuBWs6DPnCfXZyFDStmdUK0Q3makpf
2fwbGC7Dt7OhrD9pEr6Tmar4BBNzbcuQAsclpZDMyZhbcxRacPCejKcGWc5wSGql1hNjV7ywwa0u
+QEacgWEsvXQdyow7AairQI6wqg3hMIAMeKVKkv6VZ4pWiquCPgM/kZqdUeMeAI1B97kWwnNJZhj
lun3QrdE/XnfnM++nSC+8E2g7gSHdUZG3408WYrt8v4JF6u8ICxUYhSwwg0ct0aAbIuQaIuTJYXe
ocHz0jnXIidj3dSszDDOj7PXeQ45BfSZ+q9pUNd4sYIqE1j9f8pkRlFGPDHFFzR1Vg3mRXtOXUbP
JEFMQtAqgTDahzDvrW6EKFfOKh2XO8uAjI0ygs3Rzf80tmmdT9GyYbUGilVVL4SCqQTM0+SxBVjt
gCPrdMgvnCZzIkGNOQeTgV7GWA3D7q6kUNjCgxAajFFqqFlAtGUoPjxaMjc1yLnCCtAI7Bk65eQX
cxu5BbMfPmHF8RQOTWMGYPgIu4cZ1/TkeDfjQOiJvRlWF0lRTYP0kGPno04IqeaBjXx3XhHDNMVI
dNXKqE+1nESZ9gS/CNIrTn7eg92jHF+RggUUsi+e9IZtSh8yZK/WesCdEMtJ4+IKAytPkemeblQG
wdl8fn7DGIhd1wqJm8ochErb0JDYbqsOdO1Kl59zfoeJbHPX3knGwlnqe8mUMCO6SVyu3WXep7op
3Ber6RPCsV+DR2EfxuX/gbqoQqlIcniWomhcXMU74CxHa76Sx+Q3bNJ5oID948vEUsZ6GfWh7+o7
2yMLPdd1atebnQjhWlLdMVC43MiJlNxMNeVFr5ubh42mCjxqFlw7IF4AMfuREwxsSat+pkTJtxfY
Oild9vhSAN0H6076Tj+GF8hIo+Zw2ehsKj/HltjcXqGL/saiPSkJmg16SarjjIqWxLDw7WemrLhG
W0D7UvT1aEYxYp/+172YSU/o3cu+6aU9KvX9LSIngyTifs8Zii8w0Fnb13DXgRzviMwDwZ2bGcuq
b9N/Rb2z+I2CZINacQVuMRF2pEFyQHAtx9uEaxS0Zv7l234/1Y2R7vLl3weN9WrQRjgIlIuvKG+H
80/lQxPZx3kq6gYzreBl/DF5Npj0GhblEO26NlJeOxuykDUaT4OM0jND0TgZJLEKxKyqjVR24tS0
RSsRGOChnLS8qoCPbKXIr0+HTsWWuJxnS9oJj5xAEehBtfFShdiudosloA81lC/YglXDoxEHThKQ
S/l48rYldF68o6DF1GoiqRUMUWpnXwHoEZFkscimaDLvUa5tqacD+h3uu7K048s5KOoTsvDmRzJP
mwQ+D1oIIuFeaX7c1Qu29oeqtx5n5y0G6P28w/tvUowB/ImqQ7+VB8sTNdqJ1F0fIKEYvQBMPA5B
DeB7gDk24mV9N/0MACazGlf63kbOj4A84PN/c+JrqW/EdF4BIqLUdjLr5hLWICKbwvkj+rFvJEES
c9a8Vb2/rrfwMQbdd1W0z5AjDcrGJhyzIFfpV5eUAGADHhmJYMckDcAWtCcsfBeAVV3a20uvmfrV
W4xWDRg8UMAQf4zXW7ZHLQzf5vCZeo7EGF0knY1Bx391IoeDvZsOfmERczbQ4W7eTiCXwJjNqFOY
2GGeONbJkUkqgX5bRzC1dHLvb7/YlXYndFCu0h/ePVxGySZ0XmRn5Kha8XIC7g+gnhDuYPxPnxYw
lXNz0uGuR+jMIkxpZpMgqbXmghrnga9xoblmulV2af0ETmEboJKEaq6O10QCdV3gaDv/qRr+ZRE+
OH5oahadcddxgBNSANVo5l8I17weCn6uJAJJRpx+pY/Fn1Gt3LbkxuhViUH3lM44OPTO1MuSMU0L
qXhoe929yHoCLr1rgTdTMq65XxibMrxGbPBWWCWNnxCkq6jzCZpMRdUZv3d4zRej5P5dPqMZkIAQ
cOnwk0jXMyMkinf0/5YV8jSbCjCZNBjEK70fAHsqm51dTK27AfbAcvFT5JLJwTbTSZ8xp8sbgUrC
uk4nYTOGPAMpKCd0sduRHsQ81p6Kr/0gOl8ozWQqe41T6cIe3GPT8flFgLQcW9RAYq3v+H54czYQ
xLPjQScR7wC9wQI2swONQcyfoG9NnG5+BNvvQNMwyeRhibXpOooXl0CgXnEX5/0RUP5dDl9ry9jm
4m4bVan0GRFcbpV8NRf5CEohAwxFBiA51nH+V8mXkSfgpn/QdZnUCrYHqZ9sJlCqG6L4Wn7BMmY5
/ERb+xJBeNbpn2MvWCmULohUh3VuG723CMqIXZaewu+fzmkpDImGiFkxMMooZxMaqYSeX+E0k40C
jISqb1dtoPzkJgydhw8W23Nzz4uJg+K0FKwVaEk/vZACgP6jzQr+Hhu0W/8i5a2F0RcqIenqM5z6
CiZ7VKEAVNhon/VSIqOUvR/9s40triVICZr0XeGYt69lr/4u2ML6csMzrEaXvCJDx5kodituTgFu
TgZ9N1KTcZS754sBHFzHghqNNsOpNVbDdsQWcl3LkPn7BxzYcweq81BDvl4LuVP6PJP+S28aj4M1
b0LIPNg0wipfZHe2QR2JIzAduWA81BwmJTmMhYUhq52t9j3dUbFobRrzUxBtTwem6qiVlQmvcslk
H6bxomr41izHiKyaqLVL99QKwJZAQUWbSMa/97QekYCtEnDtmXz/4HbpRWyYd5DnUTzFfiE1SdeZ
Aj5qiKrWJQG0bC7tjo3v5UJwiaCIi7ic1leFa0ZlOQ76QgWyMhRPrsQlyND9Zu3loyUPhcMDra61
cSsYcep+B9JX3LKyzEi8RGno1rwJ6HpzncakikzRGTNj9DYB1RgSu+n9NJ3t+VwJdfTn7Dz8MrIM
4g6KjCt2k7XX0hF40tAGuYYlF3PrBS/JObU4z8iY2NQjSH3B5rq+PVeq1y9SQYYqw0K4R3psniqJ
qUYYAd0PqY65pP86i7r/B0vHRMIcTQ78tVkb3vlLKo1GSAa7CbnAGBFCaBhYeQl7uZr1vVhnZ6/w
7txfaeVmdjTqK2avHe9P73rECpDJANbOBsN4K18Gah/0Lh/MEdn2CE7vroBJi8Y8TlxK7UakxisC
t2RIeYIYdM7ZOP7pwMVXCQaUK38GLV1u0BvRQF+VB0VQGZMt4ayAOK2Jp8sZoRRTRhtB7K6VttvE
nWpEVimSg0HlpAo1RwlAghNcs6jNVTQJpAOtos8bL4BBAp67TLZryYfU6/glvy++BbJ10T2K3a8B
sp7/SJaEtWWLvnJ+QJ4ElKnaW/UxBYo/ln5Fi+JOEHo0xuulRbyxa4wB7c+ZNJnEiItYktInxndj
x6ZNHZRBokeqqwP0FbA4QegvpqBAh/wAyFwC7VTObrl472EqOtC04rCn+A740HfVVmzqWaKN/TjV
x6WL7foCUsg+paUqWnZvykNGXS8GuPfnruA6fF6CJDypePCXE18M2j0+pcrHUNA/vDLbVFj498Qo
q8Et5UeFofNILYEnIb0qEFMeHPHhBHGn2lFba331pNgKN6mOS2hcgXRmtmqEwfif6lj/c/2KAstg
TFj+ggWAe6E1I6defesO7ecLAuyChnRGJr/UgjpfwdO4b8uNtntI6KlZxlyQrO1KLvIiSIbVWq7X
9TweyfgdNEp28swATIPbeKr58L2JIpst9hH+d81G2z9STWzEM3YiXhLItIxuVRHj2f2LVgydDJcF
lUHDfquDC0ZxprV1TACZ31dQOlXVytXQ02arBAsCpjpUvjHX0ZBt/XUOCD2kGp27RlwBnHXhTn3H
Ox4BK2yobXC25ESUP4HF+NkbMooqWT71GckUZ4vZpzL6cV7CY9Tiq8k7t4dyXDnCqXDH0Aigmti6
MSjXGXaNB/uEust0VRZiFTrkyJ2YoqIG898cfREr4jd68HB4fAFBJuTUuGtxiS7lfIK6LoBpWomv
h/UzydlST8OhuQU2Vk4nPqt3KvjFPksBnkdIwoYVAiMcpF03MroEI6vuYk6QhY6lPdUqivUItD9o
ccETcT8GO6/MNKUoapYaXEJUBl9fKF1PxqZVNZ3wjfDjK2L6lSyOGtP7+5y3COhfLozeAeLBr+Qf
wD9GCvu2vw9eBW587No/EdCv0HKhubVTWNUDjcGfXZUA6gi+vW6xbWqHiYC5Df4DtpEJON9/wXCb
KagymJ0bAo8auXICUWbU0S5ha7xETSG1qeuE2cuGkznj9qLi17w9uFaDboaC9z4ofsqhL0+AsBJ7
VoriNQajNDgRvZaH6P+Yy2gRqGRzuYaFnD9llMntVZgfhGlOsQaQPFmpDaiutiMYXLCG1Cc2DLs3
MsK88LKudnP6vuWnIaB/GJE2PrWyjUrUtoFMeoPOYeTxSazDhFIwsjEhAyuokh5eGNWegohnW51e
JZNPHKDV3b7V7+JzC4XQcYd2nziZb8NE51mNRMZbyx/gGwTR/FbP2EyuUcnFC8MZLWnMnCkwBa+r
8RMaWMgMiIGhKuqo0CgsFULauJUkf3ciNXMZ77amffJ6odJkr7GGRwokX3QqGdcmdsStHPNTa9aQ
yc8jpKNR5PN3y+HP3qcHxiSSms0cwzz4FzFXr1SZjqBF/30DGziho4uMNqVRZnrIvCSmU3xjESxO
XL5m9bfZaU9UqJECHx7WCo9/zGJm6k9996uuim7JLFXYfzjFydaFdW5pGeoMM6hN1Uvq5t1SJwXn
8jxrRuGgs4DpAxoJph6Tz5e+YUfJobYgo58qCZnJjmGlmI6KsMxg751QnC/0g20Xvoxr94C5lbQS
Q4gF/Ad8a7Wbwgqy0ELLinur+/4tmjvSK0CcYz0kwuwnPchatrlp+7aC0+B+PIScMsL8Urrk7TD0
D+TjUR5EtLlbXbu+otJoN2IeC311xWrtonz/GvloJpv1V/4ixyW8PHOGcEe+cZnAbQQImoJBTKNa
oMp3O81fEW16A5331VwZUTZ9FGQDIOwDRNec+7YREDIucL5W+dWPhFsjo7azR7xlW37EuVPFJxYS
3NX3dXVx4TTRFcHN3DNXNDR8u3RWcwMqdztRTeKFUeyZBmh25+5DSPO799RlfAL/waKc8w04h21w
a8tq0PKmm4wK7UsJhKN9+SWF72u30LCqvzI4NqREsCcid/86mLCNRDIWdqWuZazh9kLy9S8noNGR
G8/A+qisIxlOIQ7jFOJGgq+lXP+TXiAxJ1St5J+C3dfks3Rpf4r2vOSO8Mqf3r0AOBq/opm0uKEI
UsvNhs/SKkq4vrRWu09+Y+FSWdcbahaDau5L3YNEjdMZsbealhXSr5xxiqJPbqqX03OX7/rzmi2F
SLCHGcCOgSiAoImwLeY1Nz10+qZusSTcY9okkOmC1UE9uT6RtnScLzMFoQ3GKMXTiiIORAn601jc
NVXEzJ//RPlam1xLSU9/ZzCe4I+BDQZUqq10U5w15aw511QOUuVqlb2u5NqekQPacBk4MQDBzFpK
R9hKD9mjNcS3913QIiNhauOCHVc2XsufXOw7GPoSncg1aM8hgSpohduHDJnEIBth5R5OiHFJmZld
OUfDBT/Yh4gUzJOg8idRq608UNKdqQ25FbtcaEwRJSW8PNveQRrOULngl1F1JW7MNCfLsD72Mu9f
5p60jJwv+tfE1qAAC4iwtQHmT33/vA9VN+/tbt5dnwsECsDkXfCU/9c/HNFR7MDz3mSI/CnE3nnn
9H20s8W/pM2DWWEveEde56hIIGTdFg4i8nXdI5FTELuCS1hvKPZxvYqEP3VvzkoyGgvlSvkTlUnp
+evAtgmgDOistNtxhrrUiKLuR7MktUGgvngHUYG7LpSMg2bjH2/4ckd27KTpQ564jL77VlqHzbd2
xwHf6XKvXT9NBaVkfbmmgQeQYMLwjTDxChJiTRiqhKHV92bJ/naCnTf4KIW2S6lAecfdYqg3pQ32
2+K6qLVQJUJJvt2mU4FcruTcA4X50JhdJi/sRfu3Wnvi817kXLHR6Q2xahRboKFohAmtrl1k1KKS
HN/TbzNk3iMS+1HjbLh+b/sirwIogHes1r+BFjyB7iNfYUFyjKMOqoqQnyayd0jy4dw+ENVoVd+z
kfYKJwc32zk4NKdSj6P/6IFXbvlVM+dZnyX1Pd/KgUoMvgxvS4Ov5BJ/kfMcImQ/6G/xZjWlIw4R
sQV/Fy0YRCcSMIdg3wYF0Q7Psok2OJutdokaFMRAr9KqvlFptVAYcE6GxAdXQyCOhe/SyMxX5weK
53O+8vrf5LAp/5QVNvibcwwF8nOERr+jukuQb/5FmgqoGFoBZhFWq/kw/5YrBxedE0U5jLgXrWJ/
D7hMmZFEaFK6PZjL6r8sUwH0WD5bngZIKH8hS37ugQRBhCO789DxlzGbTZ14VPPGhTKkTfRyT610
ATBbAwFLYDWxCQeOvk7UkfbydsKJufEjPZD69YvOoK/wXJXqMe7riJB1sl095nOKv7yImE/8ygWi
X9E0OC94ZjdG6Au0ElAI8kO5+fFworCFu18cEuLlGOaTJjSOppxAclSPlnBGLEQKhDenki4W09pp
8bxNrEoV23mraUBvxQoPAHHHtlop+YXkG0uH9rCY9BJOW8jwKw6wYyvFKLcDnj0jnfrGd+L97fTv
XF3Ops+QbzBSsTmRfLOpfjPDHxqLZ9cPIUEZH24GuA4JMI7c1pPYWDXMDpl9Llf5SHCHFCthWwXX
KfAsRbz8nojvb0vdPFnGM9wCr+sgYEATYhVWDRNCHtcyNATCN8vSHyyapT8Zp/LoFeUKobsHlmGS
XPSMHm3tCPZkxOvhUgzNnTLF+dOSO+1sAIlF/0vczUvPfTQ3sqhaEKHDPNxzj2tPuOSCEUg4ZkE+
XnBOyaBzVLi/qNmmWlMBYc/sfD8anzV+3shHeBvYwvB880sMDd2ivghmToyNwrAZrNtjK90PD48H
p/bRBO096/6UtTneMKnefD+lFhEqWuedgHZhO4e6SmAUtHGb06hs2h6fk2iSUBzF04zaLsNY30Xo
m0tDLcvtoBVIEMgbtrfO6mh3xESXeGKJTJ2q9xuAgWxNCUaygmCOG/fVldh1AQMp4BIFJ7/2VfGA
P6XA6pPi7wBNIBy3jX0+1Y+VecnZBOcDMePJJ/hVuBP5HaV84DRCw1/x27GhmTotDVPQvrWFCPoS
rDWwn9RLNtcvA8omgUfQEmPle3F8gc38/VPiPH3AcAg0MYUwNxyhln/ZX0lGWS5/xfA3BY/HaTX+
4QgDXxs0AwQk7DdiH8fxLqdHEIyzl6ISglHVFwQX05fVW7ntuIgQ7OwrRCm4iUfQJp9a0XHl96Kt
5ctepH83IQXI6MAgyYkkvQyl5YXkpshpYEu9X9S4wWXhMFSTs411mYJO00xmKhwmXS3jjVa6YurU
MQi0DwXVcu6nhXdQThFSjxg6+bJl2zWUqJsK6Q0nsT0Cz/PbPv8EWQMZjF/SHdNdJkoNBIlREZ6m
cVjXzfDIHYK+srMuwipu01c0b6QRF5Zg8kgmafFgciH0/OkoU/AbsqFtuDFh+ptXnJ078BmYk+wI
sTbDfMb/u4K+oEfYqSCiggW6eGS/trPcyw/w4U5ewC3X/jgKRv3HI2Eu8gDciSLen+Sgh6/1f/8X
eUdmJtlHS+QZeL6G24amzeWnyAJ7JafS+rLxQDRVjFcmI9uQuh7sA/qU+UH4KfSlD51RvjQTzb0D
qj0gRODcbuwY2tk0bwPkQAvTFY+FP5DYoMiWaNjmuwKElNZa5s6Z6yt0k5eOEZ33egAsFErPIQCK
P1V/awwU9EqEOc7u9+1PZ0dEnnPpfnSJUwvWQnUbFBFyo/r4zS2/01AvyzPlALd0jv78J+rfqKls
M8GC6TUfaf2SV+aKXWzfK7Qiw1tmFon97oZbixIgm/HBvMTTaNEyD1jlGlBulLetNQ+ptAwDTIdd
gPwVOxLowO9A1jOTZKh1sMdCR7nwDRpmrtJ8j+w/e/gWbtZKh2wGZF8x4QZ9XnVV2uq/PaRZauq2
N7r3q82TUj5clgqukMG3PPMLVVjbHdAIRqWM0qIjs14UwtbfvqS6Dhmp2A40Kv8WUSYpNodPXHQz
e3HbnGgZaDxs6gdlYXNgdEPlK9l11sBwpLs5+UECIE6MK3sC7rqZiYdUZPp6Ty6STRgsrXZbYmFe
vFu64ikugybPiLBLObv9T0Jt+pvijsVlUNGCHyxjm8Y6k9stbYuGx+P4LCCFrGAtXEWSFZHZ6XFl
cktKiFHEGt8L3lTu/9wG952xJX96m1bDbo7IRthCfmVsNKa2Qc4euYNV2DJUyRAZoJ0upHfFWp3z
/ndsK7GFITOh7twh7dPXFwKNzhqRF0/dxN260+C8nWhCgP8UZMm7lwkI9VFO7FEikQAc4RBtP+Ec
+dQA0jp3Y8N8sj00yV04+le509FIOTnMzg+BYUxToX86mUR6BwUbj5SXyIoK4k2v9iWbFYmcpOUS
PvMf7Yp+Iyf2dCnRo02pkfcJzpFHFXb/Qq1LtJCFdJVyJlXzurKcSxNQ+U8t+qEWEZmnpSubSL4K
4ZcPUOlMpNLQUOSR4+KAQGX1C2ClkIYMqrwG6yZoWzCbQQhS+UonpKag9Mrq9R4Y3qb4VvOO9gUo
KxCl4XTRO32ws6n3W3tlqpFLE1hkOKw6ODfd+Ij0rDbUxEkHsGY4yHBSQ0kbtSwQ0sbNhq2gv8kY
By3tJXw3/dhIYDk3QyM9Nh4Py58muz2HGPGyLQky/1UA3p1aKmL1csQT2c+XjY25GISdWIbzv9+L
98CSi7Ac04VH0LOVrRbYZxWYMnHaQ16Ry+aBY0cQpao23X9nxPR7B0QYLcHmQPhTDoBArj80mQrC
6sqCRrRdJO6Q0ycweD8avW/RP/hs3N1kjhu6QEjSlY9R1C7S3lJmH5fwb+NN4zGnWqGESQhVr4v6
KPr63kS/SbuXwMAKzq9t/dZGHtxXSC+LWPNLDszhsq2sFtyTW+KVwCzsWb0YAuWvBemuKFq9ArxN
k56Gtd3AfYx+UljxnpQiotK0rHVVe55xYBNDbUkJvppkX7jVD6shGSBha7QqkwfbslRmcb6lKi6I
ReVFNQi4tRgXBr+EyzRnPmkoC3joKtyOH1cVSIR3jgnTMvlk1sHiTK0/vYh4t7F9NvSzBfwkbvyr
Wzvcg1ddtUnsCGXpZQYI27GOsYQxJ+y9KzKGqPDPHC0ZlUie+kcTunDNbG9b7cdOEP7eMT4aUmjr
DMb2Wc2s/z9sHNiGDOfTM5Vqg7sM6mpeWmBNAHJfmW4fZnV3bSq6UR0D9EJD2nDIQOSBeaxnDaC+
4PDGGnzBCH5hyyBJGwo0GTMFKhE2O0HKO1zTv866XyHMWmmXvh1+R0DQjL/6npZe5FJyAfcLc/wp
9HSdzjtNb5aINQKjlnmBexSOIT0NpxPYyQMlkFgnN+V4NabTIpCotRIguiwDzeSJ1LhWzJQGDHdZ
rldJUMhVbnZ82r4vZcgHjXZuYH35OKsOxSBm8Okx+K5QqW788GCBKCnlYx2HpndlZcX8bdlPM/ZF
XK2A22ykJARJbQoh0YCLQR/m8Wh5bWy39tLlEy4IkzlU4C4IzsjlDasBjoHtDJHlj/8e70JsY0ru
HjSng28ugWIPx1rXxWFlbQUqj94xKZK9pTDA7SokkD0P/35HP7fH2i5DL7Mg3qpfynK6e64WMvZn
OA/QvyuOi0Ea7RMmWX6ZkDCluWjvA/1nOLJYNZZmY0ECuGr3UtEs8K3P7po0FIGfdoyfw3PyKgOD
KkRb7imhw2LGygiS1pXmIoC79aN2SVO90xIlaqjpbEUdi8OyNGlAkyYmgVguKqrk0ySaovFLTlxj
16tvzUj3/fqpLDEOssf4AmUdAJ4IbEEdHZ4kxs2lzSLDnjsnQKFdOMY8c7RFpJY9QmPFgiJET2u9
qU2vfYL0fny8zzGjzR+uMigJuANJHQPYTTwEob4LCbVeLEMWt7rbboljdvglY8lDPG0oNOp83xFf
h2Pa7+m/u1Lz0LQEIpwU1DB+9xueAlDYx3+Po+a3omsi/SjVoXCTfX/NMICJmLorZYxgGL87DhPr
tWjxAH0eK0Ja/dSqIGE7IJb/QQXpyW5pMkCS5UQfo7R20fwvnFOmyw9I1GfTcL9//22YpNKcg3a6
wwwVFclGqc/4guJvt/9UWrV+GxelsBY0VCpQW8Iy5IB6xjrDnh+/ZB8mEp1rszLMzwPpaL5UdmNn
1NzYi8XsuakuvHZ9yL5eJ+S8Dzu4zyzdzm7n5soJEN9IXhFMzsdkwSke+Z4gPn1/AQ2s9UxPGQV6
2KQ7FLLxw3FXH45INgutPXhU2FNjZejdh7MjLAzFeonqGbTUi0lMKsJU435mHLW6MvnkFFCVZuty
WkX7C7D7QJrCjV53jIVVhl4vHX/D20RVVC0qwGihnGJiBIz9KDSxH/H7iIA4Aq4zUWrf23IUYkQV
rSEbPvtrFjCA+jT2hyRV0fIT/Xm8gZ0jKVJBKMx7bO6Lbkt5vEKbD5KW3mt/kiFR8x1AtbTFRzx8
RVzTkCS66buXnKPkRs8bJX3G8t1dAUfab6GXFrXhuBKD+6xuwWh6h/snu/UFadDajYWQ8zG+/6ml
RqEFT9I3dyJOJKpqK9tw2ELnJkLcVofnOMHfv0zkEe+0LCUf2SmSv9upzmKh7bo4I8Ma5pOjt6RU
i0aYazH+kYlFugADQKZKc3ZDbI6s8esFsEp5og/07UCznjkg5YNuUhBUV806ZhR0w9gR70jQlasD
yq0pAzgP83Tc5rIRNpqClRt6ynyR6rbDD/aRcPcrSIRUVrjWatRRXPDK7JMu+nDEjNH8GhL4U8ur
MKNsytiOUzJTYDp4ob6l6ZbQRngUzafXf6d9wHp23L9XAaJf9cGmQG/EnkmGhxP4RYZPxtsHzL07
YmBTAwjN03WM8jjrKIUBPst2/wBuZojwdghPdXp5patXkG3UapTOFYpRIkYzocub0y913p+5uZDf
9+VA+ZHGh54u2c1TJOgjnHNLiDoHmaXhgh9JaJ4m99FUZaaV9ggtvI7g/dH9IcOU7v02ng2lZsAN
15j6U2NJM6gXHSelJxZWhdSoc+3D4FYkKsWjshV8snYd+LueOU7TlYpe+ll8/rySluMjZzFfbnge
GuYU6ByghcReyTEqWaU3EcQFKQu4ybqqDlHvjEqB+w+j+rLUdRkhjhzFLOHbCNeQNb02OTo2HXYb
9A+dhPEPEtHku4V8H5kfhBLcyQkkVmK18OSP+bbeTg3rm0ZDXLMuGwo7M1VGEmn4BtL3/sz9JqqW
VkFPtkL2hggXjmfSSkEngQTVna8ZsuIngpiOVCRrwEXH+S0yT+lPpyXOZLYnhl/G7vVOJPXA0UId
vtos5ssBKz+pF5uywX1Idx2/WtDZYxhJ/eyiLBCq0CjS7vXVsozAeTm1I76+epU5TdjrES0BhPTe
qsjDtqgTrM8HMT0hnHLOBm/Pd71NyfrnVee5faciAPKWVGEnAr+OwiJWhy3RnRXNpBF7i5imMMhj
DuewP7EmOFpCKV5lYO/FU5jRNShDkfON1DQlyFo38wGDE7pTufqmo7l91UtuLj9hSiRSL2JmXDOZ
a8/V6pfF8t4oXqa7VuG8D0Fzp3C9NRbunlgBHjqQmNzCs9bZOoKao5sKftVY+9od+ohClmkMVu0a
R4M9pK9YMkyOyDLKHvw24GtWsbhn9LrAOaylTiyy3KKCmX7XF3LuLQ4pUmwRHMhbWqt9ZPNWXYFK
XCZp8EDw4UQp6tCSzFgjYpPdgC2sQ/eRLJn8b1uRcaE9ilmz6gFte3UfAS02E2dMIBlGbKrorUQs
XGS18glrVkcXpe5XnftYL13ae7K1lRVFb35LhWlWzp8BoAfz3im+7SE0TPbSWSiYnf0fmz30S9WO
Z17eEPKNxDHls2Xu1sRzgibAOf/ICGsfbTZjmVYV1HuBdQuNXfFo6P6sBmtXXKtSnp+j9lRwXL3A
tikf+ywXF8bT6GKsm74CpVJgC9m6mwIr5UsJJzlU1ko49uXBT7LgM8nj6K/zmyp6j9D3q5r4D7Yv
xpyWjkWK4oFEXUKwpTiuxlZxMWX2BBl7WZ9IZ+6adYLavuie/p013hbAV2X6srCYM4N+3Kh1UvH0
/Qm8v29zD08lEkuF7bGj3huBfJ1tFi+7ssXxBfJHE1558PBhqyUC1AkxQ4aHOPl5/GdfJQ1AaAlC
OQzVijZu3PTVF74DvMNoz+vMfLXrjeJa2//IW66U7do/1t0CHMUCMZSQXCKCWvMuSwrNIkeT9s3Y
/VXsSsSPpk4eCbSJpAbEcIswzaArJZasUzq2ZpXEwr9MuWtzuaWdZfOTV5cRvNSnh7mRKobV/HXd
rvLJm6caOlHm553101Fiir99Zc1vjbmHR9imx3qDhb3GwDwHTSOSkY66SSbCL9X606bbCMh9fqCL
qrv1Sur45nsnK3mUom6pI8UWmI/h977bB1IpB0CbwFK3JTHT6K5ut4FLDM2/07Y4i0GPEiV/ej0k
pc4e1ZND6ifGSFIJy8hanBwf+lZwcPrD2sHEFu56JyJlMvtDlnx3KC+7qaOtIvl1kuv+hECbNUkE
jeFWZgYEv0qfvoVL47vombS1VxjqdlZv7WE3IW65+DvHIH0hipZvX3LP/c4wtBuh0g9Ssq5IJ79G
ae98W2whViLiUeJ53Aq1pDTCk/smci6hx6PJanQMfSWIyDvGDIG7NYHjCcVLYPQSupk6sXARsmLy
taMQLSfFBHDbZYvSfiHckz6inFAXGYj3QIG7KxVk/YdJe8dzocAKre2M6tza1527Z0MrksjxAtmo
w/Iecl1sdgVUheQrY7208rDRtLx5dxM0b0cyZDEGYOTVHJ/egBBkcmLOWA8/jXWZwqmI7Hgth2o7
HJomTdEAR/J7ySUWfeV+HeTu/UjO5PUFWssn3Z3mivGNKtiaIYLlQVQOsvydJPHmJSjHok0d1uJK
M1a9dmVN+TuFyRYPTqMS4nwPfokyMNx+bQp6LHUhs2DIh+fhyWBmrxF+ZmL5K10AoY1Dd/tg8wsM
7ob9V+XpQEGaKEyZ18621uANqR+TNrR5GTawyEjZdj/VlwnSngIS6lPXMq72wlrsN3q/NxiGGLac
V/XeAcdOkH+RT/dOGwPndBoxMoKY2RGlHkBwSAMHnky7BuuXceoXPVfmLomcP0rACLYvvSVyyToc
5fXmPWYk5jDg4aPDzSfNoCh1U5vNiJQ/LwskEbV/r5Uzj9FnBjWCBZtP873oqHHslvb7axHXI6El
noI+4eVEHDyOO835hCbg5cPacJ1xnR3QF9hLJRy9gd3Ysd900mCzpOyf66ygDRg3Eh2eZFztTBDd
Xaw16BLEDLn8awPYBX/8ksm9JQ1yhjKdhb9bjL5xa2ElDwOqlkEbolSWL2MIc8FmVFJOSh/v1KHT
jN9VRMLTo1KikJVHZHjHYHTDZ2WkdQ3Sq2nfKcCfMI+y5mlzPYtIxGiwacc/G3SOqbgoKix2o51l
nB+wGERLiA4zrKBI19SisF9d9eD4cSH4P8eHQo7ok4FwUurHog4wf9yd7rEcSe9hqs1yYnqep6yq
im5Cm384JkwiTXMciieoOVUDBQvJd1YoryV2wz6lbtOlEXUeiJg+9HoUFD9HPilUxQkPxGXXIA/b
fBOiCOvMucRjYOSRMeYhrtezopCEo16nZ+HNKmdIp3WP2SLAxDVgrcoYjYBxIjZS+9KcPuy9JSQ9
W5tnThIdu94YBC5L8xZ25iGLTIkhtehr5bU/XT/MmjTI+Rlzu0ILYMs09NpHWIf3EgWxhvY02dIF
ctlWC4NgxYZY9g+gC1UCf6M3SgTeyT1pUKz6id/3qHborjoY5dYSq96bQEql5fhLiaWyqmMhTBO4
ZYK1LaSTdazpsdYbEtWMf/CeHMVf+umwcYELovQHpLE91XVqgx0H2WSwJF+w+HhfUGQoYOY1NfdZ
SjkxksrmIhgRQxoNDveGQX5BnXeQeplPxYqbBjgqRAERX5hc78IsX4NR70ODeD1XOCBuywEce9Xv
ywBae13r6TITRVBg3KHECj1SWLZcmYipgijyiHAUb6vDakEYqsI5UNmmEt0Ubi380Qvlr8Rpu6mM
DG6x8Z1RHkDNbXALuwYtwptUDYf5OO69jNBaBMoNAjgIWPubYWcDF8D30RHoahEhLuQDJrwuzw1o
GpEN2SbHD8upmo4OZenC3bfkAghLpUq3JuZjiD5fw8BMvoeRY4JkVxY1lSaA/hJvWgU+ZKY6AkDW
6tb6Aa02ucYuxDcno5ZEz4zymtePFVXJMNyybVd21cxH3vDP8Ij32B5WZE40sESo9jHt4X/BDDCw
SZVjgxOr7GR3jk5QCjUx36vYJsV+mumgy4/ytrkKanCu0YxXR2zO7iAB+9RRori1sG5eG8jvZnHb
uXHfFW/AUouaODXly6ThBAMhnKmPiTXLce68g07IQLDGtiH50MwiiXjuhmfcnLfxvK/XfzUpr9CK
pf2QFO6n2YREgthL5SFwBkMot4g/fV31lv1JMKo3rfV1Cdl7V3SAcdHbyI84zFSvR5yW8Pbd77sK
gN8E6QO+b6CfKg2QLfIvqCqAUjFKhtgK0ADJ982MUZEnfciH9Xbk6wmyE9mFfSF7t//+v/TjQAsZ
W7d4BV8ZUKq+WOEvTdWeGLP9T81/yBXu4hWm7S/Jl2EybqlkqfJ89SmmhGviXPqcJ4rxRcUDS3N6
nUnUu7TAtkbuMjxadwfzw4IFtrMBbsTgJ3BpaTQmjSAnsuoRehRZ2Tjq8KM2O/n72txKCD78N68i
6kpOj0S/1va7hRHy4ebcS0cY9C6cPuB4RDp0+Sqgzw/5D6G0ywIPmqXJnnS3ZSJAeTntEm4epmRZ
YvuUMUTaN+dWaGesHo2w6nS83iLKSQ/QcCAYFxXvNxcQW9QJPYApT+ELD+kedCGVDsJj/l/gLYVR
HvYGKtSqFWhcCvUjl/azWrxlrwfCG065CeyaC5T9rBbaiQQMRPQU56/7lE5nyxHf6/Bs3A4XCjuB
FJH8gjL5MKcKhb5dH40Kvs1q3Guu/+NW/fQJMAWJRcuW3hgfR8Wg4B3FdavWDM8sv6/kJNl+/GIR
DTEue4XjTPMraJQLoodxUOebbaRMhJAS9pW6fFagZ/9OSIJIwIU4x09HgeQKAcKQXZFtkjMHMdkc
GWn39jqFdRVnrXGyRnK7eL1FTW8HQ+cAR50bq/LFopm4jTB7XN6RwCl8OWNZaun4dx1FMh7V2S6a
SNKMr6/+ab5bqC5mhKiNJvqFNnA2zmzvNtB0ryny1mir4TrR2hqv5fBXOg9KU3Xj6gIcihIIOuY1
VLN7DAHz4tVosqoZO7kYonH5GlMFhWVYYJ1llBh8mUKURPG8rFAoX6Vq5ejxEUAcNV8mzQ6QWw+6
1UY1TJSPpI0AzPkWwayV4mxV+PliTnRdnUwwMMDOLMenbNDqGTu2xxFUZCfI5d/auUc3qwgNPo3d
voA7FZ7/jGs+zE7FBydSFkql092flfx1qiCGQFoY1kpzLBsqOVRrtE/JjE0a88CzbtoJTIlkPjey
rQoaHL9Um6SvboSyEt/GxQX/7GDF1/sHRH5GlDzBDovyNAwRKaBbHHaoSNzcTdtFQh0rM62GeRJG
9hdZN0Bileortc6I7bKaEk/KCvSbtZy8FLvDtskj0VJPn/Rj04qZgN6U34UbjPsP8Uhu/QFW8Eoe
MYUdt5VqzPuqXaP3lQJHsADsYXmHA+oONN2JQYzoKkpD+IXHVxGCDM6WzzPRNkZxNOJ5X1slBb/N
zJILo4R7WylZwFDOx8kZA2K+36Uvxwc4VZmwSxpNiU0BbIe+M/OzbCke8pvtU9EF7w40afuvIYs8
AXESCHoxToMqypkza4gy40V+y3QLu1y3Cgg6ITfa2l8/iqcMj8n5ezaKKL5SQLRvcKdRvj89xgHF
mLgMKCtfccK7EvNI1g6PTBlsu6X/OUjyAN/wfeca2zJgCEpFX3FmOFd+Ouu7tnLull6aThdwB+FI
frmWSoL7BaNeD/DPDxLHtxymW1vCQm35FW69jwArentgNRzmXVrg/wGFbNbbXSXQ0ApG8Ai6yOLg
ibD/v4KxNpQGMGPrYVwx+uc/6T1gQOeQkU0pypt8TzrXBS7DIruGzVtJ9eB3kY9FuB5lZkURx0CE
p6SM88YhmJEl0sICFBIGqNYmW9YfqwdeeZ2C6jk31f1kYnUhx3UHE64XgogtAkeSj/xA4MUG2EiU
afMkRy8+r0N6GYxqTm3to1CFqFXguGj9rOH7bc3xBPDL6oNLAa29RVOoXFSBjgOg5u+ndwqSbRPG
1ixhTa2GWnzDbPTZuvhs7yWu2DxMhE5XJjCa4PZ/gOH2fTfa23tUVBiIfq9lVNvhCDOo0JQo9kRF
FPuXY4LGrMTtntkD4hC+uThzyZMYImwYfkzJrsxzxi7Ht47n7yEbX5rSc/AuPheZ6eYb3ZIh5/IZ
HGavuyb4rUOPOVMg8Lhq5KyeOrSj/niRVkhPgRNG+MdybIlNDEygZMuNElX5Zy2dqw6eCUVTi2dW
WSxXThmYr5uu3cObybZYDlW8bpQ8xpkABZFIZ87vWXisaz/dU+GZkjVyds3mHI4sAxlcmRmzbllX
EdYc2rPkWXkdZ6W31XgPvv6gCTUfTPuBOhIZcje/iupVMtSrNFjAkvXM8eNc2+F9TgeUaEScIx3l
gtD/op+2lhYqXgCkI7FMQNK2d4Go9ZqprPxH/vPng3yWFSFQUrd0QcZZYCtEwHqSiDa/J5sotyyO
8wfei5loG//wo1xx0kRutJBbJOXqOmx1HpRRwwpfhC4AnBFosMvgo28/Efc/hIqslED4TPdsttib
TAAN3RrYWhg5fiYH/yJLm4W8yd/lW+mG3ANRstKXEPbIDKnSsoiu3mksjQUnC0iQF89pdggXFEMN
f4n1qLHFgeckFt/AElV/n6p++uOU+jkQEKpeZ3myfEHUIAK23ffpcaopaHid5IKFM2ZtoVVGFLsU
6FcGOIp95U+SRbMaeS5BZyUU5vWv08Ry7ETh8+3DDHizHoxwi6IbqvXFCszCLEObbVaaG/mNNFKr
pkYTUM9YeqhTQiG67uf2LEifFsJjx6YZXeVlF9Afrla9uDNUAmCvo4LJpekLxgq5C14TadLweEMf
yyLLDsJkq15mDNxLK69/hSv07YeBJJfrb8Bg9ktfkaL3VtkIPmrkXZ6TVgs7JmQ8GqJC8FeXrY3w
hZAgOhJuoRS6+YvqOdGzUHx+55iXXqRbLmYyILkrLAc12u1g7rMGB5YoDf5Q2i4PiIrp5C1ISKBY
Ry6Qq4eekvKu9abZysAB1xSlwIclImaGHyHdiBBq2T2eMR9XApgQ+HYu1iThHZtCs/I9D0goLKUp
gpHjfZhrMpeMn1vhlPJVdsosy7iDf6Uu79hL+rqCCeWH/YCqJXm5GgbXnaY/qh1wziZHpEeuvMvu
wDpPvP4X3qibFiNOJgwo4X2XN1swrLmDE6OWd8/PqNrcTh8cYhfq8Ua3hKR7jSHqNm8E2cTmCOW1
rZbkIFnIiKnA9n5oaZCjZnUGSh6+uP8S2pufgF9W89xZmcZwovnkS/YYb75HMngKs5jF/rf1Yw71
pB/ZdicuWg3SiJZF15r5G1HdXLKyiUkDbNf6uW+rZS+cEVkfJ2p90EeJ6jnDIES90o/CFq50ITlb
oec31KnF2MIWsPjMSs+SKEjA1cuIRVG/VQC3neOuHHGYGw66UF/E/srVnWsCaOU+ZIHO4l2Wxi+n
dRJxsB5s9vbTi0102w3HhXCUsJ9mokzhWJg4e+EWvCB3Bqb9acQXtS++bl/+DmDFgfzM6N8ZxpHM
xm1jdst1/i4gOQcAbZIFcoASSOvdqDdGV2ltKyXKW8BMVEFbCy6+Y+7241Iiv0z5orlvPLAGuBcs
TzKtteLvxFcI/D+82C/ywm1SoSgZ9c1sQCG5aOMwpl/8M1WgCJCjcqiBF12PxBHhYePsNstqAxjJ
RcpxRC2+M0+z0RoG6r6xRk5vSeSM4yYaReJWL8ltkAeIqhP5etJHDRW1LLGx6mFZ/gVrasjZwWKy
j6RadldpoText+UqYUjxmG+d7E3nWCxYdXpbvIXl2NYb/OtVTYhZA/8SV0fjVVCrGWo+/B5iRuPq
RWsML+Ml3jMxVBxFoRZmJc8j6vnQiHzT2Pp2bjSSJUTB5KivvVNxAMvJ7z0hEOU4VWOuhj9EHi7b
pgRqr7z2ImkCM7me8ReKyvu79BdjnavL9ks2LMa2mCnsXzLebhPV0Vr8FEcvf8oUQCVaygFvKzS/
RNjBTIbH07fGi1DT0iNcwFE+DtmQxfgpS6zpe9cdTpQBkstatmFUG/bvpEWyuYamROU05EM4gP/M
ILniDZ8uJMNT3/kt5WAk5eDtEocsG4Ql73VXYhhzoFByfVOgaHw3V7TSza5BDZ1pXzxovss3FAch
LZ6XppPQwkKekQsQsIYV+12m9rLpYOio1C4tUf9Y7r7RrHhYte3oapHQfPK4asYYQY9cEPwadCbz
MX8NXc8aZ3fEK3osf60jzrNZWaLN8SAFgn+sxSq0nVUOBIHh4ySFryWcbwydlZ5goEGds5aHkLWd
1RU5vo4FXgnMlDiW503eZI1D+/hsTIUqtkt7dRDfSrcoXpBfTPU392AsHA1tzcT8qccQmzOJLoVw
YjT2ZytB47Nde+0CgJI1ndST40R19HdYyft5QD65wCdAxkW7xcLb6OLMgeBksK1ldXnJTBuVqlby
upNHXOLRmNoUsTt+3dgyOxac8Qs1MmzhdiLciJE0l0YaCpBnfXrn2XnqYZyaTQ8Zk4fwcQLy0107
+3mfvmcMtqWK3wwKlp8hZZS9X+iyFo7SbEPf/PW0OKyvnfpVRVJqRgr77bPU5YdmNUm5XiaZ1vEX
e7dkaKyjKnKVkXKRTai7j0d50NUeQLwznzPjAw62BNbTizl0PxgCS6QAal9aQUVcRQEhVldd+I3C
ydD2G2Y9jJOB3qICr7CNNk8KaWilIKOLvD2SeUg9nGDwDPM4fhbz63CQ+AAFL1JWGQEvdktr50L3
z/a+wpuwreW6GLGuHWalQqqGk61m3SXZc9omHW8Va68KEa8cOYdcmdaHk/arg0765rrtWCsUymV6
1D+teZ3/kb/JfFtbpqa6CSU3DMzrXyibCcN6aMugY+Mqn4dfey2xrzBsA4MaAEylIuIRI/0ZuQS7
aB0rLBq9Pia5JvAQmfJB8bfQ6siIibL/6YwrZbJemIy7bgU5s5HD6C53M8RSsxBVMu7vMnB/AAa5
BIL3RdeGfxQbuyUtdNAbOjefSWpa0cHxmGSqjfrmBy99qtD2lKD+NqnZ4QBoZCTbHOU/4tS4OqtR
tdhNFXuc+Kr7v8GsVJk4iJsD7ZF2Od66lAdnT/UOcHXQKZm3lqmVtjA5K1mP2YBDhJLY6xhguWez
cOEHXdxSebE0lmdYLUUDyMUUfThAFTL7jYSd0XruqouaoOalj2iVSI3RCu+P6ltQcqn1r9lh2Gsn
yuCq8CtIn0tS5tt4BhpGrrQfMRZQHpkGOKyEgkjIIMsYtJR/HM5NXj6NKz9EI6WfUjMMQKjqkNcz
SlfD9fPrx48H3glRY3tTkqT7Gy5bO0LxdpQYIYW0C2Dw25QoUZl2KZdKnvXXes5BBGmdMktT5OcA
NrqGnw/CtAZAldSg9kgmskbOdBMsck8VxEY6AVjtHJ2JTEkAa0IYu6fOiL+YhTJZtgsZiJndkVh8
w2ooaNxWYdyIs9tHzkFdDfcXeqDtoLGHMp/FVZuk/n8ddT0yKJfuptkq6CHGQXB9Vtjvg9vDcN7X
H2lJVivAXbDkM0Li16bfgYB/KJIv1gM4gfl0EMl46rTfa7FgMsg7+/5Zd7LTWjIL1nILxSyfo7C6
CK9bCUAOHU5lS3k11oRkS5tKrw2i6PEWBlOHj1VE+zHKFBWD/G3EV7i2x258g5kYXIhh6E+T6gIG
pFhaHYZaqmfgA/P+9Q34mC309RW7gOrAanYLHbTNXBjiuFdRckZFvmLoUiS8g3YPUeqbWHRbVHgf
oearab++9GsYIvZE/5kNqkN5Wr3VC3foJ4UQO38kUMFMzvFW3sLx51llenz+AwYCLzrSrGrGN1KX
cRIGPG4jefukliN+it4MRSKD9tnsFVG0/pGB0Xn3hHI60p/Ra2YiI0gFTgUdpkxVbH+QvqH6dfC6
2RxaeUCHJtGiKhr3DTiv+F0GOl7FQfdGqI6HhWrp4Nch7doFi0aIc61q9G+LeCOLnGhDyEiKnYa3
w1O6F6msGyQSalZvhsinJWDCu1TsaglWZl83WT89sGG2z0HakUbJnvL59kz3JEkN4H2snbvzHPTL
TrXhbb3FPwjdNS+i88K+P4JwD9MvGu4bbEuotw3eyL6V6TjFJYgYtYCtWZpsUlB/+lkuolbz3ein
7U5uNGKgh6rOA+lMkKCyVMKkbNKTfmx0n100FSVj5/+AKOvvj0Hsxi+ilXIFqrlDDYJujeiFqzRp
I31lfgvoa+JAeZ0+fB/lLAtVfXljqD28YgjbFCxtBu/xOeJ/KLyF4EbNw7PEEuisw6lFONrBzFa4
uGclQY4N0bu1zh/+IINDLW+IFVjoZdEEqQz6pfr9KX9I3QP/tRSToI1wQBTDlyKaM6iwvOtuBblQ
bYBbaluDVnwtxSbbvaEwIxmcxAJ/l+Pmc3eVdqCQOsmM4oV7WLHfXQx703VDr5yRYDCFFYkeelI0
JZI3d5a7mlo42ceCVxvVmW6QHQplhyNNuVQrJuijRwnVPfFp8B5FcmvjdGmhiWpTd2iTRKq49+qx
c1aYJ1usDnofZc7zGG0W7O+coeJG4O+3ICfLdIU7perWbzw1GXHd2QiPJztpMdoCMIfEsF/aSIZI
/7hrV4Q00T1SPrdn1d+77MV8RzTWkoqU2KtSSGLAAriHGES6T/ebXe/S5tz2QPB302H+fCBg41KR
DvwMJw8nlvJlOPNzqJHMKxT5xFDO5iE9APdVipzSeRl+1OV9FoOnMts9mps3Sa7ecBnVWl/re1Fx
eZgJrvXsVKht5hntNW/b+xL/uFFp/Oajx9wr6kzHIVQNsFgPNBA3PyCoNQokjCeCzp7/Z+FKgpJY
7fjXSGXDGTqA2nxcfWh5g5MsP0dSwhBmYy6tkpV0o/rvtXi0mTsiBk8o44K00pyGfdJov36qYa5R
dWIysUgbAzyr0pbmBOeeU6Et7brKx4S2uT/ZgvB8HDZ8WMzNSlG6i/KUFS20ww6YEDvDRtI+qRHI
vleusE+wUh3gpELfciYEB0GJrB9rAGGxVCMpKnea/UdvWKBCRoItb0Z7Fswaj1LcDgCJBqwy9Ug9
Ao4C0XCGpDGPuYOyl4P9XCI71pKDnKCgt8Zo40qT4xkPFcmpd9NgdAX/FUienkCWUyj0WTScfIrf
9JnkB9pnCXynpZSGyHvZyQ4jHRYBcQkYzDUKhMipQEO3xSasVmcbZDnIfZJXfzxBYCskfQPL42NC
Hkwxp3wuwAnazkODQrdYlvuKUO1ljVg5NliQkh2FEN2h/B0V50u+/tVAHXksAhWp4zEYlK/NGKyU
oJEmZ7VfVCDB+XGqTaJQjZ93q3aV2ekt2PXIq+DEetH2//IT7i7/RwMcOsd6mHV7Q0/MCLFV0Von
KoPTKGKVLmAqtZgb0tkWClO52mH1I1PM1JtF+WBHBmIRxZ30ar+BkkEHdvd/U1B+QzePxKXeJobs
/OPtpLB1A7bz4ittsZrR0xBcH4G2Q018IMTPUChMJZwzv3VFFr6zjXuUWylp5BjBiWX/w9A7aFUx
0gW5gElMD+EB3dYIfUTcArZeIv13rneQQg64MYWhqukzUFjh8rvqNFOequzDCeWAWSX0NEcmY9cJ
bPByuVISdpMR5ElM8SK620cgl9oRWS7FC3NZH7oS0seuJJWxN9QOFE/o9eTViJTnXkqRC1vT3dnS
Ie66nxnsIZCD3fN3ks2QFBkaBh793wQN0AJYiwlLNeHUumMfXWXfGE5bNcCMD35+aV1VYXUtAxNa
hz4ml6OIVaUSCyaYoSnneaLbVepojuWKYbtj1myYMKAvxG5jwM1F7YnAhViy4lpxwjQh6a3En+xQ
/RVGTn9Ehdk474iNREkCUe4UPmsDvDX1nIlYgS6eRR42TfCMbf7CCj8XWSFe1ij8XfZpXPu+9Xnm
RljLf/9j8RCPRaCxSN6XthqGYSYiEf9244yCNmiWMdWCU1LCGJn9ZO+IZwYr59h4c5LFpH7QLXcg
4+pWhOtBXJhricJvwnVkA/qWIYoY+TkvtBVtibAQcTT9Io/DHSUzmnxjiGz83IGfpXycOPMdHk7S
RdKSTnOjDIszsauxUa+sDHBS16cH//xa6TsUQk1b34TH1tPD63/cFs+eLOmkRHQdBwu8NWyHZkuQ
t+kbY+iyhV8/f0eh+LnpxDpNwB1gb+lTxmEFnaJyWgWQ76XegZdqilUFaXwnvhGFKUMQ1N8awT7K
CJOuDJtbs25PSjatNwHzGbVbpL8FVzhzUnohIG+Y/WgWi53sy9L/fW5lPL5EgkfC3yH/O+4Ca62D
MAIvna3A3UARIf0AW9Qkoy/985Eej6DkJ2J40+LyguATDP4j/r/OVFOcMjqtfS06ETugK23FjOb4
pYXhA0SyYw3bPz8a1AEQ3KDJX/STob3HyDs5q7d2YzWdyiRDOkgpG+GU3tp7f6kTKQZBY/YnLoub
q+diEnLy62+7vwUkKn7tnoSUfEIBEYe/m4Kk7T6A5wiaIyWK7TtqYJrKHzn+vTnOS4/i/eUbG9VL
237OBIaMijhqLT6nKyhN+EmNMAQKzZObDV3SuRGKNo8ps3CvERCFmeMz0zvW3m/tcSMLqHPU70eu
7Yt8K/ZnbnXHESQ75YZY4DfdEDtdvXkblSChK6PB0bOV/I+nm4CHYo31CS3gAHqitP2Tw64HJf5j
A5VZ7qsoCaqIOhY3Kq3QM4TZnPOuLpPuLOvNIhtwSP11Am5iErnyX38GVQNyS+mw3RPVD2Yl8HiA
PgVu8bmL+5i7Smmeg0JPBBhcQWlkUYk2BP4BwoP04N8QJk5Koekjxeu1MHmYEQgAlUh7LZNVXlyS
BvIMDzTlM6PkiVQ+Cbs5x2K4bP1kz3ixWEP3v1979FBBrDG2DWuCwy+LoLH1KMURVPXIzbWQjzrd
ghu8jXKXplNDm6UAXEfeiPXIoedyZ7u1V0MQ4+1OxbB0EPFwM8xIoAmHnCIdTe2yIO5s6TJ+JB4k
0IekFiLlqOA0ClVHPdoAbv3iT4C/kVV2D4fF0CmttYrNACeGCXHz+eJfieZWSvIT3jsj9k5+i5d7
2yO4rIuYmlPhUQasJmW5ug5XFfgur62134/yzXVipyNXuTze3lUMIhFoJ3ac2/IX6sIF2/2QPNkp
qqnHJNeazLKm74M+biV6rBNOJP6E/2O3YXCf4gU0YPQHvE3JJYGXpGQOR6egA9xs0R4VJvsI8An5
RdByWhHg4/tPsmQYAPyaZAhPYbVWEBT7Mx0rDbGjoRB9MHkq2UwI92UQOiiRz7Blqvr/WaFZny1v
1sd+6sPKrCUA3QxXZhlDlLErTpp7bB371fqTueIa6NE8107b/0kU7lajgApUvXfTpmpl1Y2fyvT4
93kFxK7g+uDgs+zcYW1hrXIrKUuQMoFZSggwFFdRL3ZL5wrLY/lJghnaZonnTk0nVmLxrfZ5ELoJ
a/cmGC5V5Pz7VKaA9VKa4ar6MBBPtqckTElz4Gy8m9e+9OcfZgmOwuJxXghpMkGdDhGHCq/mOzLg
nJ0gJQVMdK6vHXVfcjyWO1ZCW9NQ7yL+aPaDk9ydNUe4NwBSL4cx/QYXzMxUtn6BIWcyQCH6iA2R
9WyqCu7VCWYTT2w6HCaIBxZARSyjd2esdy8cEln+brs82hn78s/u8ekFxerH8V+2z0X+Qis2TYUM
Z0OX6UWhXz7xpNx0JkaqRW53ZxY0g/fh1y4evdH9czNVeOJmNIobN1emoLwlw9WHwPhbSWMaHoCE
Ww8ONYdEMbO7wE/Ok0lL22dMjmWUCpzcf7gY9xV0D4NQ2R1BqhM/XAG9SYL3KIVQDK+GJNKjcLpf
+ThdMEBYKDB4D5t1Z4+DhJmQ2vWQMZ4cjAN9GXhx9rz+DW0I6L4ZV63VYbsnYV6oh7nlVOGXiVq9
b05MFbXFagU0C+jfGIvh4w3OObMjqfN+p1gWGfaYeP40NKJ0wTp/iirMAPcpiN/VjRyqWNNOGrnZ
OrFeUxwACx2o3lgt5/S0XmZyxQmjHAw/WKyxy5mFp4cMaV0yi540Cafc6BlxCOkpErODPBwUkhqR
lERcLe8FSz7nXHUgR5AlDMtmWqrf4JvIS/9aL5wRy/8bNq1hceCp9VybItttfhov56yBHmQlnKBQ
dHadc2M5qKCy7X8w2v+yA7enbki0DAKgy0O4hvjQFtPh4JWSeEhAGdDUjVF3SY/F+1b52fUR3k1P
SeTr8xCwaZTCmewfPYGMg5IAV5SApd9yYQTWhIB5/dtiwyD/nU9phGHY+uMFnwG0yRu4O2qFyDR3
xTnsfmmnZRblNwMKoIDTar962FoP8jbQhVQiK9kaHLLlxdmOA+2TH35TAuYGjBiqWtoPiRPlU+vZ
jSuN2k6pick6DIrHYd9pc6fT5WF3HvYCjMHA0PPwG7d2FoOPYwh+/jrPleCM4Eq/NQCFFCLR31rW
LyTzRS48AFYj3jscezF9HB0SPMV7iblYjtwO94QhZr/Tr8ZT674swf0KzH/db68WPxAc24PTMhfA
jFJgtBjQ1HQ6xSSCgWCwIGpipG6c9xzHTWhA0uNe/y5hq7b12HAl09c5JBFKea8yGboIA2SPSB94
yt//TpcvhuWE7s74cLyS2gkw8oyNz5ZYRF0dXjT2byESZ7aFXroU/IAYhoyF3GUg0Xc/bJHOfUMm
EIxZ7NlM7Rcwasz7CkGlIh053SC2P1sml6kW64TiLSi4gW7qnWHMps1YWvTdJH2dWO4vs1F4lKxk
/8vD5lgieZNVmGgTMFl33dXiELXN0zvavJYK6UIKS7FW12HRQaw/4571dOKtVWAAJ+QRmqCah0ml
q+M9QF47RLWz0Vw1bwai5wrw2jNM1fwMigLHCKCdfsPk31/NzPeLBZvG/ZEAtMFBnAWMOmDt9pgX
BhIbwVB7QfSy1uffZo9NzWWy9zbSy/STcdBkP0wIO0lTVB15/x71hJwJigAAUO8iOL1IvQXwBOGR
CyI93YMxbdrpApNNWXZ1XEc1p0DJUKpqGDpGdj8jtpwX46I0DhgRFnHLm2bUaLlJc3YDSMn545qB
V5SKdsThuzKmKtYkDZbScNxmLChd7hC50MR9YStDWymB0bXqp04XrrPZ8V8+58mIBZiJo68hkZJX
YGT9llXraSkIR+8snpAT9nTzq42ziw50fZCdhB/S7dOcqUBP0/LA2HD2cLGZSvpg2gEQnRIuzXDT
ddojOaHUz2rBapRGyib1nSR/+cLcn9pCkAAtqp779NCOUxh0ZQ1xfItGhxlEKZsiwWSfwZhyUc89
ZSHlBrHHUHQwIh7Y+bOXjfWXCX4FqeSYxAKC1zSMZI7YyX6qJf1gNRHq1YxZbudwdasAZRiynKp+
gICz2A/D9qZRGX9GjE5jZJvkRH3jNcb5qS80/vRR1rOVZzf/qhOY3a3uwgOKkhhlAIXmAbts4C/Z
WaDcz8i4dS5XEqIaCHTyd7zGB3IvYDDZXDGit4qjgi623bL61cH/hpPRJb0Ok3HaMN/TbfCO8L+0
57gFXBjjVjPTftJU1kNpemx9kRpefYc5Wo2IUqNI+eMaa/ZAotzs8XarR/VKZb70EDMEnmXHsGFh
hAp3UwtNi6ZF8Vb3ABWRHNAUXzoAO6eSqZUOGA1XzonrNTUUid3YXJ8cGM4i5bXOCijpAk2z1HO9
b/WFgqDsZL0TsDuBrSBHbdyNI446VRF0lMQ702ML0RRU39apR4/vHwAjxNvKKW9DU5TC+2Qlq73V
fTQOJGGn/0K2Lphe/pYWZjkPPuhUPjZK+aaW595lx2+peGjxzHRyXtJ84R55MX3UFP3Iep8oAQjD
tye0v43F9kegXi0hyeibUJiByCBMJFF5N0q4ZPM647frVlpoabmFvxbxw+8I3YJXA4pRsqj2JrcE
4mbhZL+cZVl6UrERAVrXPMtxN98lNVb4c79w73oKk/KpwPXmKeX6lo+vgpFKQ2amy/YenI1tdP0r
XX+TPj6ylrFEljEXk5a/6tEDi3jWaTiOxvWqQpX0RFIMCfpRZbB4GT71YCuCR1DiVmXJTZVkhQsw
refAuJVa6/7VrcBebftJkYVKmHbEbqwmpXDuCj/VFSEmqYqSG9v9OExU6V2RbVdUydceT0eui711
HB3D3U87bVTD9YO8nlA9DXBdqWZBJh0n1bTFCq8empeUHOyE4KHBiemVq759CBxbUkbY2ceGbC/x
EWxGRYNZN2Jsbr0sdEglYYsp6+tjq9VoEWq4P/zFgagFAS6BUxw5X0DWll1IgRR6cdEuOjV6I8Ba
LJUffvthfVO7lfG3YCU1zpC8hcwMdy0ic631Ona+enw1wNNlDvA0Yd1WIEwsWthM1W63er8sKzJT
ibsIFnGu7mYzx6ZYWRSgWVnGCmLQRrdO3E3rumUUuRHYYBxxwzCW4lVWZXh6+4BrqfrCX8+eT+dU
cLOx2jzoyEvwqQi/tU5UpUcvWTQO/sIlwyAYyovMT8C6rvfIamxf0ZXNfGFYIIluTtj4dWeK9nmP
jDbTFRTVoZQo65iI/cQTQJY+gZ6fbIsq3xSEWEQg3O2JX8jmt1XDdfqrHmjrxPOTRfN9qqvtSBvP
YsVwiTCQtZbPlsJMIFYhoGe39g1m3MXMI8R13ppMu7Lm/y//x4QeJcPeLstNpj7R/c82gZZWTy18
klU2jx1zAPBoqxBsrSZ75bF0eGLz60jlhcmNGDU1lvqK6HAkSnlZ8L7fcJHrrWdKvC6MZjOA0T1U
6DXVKI9bcYshJX5+zo66L3Pw4/yktcK93270r4fESRwH7T85ExCvWgGhk/+BMBAZs01jQemrw+LZ
2XJO6w6M1c2CldtSvZtM2p5qr4KY/gWjw5E8jXO9EZx6MLV8brgPKMwl8Sec2vbFIOuco+HiI2oG
L1O6r9iJMn4C3bP3zddQy5ky6WoouESaSVDgsENwa5nzIqKqL2izxwrR59zedixl4sSoF3pUQ9W6
xIl7HT0c9AmU6xdQYkfL+CD5NXnNxqlhSrl4ku+h2xOqvYQ4QELgumKlaejM+6VrNSQNrOvJCjWd
41l3Y0qgnhnRHXwQBScCGYhMfrBwcEopx1+MwC6nNEdV1CIKwtfNaLSGBBq3AqhN72tezq/7PsUR
H7f8mq/EWz3GaqhnMTJ93+5Wldi2DfJWtfPHfjLkA8aAa7sVwxtQoxwO0N76gM/dPmMAkoSdVumn
0LSv7UMTYGO54gxaHAFthqnlUd6eKk91MdF4g7YZWJf+RskNtQ2gsfsYH2m5u595TPNL/wL1owlA
LOi4254Df/9VexyxbmQYBRdCUcABzcf9ygqNgvpxkCd79aIVi7U5yxGvui1ws5YXkeYjGeOKClEA
mVbLm0pqlVlYdizMPbCSnBOa7yYls6lZtZxWAbIOVd5ZXGBdn1mLZpajRnZ7eo3KMb8ONQXry2wF
Xps7W1LW+XWH7CKbpBc2esQ4g4qXpD7jLXgB8KS13KZnDgVaz2PVAW2nSwayAiFdgd/2c5R30RN8
LYGkNcY8sl6EL1HgxfUASuc5Wiqo7Q310CeDTxndRqCDz6pCrSUg+sBOwcx9/VlfD+6/Ma5PNEPJ
iMOprmastbup/8gyTB5gPFz1o8yTPH7ZUJWjfhiycpUr/vfjUobb/7IwpHzxzPkCAQcl8uaJ6R3y
80maGqzO0UfuUpfw1iKgPcKObdAF+RmHEjHar8UuzyJACX3G31hrRa8SI7BJhTCWfVSFfh8sNJmi
SYhbiRAQgxLcDr/deke5u6y/4MvBQBxSfIVmzIZGg0wNp0l/OuFGIQ4ttQgLp8qewVwbll80+Rmo
MX/Gp3UmxBdrEk8mY5/jbi8k/UHtil7CqJXj5d4tW/bEs6Sf8fw+x/B7NOCzRBT5wgtHicbJZkV+
FUOEqkiZz/JtRuWXBUZVOIkJNGvDBufjHRBUqE2ixigFwfxxuNFpabGCyNHNy4feY7MXDcQOweLq
ABz6H8+j6oGx3SvM7Dmi95mzK1iUHPTDZ4GNOtLu76oETF8mmW+nW+boSCjPutJ3njDYTrOYu6Dk
a2Sh8uUcQb8VIZpAU9kK285xwX6rIJu2g8SqG7YbzixlwjWYQOWAXRiGTiUM+0LNnzO/IClZyQ8A
JNeQR8vkaT8hB2yU270dO4Nxcr2tSefqGu3Q82X36GZho8Od+irGP4g3orsTviE4Rz7SeJtKsUZs
oFFjpzrNtcS8gIcxU6QLlL9/t/8zLClp+XFrXSOVHtBvwM0XjhLfb/NMGoyPVk3j6blUeWAgzKaz
FQtf12L8muIEMxwbWA+De9XF2yb+GBG2Z/CKi+IiXAlN3aBMLir0LVUA36r4qY8Qa2k09cwPM+j1
s/9971Fjt6oMBq7vyaZ5z6lHZvxHFY2gT+tG1bM95fYTWeeMq83BGsui4vNL5R/DeB0OTNwsXUyx
+pV2ujELXuzsPTS+eFsT5t/4/CDOu9r7GA0tp+6N0br3Zxx1QpzG9zHN1APQpuk2o04v5F+uyuaU
7AzsAYTcpnNTZ8bZ3I76tgvWN8tcAUbrSPs1B/+NUc3V08akAqetZkHEUrar+/CYYVsosQOTPpAh
J3AnRblwVyIKoLjs5zKGfFV7cJfqfrK3KE/jea7Xv2w39h20TBBtD1hvMHKS0K77osFYE5J7zQ+E
EpISn+7XMMjBC9dd/Sy9r2lPYGldBKR0CmPhti9BwuJSxJLz3CPB7u5TZIj74lRGDUNgKkzJO48P
qVMbaZMZeGRKQ45WCOQiE8/WuCO4sedjHkySneDBmyF4JHURWs+/c5bL4gcbYZJigpeAu1p+MQCM
h+FDb04JGl4/e5hz2dABju2JiteWMUlHGl9uDC+fhBdG1aSv+KctxDfkzD0cmdhrOcsJMAFjKE2W
40qhU1cqNvAlTSrQSbQbzUNKVTCbhjpvcoD/HaZiPRzPmV6IqcULk5z1ADJJoQBfGkazUiPjiNVU
nJO+dbUUZgYe//vTEFZefOeMkCk4w6UCrwfHFiLZoQSB2MeDqOJe4lNoXAqvW3rGhYCn7DPmYoo4
ce4HS6oVbq34N/rrwuZKZ0GGsXsAJkG7tyt6JfNyaH5WVnibqmWjv11aah1LboZoG4mZ+q5IFyLF
zls4fP57+GgANuMZIGfCRZ6NtL1zz7dNgi3331+2oMvJ5hLhAP06F2wDTKP+to+MbY1CAwKCfFDq
CY9fjsXDNB0e3a3H1tL/7kn7++Pk+m5gpLH7L0xp88iiK/D9D27Zaf0M55J+FLk6/uuwmFfRiR+q
5CJ9zN7IgpHAmvzf6/J9BTrxLWgH8h6/sAqXkTxKTx6SPdwe5CJ9BckfaD5svDJpSBFIMPPZw/Bk
IgfAN1vdBMAzYT059xfwb5tW5h84UEgurqxsc37yTYlDFcGv/7EZtXsFNZ3Z0gAgaAyp8Bd9urx2
2Fj3yI1Mxk0t/XgvxZRdYVNRNz0cSNBHKwWdi5Y2u1YftUHGfL1/vUOoZWH3agBfp2ZPgAPUt9sW
F4hqYtfgxqT7ClW1o5mlXUJOFKMDz8+kankjrARG0Q8dddjE6yLXMsgNDA9DtgLO4f6R6VoHMB9K
yUEUXHzxoPEWjVrVZqTDVjy0IrS3UR5MloWwrqKlY0X4i7wGV5VT9yb6+JVJan2ak8B+1HcSuVWo
wAWo3cgMJpn/ALC23KNNCZ1cTZq75CgDgknezyZDods62QGzJMTALviOWueGe+i/xV5sOUp7gYMp
+sw3PP//xAtOVT4KQj6MtLy33JIcxB7JPEdC0jFw3K8LLt2a0bNE0O51YxGa7RDz+RP5rxBmccXb
FIrYn5lHAVQbzgLS1yivdmaYO7lDk8LNyJ59f+HZYt8mp3/adou+ofJoh6MPfFMbRojsco8O25iS
fSwu2j2UDhrjf0M90AJu88YVvsWZ6CrYh0+e9zBXd/5VP4reAATQBQMWwzMBTLk4tTqxSNM5tDUs
uBdyR8DsMPVRaEFCXQOQEcqRV+8wG8Mimwb7aDIYz2MvgqwFQdAyNO+XJX2MBHmvvk/cYmhTFF30
gb/nBnVuRhwNTpgoWSB1HFgxVNlEk8j1ZQd6ffg6jeVjqjShpAdEps3jQtbwg1SDQv8jwKxBDd+B
niKJt1yQTcrKiVYgI62muuVkAHHRbeaQgJhE2omq7273bS6SfhspQSxWN+QPra0KGzdLEwmKAjeA
YVcGkQLOh7pRCpBJHHK0Isxk2dbLaX8sxx20ETifdNh8HaUPGbC1vk3qP2tI2lHU5/S8apagTDj4
z8nW0wXImBpeZ9l59STyzieCZaQq2ZTNBZ+TKtjsBx/Yot3TR1PxHEpGrutQwR4lXrwjwDBg8LWf
fZzDVEX8U+sDBW2fRnV43KBtfCdEBkpE8wHgitqLNK/BMledmlKywWvc83zaE8TYbOIiryIn9x+2
Xaqf1ipZstK0jB4gJzUpq1kJzCGWHPQHqAibDQggibyn2sCY2RvCxDxrkeTGAtGRf8/z/yy/yp2g
hjMTdaBb6jVK6nH0VdQu5dx00Or+NFf8wmJLvtOJGUTxRMkvXKNI+1taTuFMU7ybQnGF9m3iwLEk
HAjiP0MTO0ZS5aiuM0YoQjFbLHN5TSkQmr9oUDcOESyKzSddt1zTic271mxPYK0xN8cKWzq4hGm+
8nf0Ux2t5FUcRJBKwwO7mEd8l52IKLm0M7xmG1KaX4uxP6GiWX1EUfosrUDtANmOCM4icS7sODyL
Oq5t0WBeQhB5GGrATyOboAKeAXh5gdjv1HlpwhlTBYWaUhWEhrSjAVgE5K5QpA1q9VLOl0XD7/un
beHQIX63n7xtWTxp1RzKFI2UqZNfeVs3SFl1CPOd0JeH2nWyO1kg8G82h1Qr7yn/qzg0oXePhazH
sMDIuzcWLJz6j5S/ktKIyoziFD3uD03Eee2ygb62Oh7td0e/KGE8m+v/J19pXlsNnwTCMIU6TV48
w6utNxxuggDdQhm/OMEXyJ5+h1ZCwWDWk3IOhGUFSWGZRnMwmTtHmqtsF9VZ1STKUy/km0Ubi0XX
8VJkL8ZYKE3OQOHe13v+A2Yka5SH0g6Xh+QBw6n6hPFKdcQfmuNDziq6vTe7Ht4WnkrFXgQjI4mL
5R/18xJUwiC6bq5KH1PEY6oCRfbpGFEd7RelqFWv5jrlB5eX508xqah6dyernORViGlMV81KvVik
E4cOCXgTobUGlmCERPNND0EPDzmVXf8KTKRpuEd3mfeEZ5Q7Q4kV6XsN3glb27aFQlp9IYpkjlCv
vuKfBPBydnaCpQAOY5W95eBJ4HHPoz3/1QIcwnAblESqWn1vp6S4i1kXYuh5lC3+8IupVXL1TnQG
l1x6p2iXFKRaiVAs4HdKOVa79Rq2fSnqtHVVqwF0h9efcPubuC8bDBimUbtdRJUkGn1rYEsmIHeb
aJPwastbneBTbgDcKH76kh5Zxv/4acawh+55BWLM0oy2jpQRUVpP9nK3gS0zJiA0/ZaaYY5V/FJq
sJjODI1XmP6ZyMwuHJnE1Dn24bJH9ZCPe49nGKdGjo+DK8chUoEpuMoVt8cBonTIkaQRC/Vhs3ex
9BbmsPElwuG6KLXfqf9NMUGTVxv7sSe97DBnVvSWbS4i+7+BGVGFh51Dhrfmf3Z6wrD+c54o3vP0
1F+zodw+fvRkopwJU8dk+yA3RKIn/rjx+5jOhiQTOSr16hrnLeAnLp7IBd8kUUr1odMd+K9V+PgS
A1FwaDoVshZyk7rDwojbwqtCKhMFlZ4cDXOxRj5d2jlGCjR5IppTghIWDeSFeDSIkMHiwLQiJ3/v
Gt4i+vqrZTUku/qM1PFYw532D7tD9bhD/fdj1Br6nIkF9YLn4WeTB+gXUwFox664lh6i0GjU50Vh
pcfr+CuahrJU/UAf9MHPRb6f2RnAD22HY3kZbRFpwGG54SdHNkGc9y6gzYhx74hYZ0OoZcY7gOoM
5WeCT6hAgD7IFvK96L4+EXLxwJk5y/QpKDDuxg2VbWJXw2paHeCgpPhHz61xrTmAkExgMcwo0XcJ
Gpbn1DuhH6S3oAZh5MsKa2JDYZnxAo8WqcKJTM1YiICqmIcjET/DgcRMVNQn/sNfFU8vcR1Ia/7x
e2oDwNueskzKe9e35VdyrqfoM8AZHwThh289Lszn8S8LDW46RxQ5LldzPFYkXN+j/e9jC443z4SU
J8+UzHabMxIxn2SodUihNQ/xLOlaMnNdgDeMrJ1piUV5tnTZmdWGnqHgJUuaeuaIAIQhmOEgzpPo
zAyR78YuzJIQniWfR1Gi+vFukb8UcYMOAU5O4Jps/9m0yYEgZZcTe3OySt+e/tWpDQHqBG3Ld25o
LYmMbzu8ag0AViO7v1Rzbwips4OOYpn2323ppsn3pItt9KdZyIG+z9v8cHbql9oFS+crEy5OQLnp
CHoMWHJmaxgDr2ygS0g8EeghOGrAyvcaoAEhtbwmT7qPQ/6VuBWzJNhtbe5dCsnrkTIF9SZslad4
K13Y6lKOSgdGRNyq5/V9asBTfrXX4YZtzj8nHBwLYMKMhGqtZsc/gHo1lhoI82OnsV6CMgFN/TYy
CjG9JTnbpz2JaFbZScGCXiQkI3lEJwQvsICCmUHyIz+OXFE9OtAZjq5BmCSJcz6aNgT1ZX3SQBum
yjvvxnBmoRDS6DgEikPxflgbZyoERanMwi91BIHx619mWOIG0OcXnsylNoapb0nOXGsODLp2nbV0
RCUvb6dRUUrJIHJg1vv1nGP+jDDfYS77MP+V3cU8dGTEMHl0fPgaohhWJzzdZXu8QPHne+6McMXC
FUeNZdbgKNMW2AQEuZE8fJuqsEQ12kJD80mz9OQTzreJ6khwiT3ZRgL+pzHLeQ/j5iEHPlDTkuE5
GoD06iXwr9nhMOt2yEf0lNOu+f5ncsWGhDPfO3m1yBa6dq0KZwdQ1O02bmxXFMWDfiK2v1QLM6QP
j9eX0VZIAhfOk3dohSFv9+CJrh9ePgK/yeM83Uz3Sw1KM6U2cTE+gDciUvkNcXVVs8XPnczaY4Iq
qcfpSWYEkl9wY/iNksd6NBUpQXWRh4uleF2U5E1zzKsNeMN+kXKavZEGK42M9tAVWNNhtZ2Te9xD
m95kESuAj7ya1ldUfG/7x9I6GcauB+5FeBhPOAiHsUaoHDIMWHdosjwThDpMzu4ib3hJn4YvzOli
aEjyGbt/sPwhYkXhe5txqx94ttbyN4m1v8uF+LTC1rEDSxVNBw4lw+qAu2uI6q96qc+2WoWIK2Bp
/42NuRqOZ5Chq2Z4Jp3qr58YLG3qciOXuQU9f5q0tPd2XY1dywV0U0bGJ9vzvvRMQftVqpzJosWR
fUfHgV8q7tANWSJUhab3l8yma9jkxbBZjhYGb5WlK2pT5aadM32pz1x/IpDja/Q7t8oy5kwpq5nq
NO+NvxQNiFpoeVJz7M1BP+q7bu5m7/vjBJkiZ7kVVCABubd1iyoMO87YgOSkIa4WmFbw/jzIjsJV
w9RxRXp0ug6FrOEotDgqqqF4dJ9TpseXOVRjABv6qrLC5Ea4KZI6NvcUSCUcSUvOHnmMe1HXIw0E
WyFavPYSQkRN0UN275sRBoT4AxfCXySbEh5Q+CzXYRoYt8IgXq8l+SW27BLFKhEJnF8xdrBM/kbk
IognKb+YU4j1TZe/PiO5EWtkFq5skW1HB7D1xsY9i634yODv+2vRoi7XMXwMaSNFsEejxnyo9AWi
i0Ccp+hJ3qlXcrbmd3ZP8h9rZ6j0yXJzAza88GTwbueK84FxVYwgMvpWUNMSQlKxDsRQkym+WN5m
l8pp7mWb04H33SQFFiTVFfr8kLtFghg8F6/uAQt8SAz4fVzCrHYnuVJQpjt41I9GykDbFerjp7Cn
bHnPEVH9yx8JHJKsYGJhbaARng9XHZBO8N96R7LihivaSP7raHlkT/Jk3iqXke3X9CvWjLD38cvD
Uia+KHfgRNSn3ZH92vqkZoIDGxD2ENQTeODxIllsm4heAIgj+BV+kj66PJIyoB+iIWWND+oPW9jb
kDYwfF4WQw1DNGJmj8BZ5zJi3N5FGCrBKo7cxSyvcjq4JDDdiUBc0LkJ6rFOmF+ODrVQa2Xi6PQJ
CzCMHK9y9EITWA+Qak2ROPcHYpd8mnye0E1p87JaPUAijSglTPY0kel+FweHBm/tJZ2R/dckHN2U
2Y4aBf/51gqRD+l6XIeCHhBV+gTWyCXCBljpJfD1uWnaQArh1nPkOlY6njXXAfYH73P9Cgj/F7xa
bV1JLNg5VAQRK0BNvih7BvfWTXcxzNzFOPPoYiWOEH/gNqxdE4+PxNm3R25hKcEAL7dLRuSWPxI4
ygVB3IJj/fBwcSLAYPx4K9X0xBJGjHq00bWQC7dwD1St5RPvwZCcpTvReD2Mp8+JNA3rVPBTjnjB
sB3z9becYFBMxd9f0RA696Wm7sPcLlfbJNl2CQlHkhkFnld6ReJvy5uMEIXtbu/k4v+M/+T2vv3q
x1AOlPkdjlF/ihzG0a17rVjP96maHCddHYxo97L01kC3WG+z897No1lqVW1vYK4CkRsj/0AM4yBM
qpbpdxYfPEmsDd6P+SQHx6nLAXy9F6sNDTrwIm/PU3s9GhAnh9bdMnDE/qr1hPCi8Pm0REFUZGEV
MPAuC0sbu8/eIOHxHI7MpYx00oaQZpN1+XixElxO9Bvt/llgK2qAxuwAB2ogjd5TApox7i80yQgG
DXMtE5LTLWPJScmqWq454X545HtoNoUjxLKkEXYFbSsFCenSFjLxUhc/AQSD+SgCSXCo5moKY9rm
8cNwU8o3acc9u+EbM1FnpJgCjodyZpE9O82q7qmh9G6qFq9ZgPf4fXbxi+2b3BubAwaNcbp1RHi7
zijtFqkgTivxs8QPDdI8vd8napgYwBuV9+1uY6RBE3gbVOwKxlZxloBus4SN8bFQuDYh+URW244+
j8n93klYftCY5mOx4JZZAj9w0vI3/eieWzvI0GUlpjMJABfQCqNXqIoqLcZIqFSlGAbDICpkwzif
m7cT8+kHLciB4w/nZ2haG9D4tE7nNzY2/IaZDKtKFnfXT+8x1dQb6trXVSpvzBk7/ietYHYp+grj
uBsJ8FORAVFh2vE4cXgX14dENXoU4XZm6O54nFhBT+YyZ9f6ZEQ9UrLBA2vVW/ZC3zz1GGs5bVkm
zE2YOQa9KE255+5eZDuNWRecPCJ1H+ZpT1bGLjzFJgkk9xc1+jeNe76l92I6hOri0B2ltu5KP0vU
xtrGQuaO6ZsP9gKlW7zK8X+IllYPpWty+JEfgMtwkEt56hxmWCw3nKy9zRlUOUH9trwl/ELXbmWW
zLXkriOtpyTkmx9l7AX1hnb7M9GpYIUCE460NPWYrK7zsVWcpayHsMtLsB7epRkgd3QTCERxFNaZ
IBa74NkACWXE8MlgmOD3bEDjKep5ohL2QGugA4sfY9FrUpf5nrMpj51he6+WsOadkgG+YlJ++2dQ
PV3apA5Ndrgv9ZZ458gk+Vgq6GsxRgtfk11I9qNojnfuQiiDhFEZu+GnyB+Q8jm9Rf3V75Wg9yFc
zeusM67tT8C9j5entNaEuhRRQ0oZGDmKeCRhnniXxAb4d2592vu1tX1Bg8awWn6XXAP5U3qYb3/w
CKskHzoZwN++gTip4Vm4iucriXtWeDEnE03CmU2uXZnTgselIrcnseeIqn0XmGFRj/0+ftxDM91K
7YGQLVC7+/9HA6+xXTLn4QYoy19TP+zqjop3IhiuiEtjmF9oCT1DlNF76vhmxsH/avij5JvwpuSd
pa7tkqvEaU3xmxXKZNkxJamEcSwLrNNruvnvmkTK/zoQajm3qG/TTOSN5WgBKYO71vJxGxmW7N2N
BhMWEizQuO9pqCAQig5P/f+BRGcWzETMe78tReEGUFV3dYRAny4CdP99JUTT29XnQ28MDgARUmh0
0PG677sx79HqobGpt27EkGeO6nSo24cDdV0s2cPpsDDY6tTbs0RQ+TDakAeUN4KZn4wdwQRSMIPW
pzrquuwbHDKVu5VKaVI2f4siNl0XxaOwAIzTcrhFzsvY0yVD5TQOFbu7v+TlNNrxEOhem7HK2RYv
pwshAhYqc9duS4hGwR+7YigjXYPgyPojAWVkhP4sXMyn655Fl5lx4+kHNkae7SsdmlijU62rLwDG
Sx1Z5agEFOjFbh2RANQLKitHll7nyhBqktNQjwZUuU3HNsP96wN10FylTPUbiCws7Ozm4xog90Wf
GYAD0vECIsWVJV6EprzRpCM9LoXbEOS4v0f5AiCw3kXnrvbWyc0ZT1M5BmuO6uvxNYP/v/7ha21b
rG1ta+n28Ru2LnkHNfsJBJ8X24rflSl+/ICfl7nhOWtslv5QV6Fc3HRFKTzoaXJDBsm98UKJM3d6
JF7g46z2C1WynK4dnVpp5WZIFyM7+dA626NQUaU17M3uaWciswsVtlvGCcf2AXJPZpiN3H+iAw62
FkxophM1iiW/dVJtxV4x6jyikbhgypG2CgEnMz0Y9YHP3cDu/NujDM6imL92YW9vsT3fe83wuC1m
W6mKYg24wWr4S3gENh9xZfogR7BP9tppNUF6waG83Kua7+66zxPZr2CZe5bgMylOSc2uyt41vGHx
Z6QMK/mGNE75oO4sElZHpcp1y8UKk5e86JfRyI4tWh0cSBbbiGEAhS7Fwq8NghQJd/gz/D/nAWWH
eISaZJswepVZB4nAun/XVZCsRTUCz6QxqI45NlL/fY7KIZGrbking4XxUkbQ+k+WH0oRHd9Kk/2D
7NppaI8RVJWY/iDDNKbWFVEqbk/Y8jxTA4nVICqHHNQ/jlVpVcu6CxLijs+ZhXRDpxYfHOzK1kWB
Q89WAs9h5qMUsUgKqNEdTFPZASjdVy1TjmRxpcAiAwfAm14HnA0399jpQ8AUILmVXgixWv2IgCM1
k6zQbM74X883cx+wPTK85b3kWp9UDcCovT70uJFAnIlhh4uBtU4EYkBRF7mJY2GJ1VlN8XAWIybS
V6DslOgiCefayd0vcKt6LqYt5x3O125Ujtpz9jvnucs9bn2O03HgxgaSUDQ0qCUC4oR6Vi48GG2g
fXeIAmIYTD0FtO9rFCSDsa42HRECqtFxKyw9yiKfD5m1wDW0SDWZsfMzfnVESZnymEuOxZtcnZ+p
4L3LRkyHkp6lJt5Txmh65t45XYkoD5QGGioPa7e+aSZ+HMQYo2aAaoGqGQCSYVFFen3y4G8o5nnC
XggyUS7PICMWTq0pYsoZaguGIgReCDv0HdZCCljtjLT2vYwZTMLKS7XqY7z1LN1EaXMf3MissFNN
6GNanlYWNA6ukk/K9AgfxxxU4uwWBBfc3ON8Pd5fNbAFzyqskpNvjSRONPjRi14XK0+GBdoStzTr
VpWCc9mCYU/bBlmg6pVsNBD9coqQu8Gwqna+bgNCO6F5k8UKssIZXp9zM7QNBDlxxdlvNF/QsUFD
zzrTxK9BxLkZf1Er/mwOVRmaeDEcsTL64+4NLT6BA9PSt72wp6UuX0kK47RrBQc1dNYP/C7u12ZF
v/THqS0zOsp9U2aRNfZMRAM0KMU70YadZXl++NS+A/AD4fkI2pl3bmxF5q/FB3+qp8+dedL1RfJZ
Nk7FMIkvguvXFjc69Tenb43VE+j1jEKyYWruERJaJN3Bi96auCkcgBLTI7qRn4v+9kxZcY5WqEtf
wNu4cJeAppmx/qQkadLtQc3Yrj78Ka8kDKP9d0n3gHnl8D1V+x4foXfJe67eJABrGN0q4GXHr9Em
KV3M/sxwtIqLkN75WqbIG8UHbdUZYh7GSbJUv0UWV1vsCE83utN20elmdGWGDnu0JNZHdCfvAMqh
ws7X5GbF5D92NxoH8IImnAgNaqIuBYfTVUSpFmNaG3CTwqqn7nBv6GSQ9HFLvXfLDy9elmCAdsnt
+CvfluHRFXDfauohRjSnM3Xhf//BlsJ/wZH5QxzT+LY5LR1vDeDXKxus1vcA/7tsZ+v94ackjWig
r+s17X5m/lTCk8vEgDWXR5D0FcNsCTxri3DdMnDBFdcG9rOFGBLYk1rM6GCk/Wo1LUl3EJbGPO0d
JYxiXLclmsX7mJDI8zXuIryNURRDo7qdfqDQGgbW2FLsSlc/goyEeyJ8yzYpwA4zP9FX90jxmTg2
uurQ+ULN3C8rvJFwC63VN+MRNI01u6HjItbOUmKkuF2QD6VtsWpAwmOMDdF31OXyQZE99E9qWUqO
gB9quhdQDVKoqdjSFC2I2ANJ/FTz9KrkQ4fmqc492hudzeofVmweJaKSpsQv0WLKaKDxR5YNOmEp
LZ2g+aJdHH4qddlctsdGz6kmSuVTCeT7sm6k/DrjruyTkzoR6L/ctkQM3Lg02BjVIpQ+kaD1b5l0
FmgToMV3L+5EM+bxkS2pZFdDWEkBwDuJi6dAZGTyDT8IDEOnVv1scCcW1yuP1madVua3BYu32XNA
29+LCQxShB9wb9FJr5/M8Ls319Gf5bxs0rXdeCA7s1vpBoRPTXlN6R2TENoh+2BNWevQSUORvJeQ
svnzpUIMkoJbe1eoVDql8GtWfUwUzz14rlytMx+zDsA+q/MRKRnRMFHHztcB4ZP48RqFZRC7k6ui
+JRQeOdjsRyJLUSubVyUQAdXZbWAeIh3x+R65+xmnO7bDbzK1Bzt+EaB7gj/f5aujR9e5ypIi8Mi
x6/ftjXqYN7DSaO9MA21sOnE4wxy8liQpa9vX9Kshce2xiYjM18Ia0vs06aNAfeq/wfKsvfl94Lw
QjNVQaExPeZ166GWT3rWttE5Z4CyXMEgrOsExVdh8rD9E7Gk8amTE5T6MUPE1a3wQllUv7rcBQ+i
UL8u/olOPXdIy+7QiEGSb77rw2tsXNbFYP2m+GY4SNOC4J8HE7RHHFDVJNETBFfgKOf+WT1qntvq
brMtn91Jy4O5HoiG6FeH5WE3jfwiKVqCoEfsM465yP96UKqcy3LzseZPexsbRThgKCzrYC92S63d
peD5ROgEg0hukjcXz2KYzTA2clbamPZvwgaKFh+obTXZ6ScuD/rtooMVybCQV0m1W7wUxKzPlIjK
214wpx4B2UMbymO3lH6PN5hDWJhY8s7gPhiMVXzAikVA11BSJXpvdqjh423VzoVH++xrGdhdNFu0
6qB+eT90J3TGU64s156zY3vNA4QYiPHOXnXhsOwhJ89LrahK2WOvXkZkZG0ZRpgTUzPuEpp1aAdB
XDauHqZUmCKzkxZLDp8szGYcYiL6yhiTGo4NnFYWcbSNhRi6rIOu8RP2KztqO4PUzNalYt0F7syu
a/YARVftl9ZY3gjWWB7W6SWp4cZTobw+B2x2QybhwhHjPVwBG6Tia5hdw+5rK+3EgRzYMkHCmrAx
gpKhbdV1sZY9c/aPztK4jx7bWumsMw5TPN4Ssu8MbXv4ZjMpvZYeBnCtQ7k2R9gEb7SvAzW2ia8H
ljlQu+30rvhxWo72FXe/96uBn4MJ/4jwKtPdI+UkpaawLr36OnUfwnDAbjGM2kkZoSVrVNU9od+3
CAORkaH23eQ1XdXf95r1Kss/NDIEAzOEx737US/c/N8BxZ/1STyM/wU3PxjY9FpCaX4loURF7ouI
KJH6fAq8VJdnTL4VY+Ps74jJKXG/HJbQ/Paf00o/izEq5eBIpG6AyRltPPK2rN7aa5FO9qaQ1cDQ
SpYVOhYS2Ewzcx19MuKyE2y3JqxNjZh2AObYIhx51L3RjM5H1+rNlHaPaWJWoqoHjg9wZACsmXeK
yutQJqZhawwxYHEwnq0XWor0kvVUq/6h4pRkXKnpZqSZB0oE1zKayv1zO+BohL57XQtI5QjJnmJr
oMLU+5Xw6mSbg9Db0edHR7bId8B/B97/6CdQI4JOvozApCnd1aHIZ4OIF8i3o1EsLfXgyYq5ve93
z2Deu+EWF1qXZ+F0eCYOLpyKdt3RYs6sDSueJVeAgDwRkfZ6MncNZQWCcRjnvNeEc8NdIIZs7u6S
5qHUDZhcV0KlH5Njl1G5TyE7SGVq7M2QaN3et9bTL3qje95sWcDb6pTEqu+ndCrffqrHH3FgsSWb
OXHdXXig8UVzA4E7Y+CT4sM8IT2Jg5sl1YY/kZkDnlsJVejl6JfYa5y4F88V7cb/KVNRz3nZlZYB
Ip03MNXzPxjpuvbtgh2CkkM3NIYBJk24gkW4zOtJad7hU5x7mf4fDT8tPnnHJ8sJ6KZaDrR5zXPV
JOUE3mMva8VmrsjLsES5EULyAKhhRnNypALNsemhnEMOVcYX+swvHVr5tneuiDNDBfcc/nz+d+he
QsL41denkcurbCJh2vx0xTnsgsb9nxVnJgB7vd5KbELdH4XL5hMy8Co6XgFDnXao+NdfaRcBxNGA
CEQe/cPVj54phNGreC8QHE5loT7oKACkZvHnhOzC8cPc4K+TlaLaWNdG0o2lNXBQTrVLCahMx81S
oSMp9dVl/EXt+AOZ8JNML9ahUGtAo/1p8jrr/yJGksjRPiBEVvTFVfVg2/lqySKi1CRV/9mDxlrS
4WmOuYs5r167KRh4oft69zPr/ivxx75s5WOKy0z6zSvB/6Jy69Em9mFbfSx42llXzp790U8n7d7/
I/AmnLjpMmN7sSHV+z4SHQL17ONdEeAVfZCTTOCUbZchzcl0EmOkCcxRGvXuWoIB90iWacpDXuik
lj2sr/aFbXo+UPwBjgTOAquHOG0SJw0tvWAFVgTr9rhRYAafjg1PlT/tJhi+lK3dBd8KYfwH+bhs
nvYHAcoEUubIV9mMNJ1MYlEaL9NHAc7Al/m/A4pefznUxYs9mhH1pscGp10X8wHHQ0Pp2yWnmhjg
qbsyH58KiEaqPStSSU+mmdMXmbSyUMgVJKqG8wvYYmBy9w5XTwZrcoHKtpG4+dvsbib3wYPJlPen
ECKAvrzH7utccC6WwdHxASyP4NFu22c0YVb8rEaDuFAERF60x22iGR6d0yKKhPRHfQtIMjzbpy61
FYIYagnCe4Mm4rUin/6kkC5QYYxxnJaKvUW86+50sAAW0DELjcoqRpBcfgaF/mL03VhY7IGSfIXo
s0Z6EIAuYWA2iu6rXhTsgW1BHJiCzIMUUFL0ioNixBqfFuB4rMsiRtV7Kimyubrss6ESJayzdPnm
7LXcE3Apme674vzYLFvN3xAetTnROwTy/rZm/st2mPPeeTL7GbsWEq3JG+rDJNkQyuiePdbA2cBD
o+wfSOGkxCSiVzbEOyc3bFaVt56IfLliN0i755PyCTubZSJgKgWxrR2mpH4FD1KtkTxCBciVxWwJ
WjmCIewY3pSNV95xP1nn5w3E6i8DodVAN+I9YEaYYaydg4feCz4fgNKbYcVRFm8REWnF4Vk+7Lnj
OSryzrvkv/RSrwRxiJUrJIFgO5QKz1AifHJLlBR8i2Mt95BQFgGfTfIlHJxHEN66SzTacalyW6DD
dbVURJbUFCrziHWktOJb+TKB2AMQp7ogFvAuo3pn64VKkvb9+btzBCbITtWA27FbEEgDB5dRLQa2
QmklfkM9h7BBtv8eK8CvU4awA5SM7uRSzGGPe7t+DsRWYLmxArcS+5NvNRzDnP61cZxYxOiUJpU6
oFyzszy1RjKD41jUaMJceJbRcgTYHPNgvQUlpNgi7sxjrsjkyZByC0pot7HbTXWjIo5YXiQjJJLe
xk0VMKcgVFynL/KbhaLjI+1c4fP3V8eI3WllkI8zzoWmBsEZKbXMOyUHoCsE3Vd7PBDuJh7r3le8
faXHImhXRS87QEKpE/4JuJi151bqeGhSwdn+Xle+9MSlgUCGYjLdnnRvhN6yPrxDgRaV7tUkg+T7
+KQTYzZasOZC3dhBvH/Lru7Csb8UNU2aRQ58hDF6GoP9psAs39HUbCzlwX3WKNjABokvlYhIgyJW
9DwiPStROJ7pF4mDjaykRVBAxI+GezkphgTqbqCc663WywLv25DU5SUZfGqyrYKrHAxj6ZpvLeUk
09Cd6JX9uj9l3Qeh9Z7oLpsJqkamrPfaAGytN2RfYOKA2XUdPPLcV3SVOnGARG+uy67urB5WOq9M
EwVAP7i/uxVaXi29QXlkhntQxxvDzKA3iDUYJGCE7ymDephLgWAS+axJD79lhz2GWKMbrKJ52dwc
5OSI9gchUkLsotBp4qUXq1CUPQmfZqpjxzfyHxSVVzRsSSE4ZL2kRKpP14KJ6m2INmOy/QxtjpYp
cpYIElybWY48K4UwNzKr0isNoQuYD2GCHZzCrbhc258qG1W4ICfWcFOaSZ9awebslUiVBuJv6wk3
fA1yCD2rXcbFZZdBw74EqyB8+Wh2hxjm/VzYG9z9m8n4leuQcVC8QCPshsEBGGyJiboQRRNSdUx/
lRr9y6UhgujXjPrf7AZ+vMjg8dhguvMm1l9B197K9+SgZaUsSfgRn2eHpm/Ln1AdeRXhc30I5VEo
QYTrm3mXgeyJUMsaT7wNFoMZuCSBNCZIIlB9N+jsl3to48zzOdzndj4yRMkPfGOXKeqHjzA2ZYNZ
HrAlUv/yxFq/78R1B7zoctS2h3R/In8bMwwwUvPq2q3MfMn+Lc3pqhCuYjjo5kgt4CyF3JXP6Uav
Q+m+nq7mi/lWAyAzpEGRIqvZ/wN+xodeYi8oZTPPwtczDeRxiJE+MNV4x3OgdcqLyYdJDoFsGXgI
VXxvzAYtHhtFMl7UNRk3uCP3bhGdJ2RkW5RaPNPRXdVhge0nei7/T7s95ZBverWWPKhv+z4eoVu/
YgEtgkpzTr4AapSqyLvAYqYyvkDY+6cecDRagWxZQc2FyQnMojdXN5cPdyuGKJE2qUBndvDlL2jO
pBCvlkcCmacMrTZxbzc3eZ6gM8lFIZ0wk3jzG4AV+U8ykZdwvF1jAcE7sfiKY0CaEHyfWiiPhrpT
VHRTLEVp0d9P40udmI32VX2YnYu7iTfIeSwYilrFG99wpsXnPUnzUj2zpf7eoNuyAG5n3JiUrf49
CfddUOOwiOw8VqQX/XVl49O1H2+Q8hhd3V0HsxMW6VENKtKfMuCWuCFD4pqwWKeV9xRda58iOHzq
7Ec0ivFu5Og6dZvPsP4OQ820881OuksdBIZgH16pY+w17NHkf8J5dvLR9ExvNR60XE64RWx4KtA3
YzBU3OLP38vmtKiopVx5ShXeWwmSBdZeNCiRyPFYaLdrSWZDGPd0mW8pEndWy/XZNNFyjcvvJ+az
N7+5xg6peEDhESqv2i9Gak5gyT2N6CDuLxSZD8m9hsW+aPPcUry3sk44dn850Wpfm2qBweDcPY+8
x5j9pZRAe9SxgSpWkci1PJ1iA/scVte5ZsznLy4RtfJ32dB8YPglMmD/0Xsgw2eY5cTa/A/L9S3Z
kX3nHUUguqaAQEaZzUVEv+Qk98gNKMbbSFMsiiZO1A9UdTAEmu79C9QKwCPsjrLDwJ/rU6XPgN9V
Ei9EFRE1RN52DjP6SLqXhySHeX01ck8ihB9zxsBMwufzvjfyFXTpJ7g6x+Mv3MfWnn5lwGMO318h
oBmegRj4vQ4ZY4UPxxsmBq/fDbJYLVG6tGDQw+suVuzNaA1JS1LJMCGDM8FC98w0/8fJe7ui8GnR
rpXoV3deR5TgSNWNkrVa6o7RqbnuiQ706TB+4wVxy10Yq3/qFePKtwAOid1OtWX41wQaGpaMwnz8
wCdZU/cWUNBzR6JgMb89Il3qq9nJ5ShAAb0V3KsPJ05fm8TKTqgFqaY99XlrEIM6oOUa2iFzOZK5
nVMlqsMimfzP3KDermRC+y3/WMX53zPIC4eQ+RAW0Sm5svTSgB5lceQ/47i2WumhqUQCQhS8IGvS
D7G7cU1avksHMqJCe8f0pmBTyH6BQTp0V6qj8uk0Bro+ipFFutFrndt8mKO2B/Uzm/Y7FYulve6t
rJiqQJ2il3U9bJskfe7/ZOVc1cU7TPzA0jDHau79/s02R92ud3x5cpcjjWQz28nFBjPPZgvXN8yo
2xQ6yRlM8VUgw0JbWzmixF8vX83ItHcSEyXtW9mfV06jOuK7o/5eElbmIn6N5iOBwaxW9KXaaEtg
s6IW0eVin6Y8Lyrwg2ETvx5BUUHpsDYmrkc6sq5naxCSFBssCJ24QilAttPmK4mvNqY/n3niUyJc
PxQnz/0qEB0B8hEacSiS1pA+ysOvVmbxNxLajQkuZNd5jpgEb3bFhx4PbXTG5N2+G6pkuENittn0
Wh2L/shfNhToS+bbwPNH4lPM1tWSoxDM3yzUQLGRzjjUvurUOCgFe0GiIPcVxx00tJn1/1t3OyYT
mg+qEWy05Imiltc7iuFmIBKq4K2UQKBzTL8q7p5LHC8efDk4FmYZhLHzVDY2SIv6j8uyEBo+YzMH
uxR93ei0nHORYLPrGGncYqAWWC+MnLtzzW9lRVM+pv99NI4FvUOuIuR22iaQGyv8B7h83qv21AEf
oQyE8Q6AkYma0HjkiprjGhWbLG/s+BbbLw2I5gSZaqKqlHmhtlghBpEVHdAgOqsfAaEyzhEwz+kV
OXt1WnVcv6UKhRHzR66X/PvlwLnmtgZeIqw4Pxeta1/hH3AlcFeO9dT0uqR25nk59oNk4x3LadsJ
wPosFrMOZFx3rbE7CQrVqrWNblQ8BLPmTRBSzBg7O9yhNX9KwsxtdZ1GcY1vRFIf/DMu8jxQvlJW
pvt+NHn0KRGcR9ZoanVNnzB0gX47N/lRF+8L6BHOgA7UJXQoTiVavxOiSRoYLIT5bJXN/kK4qDN0
dwnxUYBGf//2mGlJLU+8CBcD17d3a3NnyC9N+avzlNhfgYQ2w/RmJ+WZefIeKqWQ2I8kOB0Bx3NW
joock0EBhPtCxY+rJBooIYPaMyLAJyZiMgWM4YsdhAwtnt4Bhn/KaPLbl9gHS1x/cs7eKcGcnPZM
SqdoPZW5AL2Uve2YOOeo6/AoM68aJHK7Aw6E/4Qhr9IAhKStaLQ86E1UP3KV7b89CcnABdSdhVcl
3Lg/D/sL0DJhECBOpXCyRZL5fm9MszdWUUsOQcht2faXy+XXkT+uWIixye/w7ahnNSupZZtJF4gs
qXY2Af1SMUOWmlX7h6tLheUYLyTmcqcKvFQ1bgpW7AFWxC+ECG2PBQ8GNu3GjPAt/GPL2zjnl2M4
FClCe/0blBspYAkd6GOMKV+B6pb159BO9Dam5Oxxmx4113fNr5omQTv0wbjQr5nrWp/ywBR6MSKY
S5oiQIkKMRcl7nFjMklaNa/RgQExtGbc7dKUzJp2Mpzo31xjfG6mXDv2eXykULu4MeX/qLrikoch
sDPekKbT2khrIWZd6jVeOp76XdbwwIn5y/F4jqWNfB29MQZsx+S2Fp4fCpx97K7/oaEuBdI6qQ/E
kX5NwvJilIlEsj6ydInuWqsZNR3GUhY0hKx7Pzu458W8k9aIDWbBxVhtymFt2IYQYuNO+md3rOB8
Xzns7pjWFeQpId5FzoyjMDFjGLk4/4onnmWzOxqlDBvcPuH6ozsz3fsIDrpm5RiVQtfRv3PvUUo9
8ZAu+RfXBjMXHXvBrobgxdIMEajeDyA6IlbBNsbuje6Da5hsBsASoW+mOmGpsVQ366otrVIVlCBl
JZZg5xZeIGUspv7ayV74YpmnDSJbRouQqrmF+4JvHkOZNv+sTJOkc8hTuXJQ5kYPuK4FAqE2mAu5
r4H7hOlZy548lVSspwHXzoBXJUd0wcs3i1eM/Dldgs4x1CFthVUUy3XMmF9ARwcUxfVQinQo7YnY
ysgALPxyTOe8F1kVpCjJOGxVLhWanRxflU2ulUCR9mkr1KIp9qKY+Ki8AI888cZm6/vR6M5PT0xV
rnDYQOtMHTftK0weKd0+XErLRLMQHJcLbvkYKaHA9f2A1FiDIbFPT30BhF5UHWbDbc/mau3EKVYP
VYrntnoYFrRUFwswhS3/f3oavSjQZRE7N1AG/n6hiFH8ss525Au5XfkmMIuS0wCdzi5Pm2IfJBRd
1Rlj/FIZgZbOZGHMw9iq+a0HDo80juh3KbKspkzaINuJYdiWPqTPiM9ccigrcKV7RRlvykoqmWy8
V15qUsEui3AMDCERgXCWnF9wUpTBB+31+2yHS8AACrEs5MvY87TTc+UGOOCCdg6ltMQ0HkqqVDeq
nMJUDP+4NVRmE+xyDvaBWL4T6CgkYgV7L5GkiKOIlPTNTu2IJLhSinW0JWpc+qKTCRukjxLqzG1f
avxfPMeLHLqLuLHQBT68YWMvPB1A7L+DPF6NBN1yiSaibH54o+ll0rmCl4NZR3TChBBvnRwAKj5A
BixD0fyjmanOJP7UAb9PWrp+P/6b6Un3CefxsfO36gFooNcM5W8NrN1ARMOr99PmyZxv4gkMby++
z9qGNYFAtMwlCzz2vBWzMBpujT5gtSTq80PyI1XU0JyJRAlnBuaDX1134fLSoNy2BDODfR5cGZgQ
U2DX7SwR3VxdXdTZY37MXRVAQfZPnkrj+40kvhCkIMuRraNIf4Ej55ZtDKAYMelT8mIvTSF7d1eI
tKKFBvfXifhcemTT2lA0Pt5bXAPrsLNLu4gocIcpAz25oFbc92+k2EWCofObZ9CGGfilvtq7ukhc
ECL8V8lXdLsQm6B+st3Fd0sl+eLD1+uFxTvY74ZuXApUH2ESVT+pZHkHYnlQXF9boeZgh+0UVhGq
ZcLgiIg9aBQcIppNIHPuH7fHvohT5ou+n6GOcHbaIba4JV419Zqwjdgwo5IV1TaVjHhgg1lGkTBJ
nKLhGW/8dK/3KaNVVmqrtUZv3ri4gGptGpzihAUXcJvvIPx4uMOGi+KbMml2jEjQYlRbf7tmOha3
Em3q1lIC6g/ogodwJKbl5HLuI/bWgUBjNJzwkxWIVrJDa5NUkEVnxX+NJgpiObWtslHIr9lJc12s
n4GquFJGijjHZlk7Rwe01cu9Wo1WocL3bXl2JLaSgsXgq6GqNAXIerai1S7pX/khx4GmcAgCRd3m
pZrZbpsJ4Ilkl5pqD/5DlSYSdByYGPhA2YdanUphJPXwaozWnTgmAdgl8HQ+bWSGSn+LHMwMrzyz
4fS5VE8SDzwa5PceWQePFLFeOwa14rLbCXFYcfjVzdhIeyfiaDlAEaXGzdrPaiIyy1MJ70rbY1v6
p5rsYL/G7cVhwr+Ny33rrDbSuwPYU6cNaGL8S7AutPkwVCcE0qfvK4i3LOMO/4Bsa/+VW6A5YRPh
3Hdj40xRPZrrQEHFo0dP9G8sS6MZ6Dc+0m4i5VEvlWvd5Ex0dy983Rlfj0JRTn/662Xz6HVPKsH8
uVjbJPIWy9H2s1HbEXjFs61eB9KFDQLiEiBGjyDClIuIIDVfja4FFZc/1PYsDY+ZyZGJLHWzzDoN
h+tocimVCQ4f64bJm5yj+2brCJKMwOqzfarSUGFDkNG7609tjlD6hhrZSYQy352wBFYk/sW8WvEi
h/7gmrOfxoqUm8JXJw7PBn1M4l4Oy9wQ9mMtvlG7V9ob3lRF1k7v6khaSmPhOTmYA9WII0GCfOkG
HOEtn+KwZhDSXhr/WUp+e3dZtYmQk4VhuR4/oMBtnOUacpUXBEfzt7hDGAzcdco4IbsFv2WQp6k1
PnviKzJuiKtCquYrIQzhNeczWLrT8cmrAf6uZL60WZ204ByotWx4coNyJOfY+J7V598hGeMURfLY
T8hFq2CI5BGIHv9z3fOtP1ysklkE7/gCiu4Nh5lHCG1ismaYpIaBVEdXN7t+E18IfprQmPXH99lj
IeTmISlzHw8T/B5SWm2V0XlMJNDPR+gPUe7EwYnWP2VZIALPNXlC+abA6CnHzTyxaEGDVJhq8Eza
qiQdQuJBz4VNAiGT54aj5GkSe4KZg6h05LMGEIknb3clr1kMb/F+PQx1MfLXPxNt9fUb5wU4B7zz
DHCYYOC//CVQUuz7d2mT3YLy4CN6DqPQRin0Ijti9rEhOjL/Mb81KTHABKvSDyk3j7/pBKqq08yK
sqd4l5V/Wf60i0F9as3Y/4N5ANxXv3Sj50opHI6HKCXCm/Wy9mVFWQxxjXB5XrMORV1XB9ItvObY
mGCVWJy2tE/6dcRiV0X9ybkaziT2tNa7nUGZEEz8Ub/wtXBYAw4veZ5e/G5NHiPiJQ/GtrJIy4Uw
7sEsibFgUb0UPw8HYLzJC2YtNhVthXHMsKrK45KVCbaXJjtZJTJCAWDh9i/RWJ7BDFPd/8ecmwDW
s28DoetL04KBwJRvZoSAIWa86XGCrcgubEarcAoWNFXCG5BI4yC9xieOL9BW8XD9p1pHTRhTOWRP
QCjPYK5oVIUbCgkTYbDpDSzvsjLdHHN3pc04YGcgD3bdQOO/fkqfJ8wJcJUtHWaw9efDI/+rKwS5
O51Vt9malOe5PQYNS/FTHjJO4q4E+wWS5BsXx84nr1m8pk/+YKHr+tiKsvhkPKnn0IWR0ImGxN/x
5eFE0dDn/Ga+mpAuGx6yvTJPrQRXG7lWqEaHMOn8wPpxdYwOQMU0xD6aatn00C8pyRG8x7Mvu83w
DAw2dUEwGk4gxn06kSxG/6XPofci9NxOPPjWo0amV+dBQRIsW1aeZwFsI9xFnOXy3j3gmoW+gEHl
2jOtepEggemaHVTBd/KOY5yGrZdIc71c/w34vNRtjZJIWYSXlbCdyMRC1oAA5diYkEWtDkaO2zIf
3C2NoHSjjo3Lu0Q4pzHqBCsOPq3RUZr2bVu5v0UkTTnePQVhn7mZGIrDHNLdAnHl/+PGb9F0C/Ff
bGfUxvQ+btsB1g/6SKX1uAjJDx3mGKH/MHw6nTLLPP8NbSM+kI6pt6c2BFP0RB2TsnPsUiOUXU0+
tjBEB859wWGHa+7XrC9YlwSzcliBmqUSMLYfNqL/GcOQ0LGqORDYEVtLeDP2Vm0VkAqW1iXBLY4o
uDaJbXdrPc4xt1fmat95eDlSqRsJixCTuIN1MeFCoWxBWLm8vFQZrVQyZZ5ZOQFMedPEBspbakWc
2RjX1tYr9fmNQeswS2M8DGmVd0k6Esb84UPZ0LViOoGkEgEhPMPMFG/u1Ytg8z7eSzQ4/xZBPUab
XCSwmDjBSLt2rvWottL1S8VPMeNIdfQInhJAO0oFmQ9VKCmYiMNeF4AGvK9zBMhcYpYktzYmqrlF
4mdnzVS505vXLemvGzbwHd8tvaSQjt4bf6u4BPL79pt7xyRjFQgcRHxLftxAw65BynlKM/j05sFD
z76e5BQFB414W5uYIaWOAmlP0XPxAtegDAEQE9Qin8+5lYvDz+nCbWUcDUYXo1R1BND3Sgzlq1oX
UVzuE19s44B6kjSLuJW1+oN9Smv1r6iL12Ydlv5ceDNybw6iK2U1Zc8kFLN24z+KmpJ3RpQWBYTM
joYK9M2AZywtwnBmaPs32DFiBos7G8ZgtsAx3ateSG04KPcPzE4VUUjMuYwmrjVzcDQe5t1ztEzn
VvFwmGdcUKwxf9kdqFTp4BWPhM0xUlgOWVZiXughv0NU4OmL0ifJbapeflRCjfGwTLH1kBe0GNQs
734qhKGqqS+gvVv3bcUggJYCfKBI1ippVqIli4wydZkRJSH9gew5r5+eJTSrufmyi+lxMgCvPduC
BIeYiCBEE8V0oVQ3aYOi63Rdp12hsPsEaw+yNODyHka1JwDV/rGX7wCgk9IHEiMZai5TJ8JzHVju
H4bkbVZbtqcYnWJkUoNg8DSrrVH2u6ORoJTl4hIdG894Z1K1oQYa5EGO2cwfNHkpucFp2Au2M0SI
w89oecnNwKQyv0RYpIXxdM4HilSgAvhjoSXPpyYVnxfOKAd5nOcA+OvOZl934x4k8x7rfYObfNnz
n0GNMO65DKhwOw0uzqnE8W73ESFY6IKxDm1+h1sA3LRnWZBK2jgK+KIBlrYPH8qtA7ONRKDHW/4M
rvgHjF1gA7GEyAKRkzegzJa7gliL7dD6ytrLccAB4TPNwSi6rqAPx6Go0iJ4cFnqU8bw2/ztSL93
JVhaSrnvdZGr0OUrjHEsAebd0TUTfWsgeHHl1NGIK4i4+2vJr1tXmdpx9dKh12UdsnygGzpEJQ91
E3nILLZrpNlZBDAbkSpbFj8G1xlxVM5U+C3/N9cYkFp/PA2xCk7ida+bhxY9d8T03ob+kj4SZvwt
7QC8E/nhDT7eZiO40il2n+aIO+5+EfPd2Y+bwsi9Y1IX2NOP5eri7PK8+xq94tSLPtqq1Y1RTAti
QwRe1+AJqvpO5G9hxUcoeljS8v41WfHEInMFTbKPt7M/9o1zddkmxjdC5eDw2KlNTpD/LNYmXvbs
mi7X5kw2zEAwp661e09+3+blhUk8Jbqy48gMcen8ROaOEO/WE4KzbyFGYvAYkg1j9rRJuEHgqCLJ
/KEKNqpaYMQqJbnDcSZQdVe0554s8dZqHySkXwOmJPT5E1y/mXkanLA+n+0BZIDKafM+Vlh+Ji4V
42u5nUImhJaxZLPclNmtzNfHzs3KrQwr536PErWnV0iAViws/4oXJkOswdrleqMmv/3DbKqFTWCh
GIDQmk5B32eIAwAlSkOywAJI591FkVKNMZfvevEvdkwWJtcOPNh0HCl7uvSpfUc/FKmb9XkkZ/FI
2li5fpslNh5Hx/8tcHAEOw1PfrM/cPv8Ps5wXnGoXYZ4LTsChy9fUAh0kPk0+34/Tz9DFEuFbNHM
fHrC5BjtOTrgj0+sf+65Ik54brAGR+K/CuLqxeBfTNaJzI7XlS9zEohMhUs3ltIYwe6FMlDujp86
WEemYsX7ynk3JR2cs0l0kmi3CHvTm814a1MbqrR/RkvhTm94kKqx9NIyOwnM01e6jIdLHIWa5cqz
ysrj9F9vPLFiHcAsHGSJHxhv6Cst0NM1DA/1vWCOXqVLkbR5ERfhQAj9N9+/gGAaCiD6U6VPGxFb
Btz1emQGsBd8YScMznjEoSIgvB2sC78/X/bSTJX/T152Kp90U69Pglc6+xf8vGlVofTJwl1MAa4g
OW1XTKEo7PApnIMNiy7naQGVtGKDANfR86/8lrY5sFQ1dDUu9OoZUK7FW/v0zIsinUGjPOmR3MUy
hEKdNKM6cPd96RnCokFrfYgKtgAkHTqGvF2kFm3hnZDXVt0x8Z6X0tREPcyhbl+rpVbLrIN7PS0N
ulZLHdad2SLotuN5ANJz429x5MDcUWVw5VsrJ+IWr0hi8NZO4SKic2Ewm3b6/6wVQJnMSErbuBHb
he58X81yIcnDADFsZ0h1kWu7c3qQQYXFq1mTUFZGj5ssugVa1XP0jJn4dkvlYsHRCxEsgOwYCDQK
L39EFn70jgTxYjDKA3uOzmzViCtaJAuC/ouxQTr254ytE6VkiQq35Ozgd9rxiyNsusrUO5icKLHd
3VVJD2JETDsymkljt9drBlxAcgOdpGMG31puJKQdwI0HjZYkhsaWAtYIhGQewbJ+CVSXoiKj7od8
MxJ/IgMK4B0BZLk4LmjY7nUoBQCpErzmn/0YvPaKe7xpQwASaXv8nMjXE4JrDpbItoHYKHiz8RNH
kmDdBCrv4zUudWomMHG4Q4Xa7fbmJg27l1I1ol6vQnemvhcUz7+eixi0Hia+5DYy8iK3FYVQMnst
RKne7BNlyySv3lehkDbR+7VL+h1DDTT9HKYld/LGkB0GBfC3kxEJpPF7P+ppx/z6Mjb+gGERY6Zs
96YnEIAAwhO40AaxwV+C8js+IzHgzP7G4e+uVBR86s208g/fmNkjkSoy4bQ1u/b4zWxPWcsrS1aZ
YS7IvjJ7hSjQE++4FqOl1xKg9Benj056dvmaprfuy7lEXMeOs22nrUBA3AOrME5sQlCH7gAm+efP
Tecx3i2g/dzA16vvBlFHDXuA6HjruHCOvJc2E9vjzD8dnYouaGFsYTtXhmT1F7q/CXZWVpCeWcik
jeVT5TcNP4/AIeLIxigN6DhsR/qhfKI/JL9SRSQyDND/QE8OxRL/R4RJdOc3YRes24TsDeBgqkhy
OT7ORzq4Nv1onHLRdd+qL49EQPi8QM5omFN4AEL9HH+uBBzjtrSZBc5TH3RzsDVMc1n8xPPEUwgi
08jnyAZasBjY5LX8lIPANfcXviX/xViubW2sW15xGuzuSK6stGtGmAROp8EehUGCmIyB1xC0g5DP
a0VjfLqqLLnmpakqvkAu2fe8uR/TeHm5k0ALhPQkfV51UdB3+XdbnbXjxjgNF4CFZZdOfxOs40VC
YuaS99uO8tHai12V0lrBc0zExo01ojAy6OgehFq8I+BbzYgw2zISBuiJ23roqzS0iM2arO0daBjW
+Df2f00ELhhEqP5jPlB2Uc/rh/41OM00gScM9h9LWlVIMRx5kFf6+cAVvfHXB5hzQE69JcbEtCZj
OdOlBPJ24ormHsVoKd8BeOgi+R/2fKP+Lqcv3dDPmPCsFS9pzAgXZnhvmDUE/vmaEaPoDAMhUx/N
TECHuExk0iaAxtd3hqtcSUxKqryfStB+k6HGqWKSHsOXDvt0nS4ltp38OBjj6aQnv4ux+fwCboA+
9JaGGxTpF2Q6mEPavIFTcQ1oHVQ3dCM3MfzyuQOoR0ulV+TFAsshFbI6G1EXuiCTPnoG222YhIYP
fPJMv+YJPN0VmEMPmnV66Zb/N0Y6klfgeicnka/ir0uXOaIXvFQv3sJ1tieEmJQEVh3bcDpOfeXz
rGQfHpTgGBwcT7dbSaFCvzSB0Pt0EDXUWWwzmFH3UyZdFjNeVqc4aMUmI6ewgsIUob6uVAtxvx8W
bTdcN40UnaBceE5Ift7usvAG9oemkF14eowCrDmLqKKe0h1OBoCLydjs2HEL8dF2tUOytlH53q+t
HOmwqlOdD06xYszXxXegLFjRxElUw1W0TKx157KxI9PufF584ZBXV0Wys6yL359uSn7S7m4JwEss
Fl9NvCTIokDNCJpZAZU5gVVHN1I8gHzMA8tAu42plhxDeKsm/ZEml3UnTfUatJsT9N3ULqtGp9Kp
bBTvqHMNyfZM9tsx5uek8ZnDGOO9vVxt6ygEO/gSqBA4XriaiFd1kEWFPuSHzXYVqM1u3l18b4BS
7fBzMUyFjOEGqL8BB2FcGZZHLk1qTKdXlG12xz7J4S/ATX5B54CSV3z5Eq2K8G7ZZqcue5xoEH80
AcIf3XqShpafm/EW5Cn7IWwhSYRXZitYZEnj3FkdwZD3Fs6/5Mx2pLLSFcv0dGSYGARNR/mjhgSR
j08B6ZnlG6IntjmAtaDFrzPQA20ZdAsvGclBUNZ0SOvZ1odWGtYAHMK9S5+O40eeiuqxtF6Zj5VN
n0MPmWboZqAAzMnZw1Kl8f5sf/HKHKjLJ5rlTuXKm8P0cb/1D5gQ5cR3gx1dOAuJJquIlquoDSDJ
WDaoNNUv1AtsuNZE3Ug1ticG2zVMPVRp1IWOkTpE2LbS+ATSYZb/aqFtHRYIEOyQ+konB5P2nBRO
yas7ud95haiFHVb3qVtMXKXfCBMstUGT2F6EI2pROEZgCFoz1fu3Tv9NtO3tEIwRL2QZkNndTlNu
y6mLaAQEg9i11+6ND1uInMxw6uesnlSCx7lUpvlnaZXevv5OTE+PVp4yWrnjyOGCTCzWy6rfpfMQ
DaJT3Cna54VkExLjLSRnpr1iymTKxgFGjYZZ/3K1BgnvwQcULJBtetSiDo/GPt5ai5Gf8bejathK
R5huf2EsPd4AifWUsfhGmBP5giJEa156luroijEzwsPbbNs8OK3ySyGxw6bbDT8yJnkcRigQhAZy
MEq1jo/Pqxm9QAscY8Eh1RIi/UDUPqzF1jM9nRqcAdCh36Ba9iPHEzBddfPsO0Eq+6GMVrp8g6ku
IpuwbccOD75qFt0TGfWdScuOhsGyuSMs4u8fGr/YHSH62+iM9X1sZTqFUVHGUMwK3gFWktAIrlPF
7RnOJ13aGkwCTV8lzMCPo0o1rbYXDtfNVEvvmSH/SFsvGFB6pyt4/g09hBw08yR3Jh6sxFlkUSos
nqG55hkfwEwQPCgfT7f8Syu8H/7YY5r+hImUOPXnJRL/ATt2exeA/OavxUBpMjdEMYRmAjaDlxia
+ybrM8899Z0UzQes2fS6l5qu53L8ClbgyRWYUJ8Lx9XJj01XgZa3b5CZtE7KSu6C9+rbDc7Ogcic
3uQ9jLiQo2XZjjFSMCC9ri08LmDiBh4vDZPyYcAWhTsePL9BH1NTN2eOh6uRhDikpGg9j80PDYPe
rKrI4AUwVFvPPIfxiM6zQLZUNhbYJsu7g3+pU258amc/pYM6MiJcruHSKXXGE1P3S2owtfrq+fwT
2gFbQLp70DI9LDqmKj6T9P/PYXR0VTUcw1QSWrjtLNfGgEa6rIWFbw9Mz3rJ3JNsIEXrhZXw8EJ3
BxmYw/vj3T2CqFLyCT7gSz/DeLmPYDXNXIfPbkymc3smm769OJ4EpqjGJxhu11pLRRWtq/Utk8tF
nI5v8GlORz7M7RTbRYZ3hs8UIQEQdcq1qqvC14AtVc0z+DcB+iDHJWAreYDFrMO2x/dMYSVf4ljz
zqS3rPOcIgKtP2kwRZcq9FfPvXmUoU+7iPv5iCs+loJt0qZnaDUQWtfx3ZO94B9vAdIRpSTKReIm
fdCgX0kRrWrqAD18quNh3s8keuSfdhZ7tdKXX6hWobj1Zb2DAAB6O1X1fV8dJ1d/RvGykFH+Yj48
DrspNV5VqBTA1TKpNEq5G8b+7eQHbqKxfT3klktjtGqHDQ+iu9hglM0G7s737zEXtSJ0ZAsQWR4+
9vYLdHHUo3J/iCphssxhkMexil/v8WqtiKv3LE1uPTx1Vneg5L3roZIGQCALWG0WvX8hMhQ0An5P
TsQaLTEzoOPW7wHfZej0H1nATqdPe2nm6tRfvAkj7CscNhIpirnjKbW09jL8JgkTlr74k1Ytn6S6
WjkSRUKnHCamrFNTL6K4/SFhMHYFnF0uaf+sNWSvk0s45DVOxQL469ERushEYz21jO9bpvZpgPT5
v7IOBoTuPtsVkRtbMY6mR7zgegUA9a248x2724I3nIYgnWoLrRmDkx+qfJaZ8IzTCVK/FXzVGtuT
F0dMm6j73ELd0BLaCLbHGjaWDcpUM0UAYqb7/7w7ZkS6pnFAaTHWT+Y4OMeTRF6FKifd2ml3NLhO
RCZCzd8SGSKZIkKPyqrYBqZ/NtpQJNnqGcWzW3WrO8YjGvCYTmGRqxA1swiIwC0wgwxIAfNJ7FV6
zlDBj00FNPbTdJnF7RvWcdO/sn8iGXxxxkqutq1T84ghoGsIYfdo0sVAnOqrxICfQqhWCS0/mzvK
nUV3+Udg4LguvjU+LjymVQdYqQOTYZIKp1IpOlLsWwOL+TUNqtBWrjfNGR5YcheepdhcTazuQP9p
fdoCCMrqWG8U4sgvg2ranwFPmutz0VqdaXrKmtRrMq/PbbWgR7HxprY/u5nbK+i9SO15awXRTbmL
1SBBb8QsxkSqSSV9AOQMt/jZNAkJqR8XH+F6jrH2IGe/f5Kj+NOAcvNQLh9C9UFYDF2BrAbZQV6/
Vw1u9Vto29WCQkjS/IyTwroD5fZoFaIV/9+9MZCo3Ix+xXfh3QpLEW9p4Yk+sIfE7ZboJ7+B+mBd
esNgD8eQm2i2UClGwpCgqx8I/n3JyugDPJ0XNZFQzM0hgoNrDTUJe5tNFOTPbI0LYYfVGwOw8o2n
GCQQfLGVMNAAQ5LFJJmcFYatPtp2ze3XgBEtXVwpvXsOy3wcJ5aBXxLNh7YhHA4l2N/CMq5wlumq
pkYGrHIcTGZCAmosQAZ46SyIjCi52I1vAApRQgyRDi9vHRwUnHu0iyppFiRFhJefrUY4K6OBzzcO
46OR5vHmQgymFmS4UhDFPyIpKh7b8V9T4BRea7oAZ0sZ8U9rpmv83fzbM2vAZTraqcMNCi8eTQvJ
UrbfDfm9FMduh5b+JTe0w6G0AYecndYEXEZrpFvYrY6/90Uk5JfU4qdimNcIsEuj/yLgmx+6JVkv
S4QPOl7kbfmOWGE9gEI4sn91ePYFFA07C679lTGlcM3WUG5sbgHi3SPYLIn9MpttNAiMaAiZyHJ6
Fi9giDIdVly7h332HB/pJlsmqvmolGqiUp8pvdSzKffJF7TSu98VBpsiJRr+v7WTyfstHHjgiWEn
car9oNrVgAtTeRcU0MHob9h0Kd+ApjGqLOaYUBVdXGMpN5S0OvjmTPdCvoEOSST+iev6DFDe1vQe
Wi3R1kMDIlcnfiUOwKyMBCODm5mmnG3oVIRnM9a4htX3yMH79byz2llg8s66WRKiOYxLfDqRMymH
VwZYsFiCqa++2mjZQRYRSS+hFlKh7WjSBtzrR9k9Tg0olRCpn++vnjvgt44gE5T6JieZ0B58Hlxf
OLgNIGsGjJjYMViFl/46qgDO8UwHPyH9CBkW0jNAV/Mzn7qqvnmYxddq+n9BIvHfWX81/3suDpdy
uJ21+lndGwms2vJ4LNigEK73NeDd5OD9Hza3WHoWuBfGuJb1UAke84D2XVIoMrS8zhwnhqSFuPPM
be0s0yapi+0prrCL6nYuO2RC6X0vVHdH4AIfwFLlIMwfzlpf0b+Z++RPYltkyVwl1nE0KEdqA51U
Bi+zobjQdn+lSsqNA6a+vPDAwJHt+3PH39wyWSIzGYEJLqE8MHYzn/rDD0V9fyGwjtedUj1aZ/ZV
2ohGZXPbCS7s8PeX/OQRjY/FB15FJeYsadgxkq29kQg6IaYhougphXrMDnV/vY3szHhnTbqZOk0b
2U83BGyWsPYqNYcNKpmrDruX1ZhUxA2+ukvGIFcOINzYw+kYCfQr1qkjIHH2xe4+rLXNpcMbHwa9
CCb6H53LGQXovxojoedKv+z/qGuimhs6q3vsJZ9HBBo7btCgs2opQb+2n5j1C5uXodipW2uibFNA
X3h6WqGpII15730TjeheP/PheX37A677CHk8jh8WwKImRxkCpVHdQa58hX/3o7tos3wdMgZknqXn
5WQjcOswLnYtOzqpcBs0XhnPmrIjoY56EbZFsIW8NrNphL2qiMBWr3gfGE+Dgy51f6H3rUhQrB8K
bzXKfP8adJpdFvrgEcta/LhvIZCGqG4fEOHaMqin+3RdO5kRUEH4EW6MEn1CHeUB88TekR7hH099
J723i3BG6bXx7njH1EoVFz/B+yZx5aDGtd4kOO6UkDZPoARipnNruun0qNKziA/GybG+JVFPoRwX
gf1c+i31jK/eQv4w2xpEcG6kCv71nn127DJf7nemAO9LP6d2QmQbeLEZnAqExsiTLsZrOdi4JyWP
jSyCK8XMj7Crnw9ne0Ptn2IGJDtGBw6eg4hSMfw8CyQh+9jcmA5iTfNmEax3VTqcUN8+/mufx7z1
d71QfaMCGAhRgTLdN8Q697Yc7tjVKv/IyX3siUR+4o1W4IDdY/FS82IXMirOalbXnm5jG2zFcNNe
N0e2pPe57ZuvGIegPcj6vWp4hmPEaoG2xzowlBlYkfYKJ2AZOUmJe9zpbEOEC/U+UbpJCOj6GR0+
hJiYNvzKcYt7A86KpJJIh9DYwJW3ornLviRVkgS3e6zn3LnK3LJ2F289FDw4Osllxmuxq1R6Uyjf
oxuEgg1DJtQnb4OKzeJRIzLgPQRwhPfe9WyDEqDXwvjqA8uxx/vomahPIvEtdH5A7WpqCg9zBjNL
Ihi4DYdsxTTyqVw9+ustl/zZpr49Y55gxvM4bP8iQg5Jd8kavt6yJB82KgyTgHc1lrXiMJRxU10e
57FKOFIDEs+KN3rvfGe8jG16ACvyfbgTCbwgr2AuliS80xukerzJLTd5j5ji0rS/+YXgANh5xA2K
6ffyQre0S4USswbXUVHe9Ma9IVuo+neFoIJOn8Bmga48seyJKMMHsvL5FifgxupsAoaCY4tsTAjJ
uo2uBtq1aHIene/6hSK+9JSsq/jm2C0c8w+XyJuTN4zse2L2b+paPTKoWHwn2gVQfEon0tPijRlN
6HFmX/PIVWDNQCKkB9hcpd5UVo4iW75RWJnIjjXucA3hUwNzppzp7OYHaZ7SOHmR4+u/Ywj9y/53
rRDywAz1qpCu4LT2uD6SNgnJ+aQw5xYICdfW8AE7JziWfgEWGGfj5m3kp3NStoDd7VGLNT7DEV24
J6rTwcigeBy7YY85vvsnocek/qweGMJfZKOfN9l3upy/20DNt4CdzYA82DPA25ObeFuDXyNOhw8+
qvHT4WgThXQJLIiR7yfXGfz+o2P/MBVZJMXUtl+dryKJvyoTebR9WX1/Lr1/Hxs1DQYgxn8Vcx7d
fuFvC+xZVNCHa8xBOb9sI8uxQdSaEgf1L5zQEnr8FGiex0gwOcDGbGT+cOQItydVlvriZ/ejriHi
opC2/hJqqPW9D00fQgEPytO1Q4S3AaZ7rm/YSZ+M9rT+xq1B7ktFfutI9/G2NPcESCTXq8T12OgG
eUgeTXdnT2UgMl1M2xWBoq4/+cHf+VwyOtoSIxvb8pZBeS6uFwDIq6J2rAcOzyhg/XjNNZo7BVHz
LG0xUOJAoBx1bg0FWcgYvQoioNGwn+NJmCg4ePRnqAOfdzOebt6Hrdt+oQjHdZ/E2uHR4k8hNA88
rvTwal1pSWbKrSddDUPWTXqVjZhEp/a+F4v7dDkY6bHchUtxLUCcB00ydLueKgbw3N9mAtHsAWFu
HnYmfBhNk/ISx/Fz4dcpvytMZa4hS2LsSF+Bx4KlhKBMvaqYjRVjJFjomkKzudaZk4aanxOdCvpK
jFy5LkTOk0oatAckQJcr7g4yMmFPFH1iuH+Qld2jkePsRke99YHjMkmDLd3NoI4OlX3HyHvXoWxN
z67Y+iVTcDWAHXVDr1xoCxMOk4PZS5Nk6X+TaEBxyWolIF+ibfa12q8qXkE/kFSsQiA1CKxCCY13
Njaq/hHyByBq68KG9g+Qa7PFHg0HDaVsQEp8kRo49waK6aMqpSyO5j8RAUWc6/b0sTHbs8uEmZLb
m33uu/4TZtZCTtoZ1cOVhuUjwvVt7SN380PdBSS8VV6C6xJg2BhlMK7W89Jj1GVtlDNXJpdiwF1x
4DSz4Z6XxpNxxfTdbDZoVawtx12YI/95VlWacOfsMa2OpI/3Mip+KSM4l9k5A+yr+uCODZSBmJwZ
N89quOHbyg0sVMuB2T37ckkAL+t3VK+ZBBgL+befGXFVodUZcUF5wDdB4g7R2lxbDNEPYoPJsCW1
+M7KFI3HQI436+sQN7fgsX2tbVfh5h2J2ItbtdPipHOega1KrthwrwrP0GS4cvDv7bRT8qg5S9wz
Xi/tk1ADiaEhoidXHRH6G7y6hv2xliZfYd91Snj6xkCXSYJpCKTZuTivjI9gNqjmbUqf5GCfjwS2
P3mPHpQ3TL+6W0sRjrlvirqh2xvTJtNI79pef0QjdA7NVTQe8siw/dwlt8V4Yv9Nacp8uoTIeUoy
yTtvM2jFhYrjY0omC2YNjjcO/qVDa7mfB3MT/LGa89DssmYJLr22votAsjet+U4tSICcgJz3PmC5
ycGV7PdyNKEIYLwx1F4eeTJgGHrqPg+Yap4vMg7fLFhGBQYs8O0Iqyqb9AVPCvxf8TNh42d5gHq1
dPg/KtRRrO+C19A63EgICAl1DWWf9zX7q0olZzlAcU29+nZYWCRZagD0dMdVKUIkEEtQrGZ0OQwQ
lAuWBzYL9J9TaAWFyhEUxZIH5bzZrojlaq1cIXR40he9MdbypH7McaPy16dllYgKilPNt9rkXuHI
NJbmr4KSYXAUzKsG1t5urwqMHNIYp01D8fPje8MzMUpG9D8mhSnW5HytkxEG9DIR3iRI2iyqw4Ua
3xfgRnF3y49tGODbjyipfBU1g1SJfrbOnYNM6+SHLD3t+TblZesIZbefveVyuRV5Qbeqv6LLsB1+
wawxMV/N9fOuf2HFB0M71d/BDH/jhR2uOYTngLdVzLV+hiCXGZvNKuPC+l5QoK6We7ybT9bAi/3u
M2zXIgceRYAWfMy5/UGKJL1REmxifRHWjvHZqp+V2H3kQYB/QhS0A+4pVvFnHW0gm+z+SNEDkTrY
Ac+72XHx7YZ8KzRP6aBlKSezmNdHQLHDWuAOvSdOObVl4RTM/+TS0tgcTrJcZ8l+tpJ60BMyniGH
kUOMn7I80roaDOgKR0DB9mlV0TzyTANcQFG6s2WX0LdpHjKyLPOxmLiY3TUV9RgEegeuplPZv5lu
7paGKCKzmk/fRUlTVL1ZaBzu3/+RXp9AOV1rsomLQjcY1aKkSdW3NVE7gbksfsFqpYqBliMTDu1G
jfbyyFHkO44n1Of2JMGunL1VjQK/Q8Ly0r9RlQ5kNmanHUImL9gU+thf9YvGBMZI6CW7KV8yOfOH
uV8Ecc/rD4W16zg39eJTO/fP6j0IJeD4VcEgi+N9j8PrSHT35zyl7awo22vjQ7VI/y1R5SpUC4MK
a2W8TqgiNxMIXGTNqJZbacqpI4fyfUaHYO3DybNGaWT3JyRfSKdiwyOAqHAZBPuaniGnzOhlqNdV
DRYR+6htHJIH7QTziQeDJF63XTYUG47s3SxfsUUWyCGosbU9qrnD+UFkjORhTYR89PsgPQFl+mv/
WrG97btzMjhQKROYaHbtevmrYHN7gkelzbsZyoT6k6hJB7Uq2J0c6xhf5gWL4Qb0/BQM2pUvWfnZ
A9Ijf4gsmUYgX4ZyEkOrqz2+S+sXKc+zr5Lr7X7/mTxbYBse/hVvu4vx6wwxJgvIhXLKlqO1xHMA
xSTyyHgPFHyPUdV5nHr6U3jySv4vx5v3NC549uznFkcVPOeZkVbjkoafzB0WXnnZJjZ4f3wx6c5b
vRKV0zA/+pCqnq1DEReYQ+TKzWLnBH23x10IN8NtiCBa0No7M2TIbgOTXGHkczzHuxebArIjABE3
ARcXs0EcW7mStia2Hm61dab3gKJ5joXPzqkIFkMXjMMO0JtlXptDMTJc8jkdn4kZ3YvzdBOzJkfR
z8gteZ9RfxsXDAdXbjFZgtBUoRtWlGNKr745G3c1mqBBB+0AmV9UyjYPzSBZHM7xCnjoZB3KXYTz
Kiqr5x+xeNUqOCWDiKEs05DRqhtfYkwKhISkcDxZk82tpiU72ZSjh88B3tec8ujY+wAuHHir8KXO
AQ2YJP6VUCbdngLpV29S3RlcXA5ysN1nuDBD5gRRR7T7aT41HF83GxLg6yAL0X0Ye73GwU76ZTti
rxKEp6sFmQQE7TNC5LxgfGNcGq7zujF0PikvGaqTx7/zHXyEg+6Xu1m2hHhkXXWzOR4nJMK+Fn4p
5GfShTB5axLLKcrtSZl/wGn4PQdYf/BjzjgC/pQJD2ndk1ien1n8kNqSRDX8ln3IQC5u0FocCNO6
2y5jru1/mEIg50UzVa+xBPdpZXbZX1R722nq2hnok7k0fc45SEgyDmzeB8aotX4D0VGukU/I1IfP
cxpbXjLbeiErd9R50nsgKreNwx6nMHjsO9RXqs6qsaJlFNqvWQRmig8n4M69joUpbNnWcmNCmQdX
au4LrnJ4vSBzsQuhcx7qhVf8WpCv1FPiANE2nmq96tkPHUIfwPwUsG3VSWVWFr76kd0T1WwWO4PA
iS2wNvu7LSLOK6ucYLyJuiDVE4Qa7xA+pkBUoEOCPdV/MwTxDiUNeRcKEyCz0SFQEBTaxX3SOPeO
MJ/asG/1gD34/Cer4TIgYME73hIvuUKBRNpNuc7U3uYNubv8GAtEof0KS/ROuDTkkFpdwai7ufUe
93g2SOoNw2QxabzekqcChLL4CM0+CNZVRjoD0HuuNW2Ub3Qp2HyPW/sPZtLA8fkHq3jemltnimJL
fRwu7O3Y5ehs3XSg2CWy+Rwa8paezkILZIcHEYdjej+NGZ2xlN3985Y86eT9uAI5l77xDP1JSzJ4
VF9w0tKPri7LYJUSwYiUjSOhWV69UgHwYv53rKWFvHqT6DJAxosz+xqXe1FlVs3C5pgrhldTzHO1
q3SRIfv65AnqNuKjWngNFfBaVLrgyQNFwo8rm8yILmL6fIY9vl4FuXHAvpa8oZy86JKFi02p5jNB
aknXxVJCofhOhFQd7EDnljblqNavpRMNXEMhgIyxSWDVKTEUbpRk/juoryQJsIFkKQNBYY4qmUeX
iObrnApS8+aqama59Nkttw+NiMaTbSj7xKICrLo6AI5ggzrOy7+ifC9Wne+cZvT4oC0jbSyw42/M
IbcbI6ba3cfODNK+xDSL+QIpd0jyzRKnq4BZU+TK1zxXdtg2Gs6cj3NqKLloa2I1OMPnBMjDBGyQ
Gjz7isF4hcts4gPbFJSNSp8sKQtW9fM+fbma14ioRTROD6Tm9WOLxSqHzGFc9ZqpfMnt+UDhACPV
xFUyM8gvp+/UwcXjkd31Jdp7Wst4fI9pSwy2mER1x2Zt8HmxaF/ik5IXxhvl6xmPfTwJY/Qw8T6J
KXShk46yHd1DelmhZiv+QxBNL8zaVa4I6WVPGesAVlMZ5P63A9KgwVKzqRecbDoM+aPJgC2f3hbe
0GUzGSe/kqscM+ldLums7tzaOEgfngmg0A2hd70w267Hd/jBzzcys5JYVGNMYXgnjyXmz4NQpD4i
Hvnl5Paf2pP57sxTaraxkawCw27bK51dMf+iSLodf14Sb10kYp2DRmIOEhyUBFo2l2cPbjayEwwg
yeAHQhKYvHVNuY1Q6pm9zSCoy9bL0ZuutwQcP8IBAKzzRHRDObtAiZQ3agLCFgvEfZqYdzze5Jml
oUtCiUelPjZiRnUghIddojvJ/y/8qUnN7FRvsqBee75W+olAoGLAQ+ay4ShHH3m2jiU2+Qu8laoK
KMrdDg8CAu2w8rl6dqXBN+ZmeRQVKHHQUqnIfIipN0HR61GrfP/WbK8wEogKTGDGtYVoV0nhZcy4
RZ1CoFfwhYGjZz5+KYIE28KFHkfPzR7JWzEADYu6bLZ8v4GCNON4goADNgTrWNk7j57zCrgzUrJw
DfyWPDg8v1QnEWHxHzI5D7NU7dGqrkwtZzRIi3/Vv/zyHIpHKZmpveBYZi24eZB5zgqMONDjEcxL
v7lI/9Ez29TQAA4dFkgFzeP9zCm3IqLNlbYY0cEfJ/xPDFbGJeVAYAmiZ56vdDpz0vmde8CEHTb4
WkkcupoxkFjkek5MAzqqUgDyIhsJdFe0F7nfGs2HKFsGVZJPYrPtJdvxUHgdGoZv3S7so+il/cXm
w50PuGRSQQEkptv/taSQBAIiDYpRaJPO/913soGAKuT09zc05+J9e5tXVX7Lu0W6sOE4mTFHi09r
V7WbK7OpCIKgPEjgJVZPOPEkPwmSvSn0U6U6Wy3gkBkDWCKRrP4i2nSdoXo8HBVIay4AiGwOwFCF
M9pQaOvJafEMwkcZGBdqAv8njUc6IK8lrf/y0k4eoIgzJ51BN1lDO2ou7iyTX/IZTMCKQhWwn7V7
sqwLXO7TxLd2kkVmK3TRjkzHlnby4xaWmB/10ozo7dEAgcOF2Yzir5hBecgTF/k7qyJUjG6l/NEO
GInqpbR/daUui0AaQY/nZuYtkUWL74h1qKot1hIA8SJOas14roIQ+ktlcI3eGHPUzhtm/jpexH1X
Izi6ODbdu/vE52sebaGEAezOwnc0MXDFKmFZeNlp0VKI5fr75HBrasRGtx4HmT3BTS0f5oAj1/zl
81YUiuP7poGSE4mYsV+y3DBNqkf/ObMyfuucFCmv7/yVz9z0TS1FT16lh8bZc7AT5utBq+ypK046
s3wCcISFr//+P66tsSb1dOi2BIMFcSP3YQxUzj+XGLJKYoGJPJlIBjOPhlEsIk3MLIoT7MDQYZqP
2Z4K4okjLgF+Ds9mT0F10EUeAzmczh53G23KzWgKLr6j3pu2cHQukIxO+Fr9C4l5mjOkxIRFT38l
JPvwJkZoC3jBuc6TDdC1fBw9VtNEcZ7XHQYU0AlD/3ZgnSivV3TEmthdcbmzOUeiP6fP1t2xyzIS
vrj33E5bdgg/XaV6dIkUQKOyPjjRlIPI5OKiKd78x0eLX+6n/RUYT03OemwsPmMzc4yrLS74Bdtj
vsIDpWk2JnTueGzNtg6k5ZjgeVLPY6UhchxFRZnJYihiSG9sv4G+8+FMBmwV7rcjrbZ4UYXC4Jre
hp+FWhYjwJ7N5cQskAiIkA2l0ZMTAyOwxpY+qii2clk+b3Qp26ANUQvS9m06jAYzHZ8ijBwbfYMX
QqkLq7RdjeP0Yk6ycf1IzIdDqe5sfuKU6fgqHHOSDk8D4UeBkaPFGS/txQH051J+jTbrPbI3Bg7y
LugHzAcjQvXsNBmzn4726GkEJf05OrQ8H31KE/uiI9dvWgJLlihzwjkNZvM8WVte86WD1jjsobV7
lmAKYtxGfoiITlzfzdoqLlWrXxIsfKMdN++fYCO4lAaqhmgecx3iwjkMN9nAqp9X3dgBqMu5J3b9
vfuMdHuXYcUORJPpWwtw8QR1u+vTWvnOw9ow4N1h+yv38xONaBJxsaBJA8R4s3Gl1jN2SBEquDHg
i90e1oR18rQERHONI72XHhXA02yeF0tfkqzc9NSpTHBBzyFblB/1FrMX24uKnZpMraJGUVxWjUIp
V3ilkukEf+FSm/Iz+9p7X4sJNZJiXpRkt/3SsJhXriuD3KoWYxuIgCp9Mxuucz+IAIXkH7n7Mqeq
CG8RNcpxMJZ5r9T1AVkBQryWvwo2tOIZBPo6GVRXrUY2UvC2jm0037o8B2o+ALyWseM2MUvk5SGW
7784bcPw3KB59bxaa5lyKMyQSvPRLEiZjnWw8JJD5WOmepjv6WGEt6k9NEh5HF948YHIz/Hu7Ibz
6wZQiGvHNBb5GZnqqBG82lZOcI3uIavdNwLle0peuzQOSX0Pf3jlrikQE2bYQhLGO2Qn5UAT4Q5Y
ooZJ/vRumYfL7f3siTiDOj9nxCnWixITJokBOw9NNvrIwLxX/x8umfmmQbD78735rDHMhjto9U/W
ll/mldhcFXz5QIIaR5frZReIw3NN1eEWJloPbId/eR14YgvGX3nMD7gDuXoX1aYkDsGCXbWeE5mB
3lxGCuQk0eygx0q3vYITZSaCXNH02kHcDewYxwbVx8fnMNAyoHzQFrbFhDCwKkTF8hVqh9YZ4s3E
IXHBoYxxmNe+UCku+HC9tI3TO4tRFoQSjFEf+BMI6+0aESwdrujLGBoUWVZcXNAthVpY/A3RWtaP
whzMW/UwTCLlRQ2WrndtyWvy4/8T9gqHNkI5HsHl+u24ylrydx49o/t+ig/aM2baq7lrdsH5AtYx
UKYD+Z0hqHBT02XWIhehkA6aA9jWLcerwdKXk2UWF/oQhrK1XTgkRbMYjY59frL0tXqNxoK0eHJI
5A3ANzifY+hdTQdBygE767CJggyykH5I0lVcVHQRB3PfpEInauDHc/D/a/Mm7uuLY968ZEQXi6+j
3wAJuKrXI0hScULWFwYoQXPqyAP/WF5kddmadBt8iZTkTvuqnv3j5Tdb2r3aEHBE2RETrey/frS9
LeiAmpT5Gv0meU4XHzuDrUwMxj5RgtzErkQJ1A4JdMIPlWU2S84ghhfjHwFsxKzFnRhgqCRo+mim
4K6A47XfU3w1Y9SCxOIdzrwP9Bf2iAsSW7+WGhmLTSoMog+wBJEV79rTsrwilZF1+soYU8K/8exc
vNbVyXndCkOX7zZm3i+q0diPGEFtwF48nEmN3VUrbEhPpmTbjHf5LJeieCeYY79P1K4rO9f/IyJJ
hyjlaJojMBjv0q/w3uLvpt64X3eP/9CJNAqiwxXMR1eEwo+IjIUbVmPYZOqm14NBbhWUG3tT18Yh
u1OlULjmLblfDU1mlBD7ZgXLTX7fpbz0uktt8Z6LqC2rVy/q2LNHNBxJt0QCyWiZpaMryfn/V8kS
/IfdDgVBW+ysaDlDbdZc5D6QJAWat6cn+geAt2tvNKSXluqAi7mr1y3A9DzDV0UL+men2CU4Mc9D
NbENB4j+gw4X+LjWlRZplv0GCbnERY+pvI9P03+B1QAXJbkACtVZujISE0hK971gVbo4AJqSZ64b
omwisCDQ4cV32b+ahfvjk/jSaM61wLbsEZ/2Q1SXQqBu03R9iGN5O5Lye6DWLlIqBFldrwdxopVb
YSQ3nywGx58veV12gQZF8bghv+Z36VD+oFhDWhpQKX5q2ULBe6u3sRVGkpUOUW1f7c1IXpED6T2W
/HdHXEmb3doGInCVdb+roSbgPTqxUKjIhyoS9ZSp478Y/OxfqhSY6D8Pfk8gbwRH0/76YtPaFbBs
Dy91ezrx3zTwbYUo7EK8ov4N8p8+qarHs/5oj1QahaVqnt2JcDM/MrjgH/owVPP4XDJltyK51b8+
gh8Qp0LZwI+RV7qBZIbWKLm08Re61o4GanlQg5eJLKsVOQxkh9AaEHeucVHqe0HGcaCYIRJ3WC0Q
pkXV/rrUImcIPiizGOTNj9iYz5EzM4PCLYj/1fWO01BzdwmQOW9B8lgphVXs5WPCSj+FnM3bM5s8
liP7z7FFe41o1b3haA7OJuu0/c9knoWYFDLUUpVR9R9S63ZqWSo9UCBCWcXAC4tv1x5ibXc2oWJ4
vedVAPH4D4J3uzcjmymcQ4odV0w6bfleFRnavJzIpzM96ac9HSOjIlsyXbHJAhSvHV/yowkoOSCC
ExPVmC/CrJNUz+B5W3tJRe51pMNXM5oDrGRBPp3GlZWPRHM926bqFkijeu09sh5Z3+hVvBDCtYGO
HRYRJ9lRKMv7YYhZ9DyCb9LxW+Fp6zqRlE4G2npVML2Q9uCQGvz/ALe1eaY7kmqX4ML/fmnK7e/H
N+IOI8OHthH89riAFKiZ4GJM5MBtN4YY21ac+c83fkPMtikUSIJVxQtmfYi7TtLIN1w/VvlQaA1L
0bC44qF7kesYRJjIkDHI7riMnXfZEXkBFufHsDjB8jsWbsN/cDEH7pG7Qh3cjS8OrULqjS0wXuLv
yeVl8HC2qN5lQ1KXLI4TowHdae01gU9ID9yxotjHKrpuKUJ7BWNwHxZtwy13wlWdzq0qdVM+kdgp
fhv/OEplWU+lasyNDb4q9A0pyNYSn//5EED6xrIAHUyuugs+9vVcLYHOia85ve9rIu59iO35UB/V
qYX8xiqWf7zI0W6/zi96H5t8uFzL0b6B9SYdTeOtZKH9/YK+dJmxsO0AybMruDqpkSjB05F20kV2
7tWNOy1TD0jRPj2jsiBYMsJJ837zwlaDMZwYKLFoWDPgsLbO24HY+dRmahwhzhQqX7w0FuxtZSR1
uepTkyoczlVxexrgQ5k8hmfajef4hck8XInXLR3cq6qAoEsupL5iDCpxNxkY44YN9eVtWZT1m22U
+lIT/ofT5Bd7d32QcYwGZPH8J/c9dxtkWuvpX//e8meYnpqH56SjfbXpPgJ4vSKkC5g683xvVAHr
gBu1wjdWjvx9DrkAnrGXND+Oy1z9ZBkjDoJ6iK1NwOYj8J+xnd2WLqCSzmCqDaNTMT1yW3J0xtcx
u5t7yGmTZyCYRI3NmWExH+zEQoP5X5iHpfzLrKdPP2ZWdUzSG7hPrVvy+mH1rqXbnN+XpR3Htz5p
g+XptXxwh3Nd2yJzjdyqB+cuDXc7cHtVxsOpRH7v5s5WiLb8XtriSu5kXVW9rDA5f+H8Ji2f+XUV
nyAutPjosSTi/LfaKpyppoYqfved1l7TeVI+A4k44fkzUJt5aX6tETBHnwDxvWwBMXNJX5XjxwsK
ozhvoOLhlEbCviUdXlaADIe+nVVPLp9cwWs5npg/jIL9ghIeS08DUXe568CJWXR6P+xKkUXVrUut
U3y/HqPjTuogMwF8QUCPB9ZLZLkOtyDOFTy2GoZAIqwcMg8dJzbGw3/ZX6ohg6VWFHrrz+gYvpns
BR874QKdB8lAuFrCyRQEsognEcJ44CZaNMJUOA9c/CImcsu9UGjHttXqmXbz3OiE9QgkIN/rrikh
Xsf0EcdHJxc+DGXgDxHwSQvglFrL4Jsi2KfppznNlp84qwIUmcwQrG5YtX4lhSbK+gyevUbqRUM4
pLqomW4XULI8OtB+ps7hdejXDh1D+5fahW9lHZk8f/uEPzlwCLePmwItN6NsiWbUJd70Z2zJvmmn
V0njNVCLDVPk6fYg2ZfmkCkzsIcTYz60VUIjxRohGEVxM22A20O+/40DnGPVFkgpFhlmS6NZBGp4
r+9bwtdFH4/gLv5sptd7AytqnCqDYxlkA4boBd+7/IQfRsAMQ7OSudcuQKK0Ttq+81RCIDGVhqiK
P1F4h1Vhft8ejsqeRWJwfSBtjlAUW1oygBoH+0NRk+q1Bjcb+gMvv8Qfuspm24U/rM3wDnZ3Ifv9
GbYFmU0Ph2EAyH7oRdqAy05IlTefxR9+vcajpkejGWwQ/SmFzCkTzW8A+r2A6bAt43+ToZX8PfHc
Fe5z8whUWXYzq32grPtL5j8TwMgBYVZEilkP6AtR3J+9gs9uYok9yfPrTw29JFJyd4uUBME2Vxgl
3uKcc3P9/UP5g87QYoOAyuX8LWO+NOYr2T/c+3dqqEPHImGJnAD+jWRKFKYp0tXXOTD+fP4PaLZU
Ir95NJnVn7U4mbrbrYcRF0Pk8dxz5HaL5o2ccnp0a1080OdX6fko0Zss6iF5FaUw8eWDKka+13jT
D5m3uHlHmjDNFsuIXxaWpdrj6b0iVXj02IqkKXYZXE/5M8wRbEwZ+ylih6pgQ0804GiAIdwUhTpa
DWuFTkp7HLDD9NwtPgzbzCJvhpar74u0rE/OH0lKxgXja0QlG+cgMvc4/RWiPGIgz+3W050c4ZzN
3KIkUkW7yLL9HAO3WVR/ARgYnWd8+/4AwejjvJqYeg8Pefow1WkCyxG1GzjZs5ag8BiKzILxHZHV
xrLyMZdwmKdXgSlgqL9VNs4ODrTA+gfm7WvKwLFtbrQ88YXRzKFqYdqyp0rLXfjIFil0qcsQTRjK
uwpht/bpGR1kbpD4vJVGQdE3IS06a03vHRGD/fHeBDC9pHSAE5hWBNBFzBqA9uYBhwXqHp1ZvsRH
CSkj/3BQISR5HsQg8uv6tSmkATRQBVehp+8T12sNW2hmid30n81PdgHcrlRn6ohok5AMIDBmL+2A
C1y/Cjvcz5oNA8FF2CjGMB/gze4TFbzcRDVYeiGtiWAHtxS2Gt1LpII7ouCwUfi/JhM8LOzQXssd
IeeCPfAjkxIK4Y6RynYgZ84D6rxBLaHsNFcDYh/7Gt+03UEv3BPWWijXJF1EImBFFZt+QTQ+blSI
0Vterwcoe6eq6YvVgN7+v+q7iddIkw+tpFuoEuRFLIhu0bEN/FrWz9YHpD9SeJQ7HjT6X0DYg0md
+t8rsjiIiF0zGTNuFvhQDUKHruN5FE8FViDf19tn1unbeyXEIRmRLJ+PblEjti21UrmD0feZScJY
yHJzkHnjH8ZICy/HvPBEGuHXHe5maL5zjj+uPaUdUmuSi/IqSgfh0125MjN8EGSnAp/pAXCNYEbD
k0Qcb24ijC9HYUxtiT92HiB5HdxCT1YnOZ+5myEXY9ekLzu8Fi4jk7oJ0dUNb/0DcP7yX3WKrmg0
DFfb9iYGNitRPnDVgUdWNjwnovY2iq/D1Z0731LpqJuq3541PlG355NK6ZIFM+IxTlzAAQ6/5CMh
lcjRcXbqxRtSvJrJ8jFibTHFOi4dFi3qyTOP6cGE/QuqFPLnNKlNetPoHNL1GZbYxXaIqgtMVmQW
iEqiqyyozPHGyy3/9niVGPeOga4AMmLhJYZD5OAcVh/qG8TLZUfoTNG0eJAZs9BZLgVe1KGJMeF6
rneOYF50aCUTtrrJKfCdE0TnJx9Alu3JtOdFdedllQY9BfUaZdJ75Kpq7omIN2gc6qPTKhl8IC0/
dsqUQqUSiFx6x0xuO+jilqF3n+Odmq1dImrvI62Lby9YUeQ789PE7bVAs39mJUqFsB30wr61A37k
YimZyk8AbsDsTLXEOy+R5c/ik5XKoZ3+UEHDM+XEWQ0GJLKEmsSHC+VMyhApOSpanNuFkbvs6j7I
MGfKFSOxbFkPdHJFqhh2p+Rq+BfLbT2b/k28t2Bfkd4mBp8fgLjDiOasE2t/Yu9IrZnCtsAaDBaf
i0cjMyt7crxek+8yS0ZOCLKIwe0JizgMSEwhyiGFv+PotNChe8p1yq+KsTpIV9S9eCktB+tH/xHo
9Wx69wv1tELUm34q9W9+XIDgg2l4C0HyjJHe+sxrJe9YNQB4pVEcyFlVtqq6SRCTk8XOEkzKRZ26
Swfca9U+ch8VLNXuzlUL2m6wVYasikRAldx7ZHeJIAIBPa2ZLGVyES6bYITT5YybsakHFxIu+lyL
twbGZABH6IbadXNhsrFMYcDR5DdmKGIreYSqWN37FMU0J8zPz26iglMrtc2t86hEQraN2fToTEXi
QAOGWsw6Qs1X7CLLefsGgOzH3iclAt8LRX7H7o8WeQi9FI2PNZxjtZ85thB3ggwT68EKKphi+qwb
rNSPBqppGQoMeF7oSGOQYCnqOV61ih8vsn3c8AAAW/fi4ivarkXw3wAg5r+hogglVEE5ucj3QhfY
u8ADSQ+pxnrldwM/NmKGXYs0X1FdIVzEN/uJSmancSh3kCMNnDco85xWrwY1BwmKfo+7WA5J6nlM
6oSSMbBD3FA2lcqFGZYAA/bezfib44nzMopz4HnhHTi9UrVuy41KB5o8SYA+zP2VqX7lL+u8pRBb
9ZWCYDIfGsSna6RrzsoGYTgkfFrmIuHq9NkC5pjVBWD16zQzozr5+Zw7xwlVM0zTf/r9H35VXWeL
zNlkSBTnUa+mWGE5U0QRFdk7w75HP6Ugb7c6dyA05T5elO0CQ8DrJE0Z8cskMnJ60NEG4horrond
2H/+Mk2TYSwTD4fQa8793LQy+smlZrP2BOyhOmEY7EVhw0FF5MWzoyOwndAjNeGiEJtYe5bgxmRV
huXwwLBUVsXBVtYP/wx4fLB0Cck9zKcCf9fIBs4cG3/jytaHwsQ3cPdeCvjAOyikjhRll92iP58q
33Og/s9hs94rv0/mPwhWCZJGgNdrK5u+zucTHkxJdJoX5ZYlsyJQ3/zcEB/437DtUk+P0m3J0NuT
8N5HNMA13Ae8RDtOsKPfFrqBj6/ykuGoV+attowwRP8oWXzz9/Nwgq0oPF6ddzoIsM4IEN2HUE68
ZFdFtH3s7rRwHo6mX1n6oaUMyio8StJO8okiq3ZnxHbBXRJGzrl/ttexMCqFjzyTZ6SleKVbfsA3
Tb2BNIjGZt6rOiO1BayA3pKBjh+JO5v1k/O9c0Ch6Mm3RV4JT2aoAl0Nb3WXJHtLc9RfJ8LWWVtP
hxzwjFffbMIVSVIPbrdzv4T2hPEuVap3r9d7nI1LTDsVhE7QjkAXqOfUSWVZ2smTnYEz6kKfhJUV
8NpbzMeepF8uqMytpZTjOJFctpS9+y4thDZluiBOusLYvK6srP57UNlnibRliivEUB4JCQw/rB4b
bg8zCnnzZ7iPedYk7zASPGx+4ZDeAtMP+sc59ig0IizupV1zSjYrc4KRPPkrPxPkR2LUm7d+SwjR
9JM/E66kqUSQXZF+0izHwkbLLuoQyi+Jmp0TV/PYzaWxpBxSWM2DFSRdRen/TXmTI37/N+n6Bsc/
C+k+zqwCDN2lVWqVGkA7Bb5khW34U+Qhi2ndjxYRUhm82f+7UGZaffKKG0SVDPo5iSTBNMifr8ym
i2ZpZ/FNtc5JAFNsrhxsQn/TaYuDQe9ky4dJhnAXvUXTL+Lp+jsYsJ2U5uPTH2DUcfFXIPLpoBpD
btL06lOLY7XPPvHlUwr2I5BwsB8mGfhrr1tlhaiLxvbTH1tY6vwur41vC+GxYuqNVIhVyT6UUAlr
e58Jo97igyOrmdyCmg86HeoejCtsrjVX7jLrhQog4eqTPQ2lI01cBN8OUbdoisdJKiTK8KgMwl6A
JTlt0CESOMORxyMG4WZTdLzt2wTH/EmT6pkCILLArFDPrqA1U4YEG4w1l8oKMi7i+L34PpLf61r4
equWWTqgn2nfLWOdCnL3VaAf9uGg0yLdr3XIEGAti4dsuGt2zLHJY8TYZ0MhjJzvhl0WkFYDHiSH
0Kd6v07iH7AELn8TOuAqnSgWlQBkNOXh+05SVA5dNIvtcPF4w2TTLUxuuA0Ww5tYzpl+76hnZ6jS
m0ZY8zriL2+JLBMUQECSVfkA5R4QzidWgrHQ0wjFRWDw/V3WDaxBTUR7aURLIQTHfFOAhoY54AUP
y90kpLRlKgk+YJdMnpmDPZaTlhGVdltvwy0zbIAgFaCP6JxezwYFryYqZaPTI5QLyFdZpGHWjLpL
bpRELsvUAtUNEo1kQ9whd61QYAF5+CyD27Kn7GO+ZAHOHklviPJsP62SNmU6BtsFKGXoZyWmBZth
62U0p5UoMjH0QjkQPwDcXqm1aPY1dQ6XfXpVhYdY24jvneJWIeRNTNoK1P6DgAEpy4UFzeGQghO3
0zKUskrrtzHHvwfT6F5T99w3OTUxBRfLnipsyTINBjfRpNhdNHoL9yBf1qUVw4417kV2hyYyD5oV
o9cCVWv6I3aH483maihmyCgXKWaoHruL5HIHeIXb/aejyKXGSTYT7kGstSzr44KkFcFxTWt1ys0D
xwW7/GwEDs7xY8BLX3XKe1r0o+o+BNANabcK+pobcgfSa1OmBr8YtMSO5vuQk6UTj+Zt6XtxYnty
xZ6ZiCTuvtZERYKZL5oGS3V5ogrTYU3BqZARfNmWvjcU2G5ivj9wWWYhsvzf0pBAyOzvbaa6ilfP
xSI1vsR1Zm3vs1U5VjicszCW0uoAqLRDHx4jHu/ciBQIPCD7sIgH486fIRBD0J1axz20lZbNTX7S
9v6Pt4bYoN3g+8FfcrlOzTMc7hkJuWpMfmJOMB6c7fwwisaK1yfnVMKgeMZ2xXtAppYVr1zJ5ps1
KVU8rDr76IqA3QjB8PO9XPnBVqpZFbsB5cwYHEep74WjJ+Ezn1XSkz7i6ngKfn1O7gK1PjL7GnS2
cBI9SuFkX1AjqrFphvWEi1zx8qVzRuCtyfZ0VN6U3lZie+u46RwySDx+cBTgBscnW4MG1nPn7rki
trcMVTTTH1KlwlNI3qqlMhhjTEpkrV9SQWnHBxLmaxf5qZiv9cc1ozQ80l76BkK+dekG4pzVjDoi
QP268qYGl15bl/gfwYpHbPPY7gWhFPcbZ+4H2ek9QpgQLIKRSRqPJBXWjDbwsw8JBC/qBVh7Ygp6
39OX6DqG1ntrtwC18oaSBKsytDO8OdzClUOlmDjSHqT7Tv7PKX7aQFkND13gSkBJZNxKcmveDNcM
NHIWTdqu/v/L6ledEZpVHirBdDFoDQwkQPIevKNzrgS2KKDjQxWm+an0kfdZr6Q8/Wjm3lIq4fgF
J9Vpk19SfRP4uguJKHOjWyeH5psmgzYkyaC1l0n61rc2eS026oFdAX7Jh3/A16kCiHa8A1Pwpety
+ZiRqMVfz5L8gzZLC3awgJG91HgEGtRdUSCjYdX1p9T+xSfvlHrdtpLv2Q/KsLxC+3YOcVMed8mT
gtt0ic4xMOi9ZT7wByty7cC1De31DHUaW2o59rZR+BjqYfhfWLyqjN9wMxQsP/dQz5VwRNPZvqLu
qc/HgL4ThnzugLZvKANZ/7LNpvdNAPyWLFb7xio8aUqm+gHXUmnfMMo4pemhm5BNZCpbqfj+3N6Y
5wr7cF9QQAv2IEpzUC3d3elzCqB6ihWk3ZMwPZ1iQP3RqPcR0Qrm5Nb2CeY6oGlk38D/dugu1bGM
xA6b92zB3KdbvdHwuVJa/y52D1KNBHLWQsQvdsp0CIRrJAAtsI2wovIuNUt3HgSYaoiSG4VjmNCZ
LvuiAvkJKGJz/QAPa+aRHHiYIAGI7T3khDpOQuNh45f/uUao2uJHtR5AdbDdTffRXBg2EPKj8Bek
SubN11QylFkCqbmD2jrQK7QcQsH8t0mWVBAPf2OsznftdA7zi/cPstIZvPcK9yTP9HGMWQb2FqD1
u6NorObwNI+l/mUe1vUKVCdtiZBbo6ylSAg0irWHG5HxR/Lrz9ur7kcprVw+3Z6cg2EjicTrT3qo
j77kN0TLssAnDA8lT42d3PCrHABgvYirwFogTvtkFnCQRcRp3ewMMxoOPh+ojUe9ez9fcNMf4M6E
X7uIjrjhXfm/Beea7tSOFQykOaR00D1X966z7hLmo+Zu4Ozd3wxe5SkJ5669QBnnqPV5dLav3LVG
gzPDfSxcR1eSntkZSUsP8A1JB9Khr6NNz7cGQeRy4fECuT/Coe69q2trv8TSql00wnfIY1F5fLOi
IWaVI+Sx4/sm1uzPHU47X69Qk/ypOhRrwqXIZyNDCVQBKfglop6qI/nuOedRLBsuD5nLxPzrnnPa
GiQpE3uCM2PJIy6QEf2gVBn4/IANA9Ip7YMZ8iK5tmC44E5RFcJA2cyRCK4HzR9OeAz+2RTUxbkR
Mdl6J6p2QaUu7zvrCKkkKc/sGbyRGP/x8oQ4Rs+6A32MnSV5m7FuLks+5U0Y7v7n90tces0qTHOX
WScx3vS0bjvzBE5gMEWEacYcYGfgmtMpFT+g7qurYfvE82nHvaJL8/VzllnbnVj7R31xyjuNEsVS
y/QPzBGAa983SAe1ES5p0RGQX/GiUpe6FGSlIaJebmksoD1PuQsS3gqSDmWnzniUBNuquktwgJ0G
6luifUlwOgLnmIgNjTlCa0zxWrAwFr8JczHOaDFJQJ3OU4AP7OihhpcX2yfmV0iJOzUFWJ4+Lvzx
8bQDE55d8s9fieK4Mc+020CAlvTvMeZs99oPGc8P5zqI8KBAbmxfRXm133T90NHnMlstzNpNlh3X
gm0eYqtye7DqqBz2lX7h6xvqKb4w0pjo0lcQ0NlZazaunSAQc6RRvw/Aq6H09G03B2QwgTQklyqv
bcSrO9ssEUWsoxsL3fR1rwg1TXP7C1ryoQ/oWQSmQxmKPrppg5/i2nUmOrqzoj7GI7Ybfcizkq/8
tniMmfIZDcYDHeQSBFG4EV5GySKNp34uVZpZiE38fuz/0Sdk6VdTwC57fR2SZx8LMV1M7Dc1DILw
aDDrKcgw8BnfBs2G/oGrBulH6++G9XEQiA6py71NDz+/MuScKxmwJdteKMIEpcFRn6VDBiWbb4Bp
A/+yAFggc5s0+lsGcyyGECeGvxvfuAucC+bu6PTXy77Yel1pbqlPhs0+onNZZeYhujgsaRxygstm
ReuI6k6np3NC4cEhJVRydl7MeD5LHwPTAzZuUa9UcfnRQ5KDf1lGM2tX9wqhiObR/dAdbTIjK3/6
ILLp2N5soDZBMLObLZEslh95xuIeyd1ZXrQWCO5fYReQZSgv2NyWMs5Qjp+VDXGNDptJtsIMBGbA
ikB4PQgcl0/21tcJEbSBmHB7D8MQT6cpQ1/yo+IE0Ztu40KaD1bQZI9d6P4FYKWUCe7SciVLKzzF
t2HG3r4Mt2sdeZBkvUtnpW5y9gJuxJG8oJUv/LgSVkeLbeC4Qswqs2d+nDs7Fc+aChV0//NGxUjM
w+U3c+Qy06mGs+t1kUEbZ5jtTRy9LogdC72ekT0NgJ5QbaxXdmIryoMTi5N4gAiKdg3k//TdIENP
UizGZc56neBba5RrtACbG5k/nVd6Gtp2GjFo+NDNRNWcYvhuK6lxmyDysMTjAzYalwAG5KkmLg6w
abjEAs0KfIp1Sjbp00YunY6ntg/gIyaXSv7ywJiJm4MsTVJJSNKExa/GfgG7qg+q+iD9fbaj0Rvk
+ef60A+0F0T0ikiHAKCk3eXkrWHePE6VP02P33AgWpmQ+zAr0lBJkyfE/+EfMIsCp1Wol/3I0kb5
9pER/lKr6mvs0Aqbb+lj6UqRjCtU3Se6Kdte/e+9Ev6jeWfs150IwQY2KxXoR+z6GmpQMqp2l2VZ
P7gUz36/iXYhpIv4FcrBgDwG5twjjx029Z9d98FdjNMi1lKOnILnG9qifCKqoV8Cjj5C8x3b17Ua
YRse+TgA5f0STQ3aHgCis0vVUSe+9GqHMbISR0fAEtb8caGB7EUhjk95jVzsECJMMasAeK6Z/02C
LVLXvg4kfH4mGysjA55DyoyeRPLMaKbhQImIBZYAD8s3oDURpw4lidP52h4q1o57dDGnMHW9OrBG
lX/E4tu4N6m5cOB/UJnptzKmbATPSJ80dQXOzcoWNVBZ4FGrSLL9o0eEKBBrPga8uv7AndGOB10e
ZlTVU3sT1P/63dFHN1sDJonSkaCJy18/7gpohC8KLeQeUJBGEY/9l2xK/Q4wuRVi4rZFXkZlNXRQ
+WelJAPXDZ8s9yLo4boZ29bEP1iRyR+8r3Qwerk5yNkVB3l2rwTxCNWX/iYHZldQRq78wqduyGvh
09RVpy7wknfdcV2P5Udsq49EzgCExFuSVsDl7QhVWymmruUGTx9t3Xxyh5xzCpob3nvfXIzjdGt5
CP5GpscY5abtaHF1ORBA1D56eMkUnoiPsWV65wPKckC6TzgsXhuRGjeTzrwV8ozy8xHcjjf8oHM3
WF8KPw9zBM+4tIAkl3XILIpxTHnx6JlSTrozb+YtjJMvcpasnRnCnfRVHI0ahRTWQB688x8X9c3T
urEjX2MTyPkUtI4f6Qr2IWmkDQWxls4GumjmAuDBxY+8vtkTVOjdQs5dqPIhIzhYGJaoYBcAIhXz
TROip6XzLmOX7iO5OXX03QJm8nZMXiuDV14MRFd/4o6GEb+Y3Ti4hJHeG6SxbGby+xXiPe29tPCk
W6dYwtwLX5CirWsA42UFJY63jgsfF0mg2WRy86u45cRK8ufXEy/F0ZO4ql68IUQJays7n74ItVBh
acltw+spofN3uW78+E9YjjARS17sI1KrOlpQ6Xs01IN/doYPJqwQ6E2AbB/7EfTDfPyOUVSBMXJ/
XLMO1f04NbISRW02FpCdbrPAPV7JPxSIxq72HiQkhKLQndYM8g59Tzq9ODPoNESRmmoUinu9pRvF
266MDdxUFyp5RB63Jznw4FPk//tyUH5ic37dnsDcXEEqynJYtovy1z4pKpCPtgoA90z3mpzUXNpN
p3HyBDHXniy0lCfUkedttrvI+U6SzQIZLDR5/Ifs2rUeK4F1nVd46JcGwjl8GQVStYQEu9HmLQZo
01T9U0jHCr2CvFNWIfDgdOAYXf8gceUUb2Hooh6W56iyRd3FaCtZAQex6rd7BXkAlemwEBqexAYr
XMxrvkxcsRENtOWgc8KzQn/iwVffzRdzXXMqgXUl8a/eifN+/3amQ++H951wguc90gc1eT7LhJKi
qpM7o8hlYt8BqllJFZK7v0PcqigaBYBe6euB51H8csKd3NajIWexS1QfjMdwHr3pWW3mxIRkECvI
w7DUabEEk98bOoVRd9CidjZUJlk/42pbin4xEZF3KTuF6AGYdFXHxAN+oPVV4DdIXcPq2aRquzdW
ryDw06jQXohoJLXaVXQOcY7lgMo5U+F3AeiJ1PBXdfxTQVJXzaB8BL12tzcqljiQHXwdKezdeueT
+rR2AVp5xtNV665yspW/vfok/x/MniVDGSPxBgm151uynJhaXShxHkVsh8pdNdzhRS26k/lzco4R
e6alw6vKwR43GXGYC/rZ4jTbBILmzhH9aws4H6fHM/Ah3SM1c1ocxHBRhIgI75pFAKa0WWykY1Yo
CthTAYXBhihvRIon8c/q2fb2nV7yANm2pyB7w1esI+/PIk62jOYz+60H4o08GbEuqzltyNO6Ijil
JPLynSvEC0U6koq35iCkELon4FZcSpNJrIT3WwNFMQEweaHlVVw3Ur3RBF5kR9X0l8761IbF/Qst
qkWyIP5IS9K7GPpDNvSCHJSSf4UIjwfKsSMc2hr1iIcsa7DgTwsARDrS2UuHev+F3VzDj8BWllY4
PgqNmeyYymp46lUS0cHIiNa/6r6Gm1GDSzq+uBPkuz9mcR68sal9UFe7OK8qP1sE/HwLvSnJOL5j
xrnmxkVYb/0VC8fP0QN0EFic5S39CakvutOEqHctBMUvmmnBF+lmsgL92Ph1tzkzTTcuKSPv86Px
ZpOVEFZ6ZJ04LV14jDJLMYRxmVVT5Se9lklulgnL3RodoVUuk0UzPBmXc+YxsyXwqu1EBYg8Gk2Q
osHULlEqhiCUViZDANDyahAFC06KjdJw2cKXprP7lb9k4BNrbSK9f5BDIXcuCpVVTzyG8Wp+QcWB
GWZ/2xnx6c8pH5QzIpB9qBlr3lsTuOjVcoQ9Zj71CHJcYwK9PROhq3+1VtVMhofT/odsdu94yH5c
QMuvMIb6Hi59ZGGT0xKEiuHhT9aH91MFSA/OY+6Blsa3R8YTFJT6LLGLpafa90bIkLRjwKGV3HVf
sNZ4jtXq+AK237eDtYBMnXbhjHgpEOhZM/fxicW93BEtm2a31W9UojmF54K4aPOgPcxqNKnDPBHs
S+kU0kA98AjR6Ugn0lTTa3jURo2NxdBIog98udjWSuswB0Njxeapiado3qXvmCEH3WTf2VZlOOFY
IIffrblc/XMcHhwIFIg4xFmFLQDfLOIZD9BMZu7Pzq/2Q0aozh7UuKoHtuA5UiXOK5E1SxqwT/A1
vunW9cgOluA0fYObq8XrZ3A5swwTIO+tvDJIjYfknzId75FhbcONMD9QQ3Sn7j5HKGPidRWTcaZQ
R64hy4jmSr44hfXMzOqUKU98S7BkBc3bwCNT/b37mHQlQLGDywAU0k+z904ItdiYhqlhP84ELB1A
dlJq/rnAD1QPQVnNXzCEdHErylKeeaCRhyhA+zoOiJ3yt4YUtFVoyLQZuO7yAHx/wkFBKMcJp2RP
32bvbLxHExI0ud7y0PKSUdIIDQaS+ysLOk4AJLVcmEeBbm/aXzbB1Ug/ZbMvQl0R8monaTlMFjWx
HTQKngQzFdkapeaOLJ7mOJaJetB9Eg+pPrwVlx950Md86mjbKxBGZBWcCcTKHIdAu71QXN/RmleD
j6g1goQug6yVQkovtVR+l5/LbEHp7OmGd+x0XPd0eaaMCnfADTrjz7V6kWYIxGH1X6r6+Pw4lEs6
5yZAgDo75SsQ9H3T5tv0nSYyzGdaIlJ3/pjHLzdRJFBiyBQ0N+jgxDAM/elK+KRg1wOtPsKKFk4s
S2O751vAT6UPiezD7XBgdcpH906jvew581hj9c0lCg2dLHrCXvG77RruGZvxze0ofkFOYdCOBa3u
ZscTLST+W+kjByAaYa7Yuf5DcpXYTGXKOEF0COh7SFNZD7hZyXJvZZwLSPYUiTmmX11MOXJhS8k6
rs9zzNjn41NQq9irD/u1BLxEEovYlXi1paSgsDsRIsBfRSWQ/qymgqe9g7zN4ZQGa2HgLUqkSbhX
1ma8s97NYoh+TcJdbvMy9ZmwcFyXaSCIroGBbaW1bhQpvT8liXrcRcmiryunOGc64OK8efJBEF85
Qi7nVY+W0Ty5UuKKJ2bYuX3B2dviOFNtGRnHqjrb8yWOxFjhkf8egRik+3c9DVUsX6schx+9PxbA
BqAiImN2RH0fsLJF8C3gwpqcDP/d9JEd1As7FN/PL/c7e7/JFvr1E7KzPunx7SVN0qd5jffdMTXF
4OuVr3jcNQZIqgbtVvPBAQQrBRbECKNVgsT3NCkR9yMNHVh+OivAlSbTBoF8TLkcHm2omcXA1ABQ
zH9kXJmanmVrHpzqcfOzNPqVjxSCe+D6DdqILAnwTkiOvOeyuJG0oBeCzphUzkDuv4Kf8RvmBltx
rYjynayoMw46rVSQnbl5hNjpiwjqqS1zcCAAEsA0aBW2n1VHMYTk4k7R7ueZF7rWKiINQ22+NRFg
ig4T42OITzvLkuFMSJiApvXqybz5aelxI+UVyXeMkHC0vdJQRRNSoaRUJrTrYMdpgeWKFnl8Rgtr
INbIVjP/dJpCksd+ALD9Z/bZAu3MnSFkrOztMlYIq3T5hutLcpApyPROq9qZrFhYn8oM25CFquxe
yNcvBJ5sUzDr2k1ELtgbvUS261rwVWAxjF05IzqhFNVSkZyYGsFu077Jd8j5ZVYq3ezqHZiBCP2S
SC2xCQmJkZJvoB1M6CgF9PBVV+Ff1tdX77azpdMTlLtGu1xqfJIkAYwKzthS/cYFzufEuz/9rLuy
EACTC3HSK4dcXGE1CUW5G0fENXImm93wEx83XLNPtZ6o+UZtxLBWTBklMmwbaPMSCLF5I/9gnRF/
4lKvsqJpvtmfTArj8xFGdifuTrSe4dUO2HXxcH20H1aREzVHKryIqZn5cMCDnztaG7PBW8ph6rgo
jm9/CuH7VsC4GOYlH3fwe3iGKeKDeAVfBBjb0+g7CLcjWLv7oOwijPP4RXPWsxNzJ8piK3l9bqhp
KCpPU4WagNejwfMVxojKIKACTRj2mnnGga2fteSGh8I38Ygz7kxjMvx2yfHHxLN50FKcZlmJPWqV
CAYzXWXK9RN/K5htVQ82jWPO11s1RR3iMMSn1uZmjVO3TpQsordwHvRfudxgiD6TclaGNbvGa1p4
eGeXs+DSmSvhxxzFb7BNM/rg+dFCDgDqaLtdM4u1G7lJ6EcyFSi9tfIkU+V5qEdbbsVUi4nt7d3d
wsQeIThHP93gB7eXizj4Qgt7/xPGCcIY+XkjB7bpv/cRaNgLKZ27PBg9uY0TeVhZwRPIyfK0mPCA
hNadK5utUHtIdFj9sj0g/j98pEa2DlPx2vSKypmGbxP4+B0rhtfaKH66CurXrdVIQlcKTWs5sn1E
7HdhuUDk1wA+V2rNPQZLvYUE3jP76s/kUzwwrm7rJ3jKiroWMjmBjuklfoBypagB2To4laZiUZxJ
M9F+BIsbaNGBhmuOHqvRe3BFjo7WQ35hlNqp0fg9hZVrV5VZc2tdzmktPljCJ7kOUZgVg6D4Enep
3QV2JNkZ4DD0bgYk8zFffmcdKHmi2TR4ePp+xzTRj2Yir/bQ5KVDcGPGeCGmMPCjsJsAf1tZZ5TK
x55cy0n5zTLKf8crzKk9i6ptscnZfV9bbFP7OQbK03ibgduWs8XDQ6lnyfhA9Z7RU3DU+xemFwnX
7FN845c2czJb/DQzJo4uC+mo2tA4CL/PkyODhY8EjuvRzHOckpTv9O+3qY+rafgB8I65PgFCovhj
t2xmMTQ17udz6zsQ1rJaOR/Xx4d1DKTdZjx2xTvvUmWYIkvrgb/yxRiJLAcTAEG5L6thl/zJhCeG
Y4sVVJQZ+hDu+kuiC1OYvoF9NHtQzA1dlV6807cYhXDKJvePuIKP0oQsqB11jxBOb64cFiurqpr7
LqGxWREGaPkQ5dwBYkKn3ebgkIwjxCCIC1KGTz6ueBaec5xQfaLKUsTyVzljJeJkr8qC733PbmHz
vp4nnkLohDb63SCq0QB2GivIeshU2DUaWAR3ZbdkeJJ05JNzfdTA6l9a17zG5lXDSVxqHf3dlkYc
mMTx40H4Q2ewXT0x7//gJlxMpZf4PFiDIkJFQKUEqgmZ/tE6Ufdw9Mb9674xDXdvvEnzYuDQTBeR
03xWrb76S0x4o9efWjLuf2gQyZOE5aUVpqt+2WdqszfmtuVjHfwUmNk0GROOlUkXJWs5Kh/woibq
US+sfNnKqtp1ez7Z8WzrASmrTCPuE7eYbcbFjoOALp7UcG6yMspkpNDghqHAweosW2eYs3o4q4At
ZXhvL10BCBsTzjgji04p282kl4JwRBbBF1USe2dAJCkoj1u80ZX19o2lZ4w8upA2RQp5GWOALzEc
xH+CNZwDdgHU0cqAIBeZgQM0Hf8xQrBLkjg6uhbiogKYcLgajg0dZWshHkYdvmlRxnrr78+qqVM7
0Jyi48L05IDV1C/2GLJqVx2sQ18LUaYylrkEe2Zei/EzGCfA90KkZA5g2SPyFDf/Wxsyz6endt9E
LTYpn714nlw6HuqVt+rxDjfATPgZhIKUDyLDo6wGmxaqgyl5Yk5WMCqhclaZbCBuz2G6Uk6iBeTD
90m41TSpxIHiZTsl6z0bQHVl/R9Rpsa5OoBMRRUsgeYuzudLGZaBriNImeA/fy3XNhEPm/UDEZvE
0dQ8Oh8etBhcPeQuutdQ6G3KejzAGYGtXyu9HW/qqhMU7+wcYRmZCvEaUqN0pnIRUEvh8U3qvCvu
G1HkmXf6q7/mR3nQo0cO4Q/msSTp9vrnC2JH3nO0POXsbb+2/aZFzEsneF0n8+YZf2BqA0aonoNi
S4Kzj91ab/C1L8E9E9l896jYHq03jBHl1vJ3zF1n2wKiwV5S8+6X3V8QXJKJ05zCk9etAcDobOQh
DPI2iiQEIWvdF4PJRR3IeV6BaNmRDGrFsVfGe7SizPloUWmdT4uKVN8Zu1DOu2nhuu03sqBSQe3z
uiX4cynkXgLC647UZtGjPF3GOaX9HJqxVaCFyUV+nJd+QsLAkP4M47w9R+zW0NJ3z09HZbZcSQx3
+nnFfWQremvSSSJFuVcSl6cKJmSJ8LSP7f4CvLFvv9lLc72TWfdPZfj7No2SRigGIFdUcrjTlm3d
OtKzbLgAyUgWGU0/SwjR2YDbZZ4IJ89Uo7sk5XtZlUycNHOraDoH424eDxnT7cmIeYrfwn6InVzV
j19W/OPmxMwloDM0qu5CJ8K2qvyjLLU6JIGGqAJz/9sOrqoj83DN+RxvVFAQ2Cpg2GG9LXJMcEq+
NAPwDHcV4tIf5saBB+lUJInh4H751rECmgAPmEeVrKWg0qzSK5diWWx4kiAXW0eglbpUghVdiOME
fRRuP0vi6mAaBAeubsRYIPrwAS644bIjwg8/7PmXBygJex0cUM19X+xVJbzmrWrJbBQp1u2x3RH7
kKeKp7N7BmqUW8YYWNL//QFdzQm3pUFV/0qAAXoy9ujEVCeRH/g2APzPlMvIFg0iI9f8yy9eCevr
2T2gT0W/q3SajmSBqFEdIB9sZAXiAW2jbg+R1ICFgfYTc5a43ayFgHZ3Dv2WSedz8DGpC9bhhkeQ
gXH5Xh/ypKLsuZrpozwsmfXha64ZrAqnX/lAa4rJ5eCIj4a0pCPiCdQcRhQcDDagKrXkh+A86uRB
jm7bBG7/CL2iV620D+Qm55TfGCbgPeTN53K/QQBq8YmHqulBEaejQheU9yu5W6Hyt67/9oM7Kc9C
goMwEPqFJ/AzaRyMM42JYv2+kOFo42XfYSNcZYV7/4tPW7PZ2os8am08KRZo9dftxorLfmT3q7E8
91/+BUsZPVnOOc+t2zbyXKo5SdqvDeJT4ozB1sRa2eqkWhe1/4OXRNzxB8fwEfzyFloHR7NV7nZo
dUHvXeouRaIq0J6LiYI/68Jy4RyA/qGpqiSbEJ6VXtKIbO+5nW8ntoztRQplS9RuvyvysjxkJO+C
yxcvuPfuo9T7oaKRKjtY0xNql+Er97nxmCt9mhyC/Hymvqst/Tiqyz2EINWz/0nWRvAGVt10pnsv
JbKGG7XzCF+CcMwme2zI7V6xVDXxZtTIm1G/WpMtmY8akoEESK54TNI6guBj6ZdQFbwEPSzukQEL
O2+P8TixYtlNFTexXSnkTQmAkw/1AX3pwRik9LtatJ3MlyRpUr5VB+/uxn5PdQ0cJjaJCSHahsDv
ghmzvX/PCdU8eHvUri8/DM5w4Vd1k+WDwD3T50z/EfmbjYKOm877vwCS2m5D5M1iTteFX3Urd/6a
I0Cd/OebJW0LU90p9ip0QqDlrrhthnrKmnwVwVpzQ6eGWKVMt4+gTOIoxLpF8WRyUmf5bya9wB/5
hNky7x6zvAqchrTu7N9PWheJvG4OELdZY+hIOgVB9fODGhgIy4/hPdjiR6QXruoLfAHSfojFEs8E
5DyNGjmpEthjpLgvbpFSHrlK0ORsIrKZQrl/CLCTZ5E9d6kmnWjkYlVwzbrxvmrpddfsBlEnEZKb
rB2SJJN2UszZiXPWPVn0ZuPE4lqPvsazd7pnSj43CXjlWX4l27jwFFrurQ35xOdF70/UDW9UlsL5
nM6WNdEYY+5jPfhdgxNHK419Oy8NCJRrwTWQwO1xQy90wyIYB0ciFy/ApURgQ8nToHNXSbgGY+jE
FDk7TwQXwU2gd0ylYhoefcV5kNdjEzroRj94jUQyFoGEC1E/bNZK86BhWVahb81W0oQRSv8d5dTs
oDlfCos25WxpSCaTFsyXTuwbeAou81syUNmnc053BHy0Cg3QbxjvV7gAUYHX92cI31GtzZ87Up6b
H7Ek0rVhPItW4TLJEvz1oGQSFVDxX1mca3yFAoimhLjikL2sbJtEJ/KevWyRdlOsc7VR2y7Nm03p
fO/XDc+H5UaHlzoNNxuxsnHTH2ccocgQH8D0wuUhCDyiGZOEFv3tCJEpXF94kMGPpks3tXxBmy48
D5XVQKd0fXLgagHZjcwRSKsI5glJzUwnshcbSbyRB5HIP1E8K6PQUZ6xfq33fyWh+wDq7vIY+uWC
tAc9a2SK41FuJpmBrH8Mb2U0X9O0hoPU2Ir0xATlJAwTrnd6Dg8jkpaYH+adFIb7Hd3KmstI4zpT
+iSkSNa9fWBPZJvKa/PhSoLgUfjPCQTXvOO15RuewASegv41oTxVfI0SWW9Q+OOG4UapiZXHCl6B
j/FlfTQRBQkgOci9WsYH54XzMcNcFAHbAkwI2uASdCg2YibVqZCF6/KT3H7N1RtaGg5TkLs6Vw84
PCsdj0JyKACcZsYEjES78Oi++dayA0/b99LvIi/INB7qd1kckwMRkb371wsUqfmK1Wb+sfeMASAp
jy5xr/abvRMFO6poc6OP8Ai5CmBNFgzZ+ssM1vtTR69DQhp2QN6jUXiEWrN6sk9hNQyRt88br0VR
2Yt594/Emvu5j9ZUd3CvC+klsh7uhp5MHnyHRD1Ht+XHDPoJIECf2NrXORcrjTvNq5kx9Ianaubu
g2VvkJJljIgKmkGafy0yhS8Exjua+SAbD+FB3gp5DOOBU2iFCnZXEFpB9I1TASxMRChoYUGfiBTZ
ddA7cVm6hPiSBz1siDjZhLbgKw6BEFb6oNTcTmaSgMnj8LWY7PRRpF259TisO10VumdH618vVNOr
XMjs6oUkxqUHYTiJWO5doPm0TuIlFui/iO4Od5QCwhLNNFHZX5XecbxHSYkPK6jgIEjO251ONRjf
GvU/YVvsrdB1wIZf6iP88Ex+sXzYUS0SqMOlkyILbkhg+QltLxhIseItYtivsUYOh6LNHqF1UEI6
cf2RoiUkAu2Ff7WPYG4yBwPv/2Lavkss0cZD09fYCqLGD+8dUdR2F6/GlABMyadFKBdNaxXo2zuj
9+sDKjh9rqg0swUi+FRi80MncXohlbWA8hBXiHlVJI3VZhWb28aA1OHCrAZtW3lfpUkKJTSWwt8s
FB0quES2WRSKN6Mvd1m9uqkPGW/e07Zau/0/VnjgdjxX90fS2a6EFUMz11cjw8F4RjAiKB4W+kJq
tpuVz13lT+SZ4PPOGC2/e6Xvxi5PM9K3Zjxal7eVCDYVXd7+fwc4R9HeP4jlpGWSd9sTkztb+TvV
1fzTdhCAhuIOmfsWM6AfzrKhMMDTRkqy/R5w1Amhin55UthdXsTIhChnehzjEvPWFnrP2H5oHq+p
hwf5l4S9TIlNSP4N1ghHnSvE4q5yzI/qqIeVndm+qewU3N3y2wb/0EYOXYizWeD6kRlE29Jvf9vN
uwZ3jAdFhBYGkoaTy1SFShbXMY/tLVp6kFbClTIjTzpvp/Q8ZwlrV+DJY2nj35I0fBJouucJtWmU
O+PXztAWpTCZQsTnAEgpFpWMLr1cz/yqr2DphM83/XXo5G0LUd9S0d4gi9SqkEite5nwrFxIYGp9
DR4viI32SP3nN6QDeBxzB4SO86ffzlWaTEJX/58ffy3GlTbiQND5p3h9FAoRIrwyz3rRn8LNYNhy
nXtu2VUe2L5KCKrettb9HIAwjlssPC9KpiKgiBkn+DNSjGFLZBuGEEyrRJh3qj+slc1HHvGRUF0U
+pT5LuVVQkGE5kJSjorHdh5sDN11f0IzyE89d3DwzRTXFdnX/ISIzO6qcReMUYzV4EwSZc9hFm3E
LWj2DfsMestrbR0tQ2ps2msV02FPxdbz3h7bh3Q7gQlIWjioQMBKtMxNTkn6THux9Ys499A4HwmP
78JzCY7mKVctrggMgsnbLIeZ2ur6OJ5AjHlRcDA/EA+5ee0wPIrSUxg9ljzfmSovX3WZ0eJHtR56
upEyaW982cq3j3SFzbYDrZMUNkZx/y//OX0qhQw0JysqcaitAq9AoAhHx2MVa4mVcDhZDARzyW5i
1nbAmDFBLRGyhlYhmq18uoUniZjVa4PAeqvihJ2C0HoRkgfC7uyNUThUajnfmWwiw0rTDiSNMoD7
CCRK8Grkt7YcJeJ31GBtEky0olUKQ4NSJ8LRG+La06t1b+RexWYBxCcaZIrqJEP0v37QHA6Av1R8
HsHVL1rBRdnH4MrGVCVWanXHXhQ4LWj5++6RxXLSzOcSQnUbpPVebJam/nNKOR3FVSLZDfIesvUH
Ac+OEt3hKm2gQBIBGfHB2VwNTqlhIxqVCyatsnMtp/KlA+2sO11Xg5SOTGhop4j12qaZm4AJ1nNE
nMX9An5LezVaseFOeE5rsxUV407ANyMwZcVbv5WIR0It4lrA9NTf1CxGwdaqds3iBZamQkdh73MU
H7TDIZKW9USwaKa/7fXQwH0FK6v3RZhbSGpoagkUHi9r4lLvoi3DbKuPqyruFwbQwv4nPhc3WRcc
pUMSCfizr9zV/LzYbBKct1DZ2rLRsv2Hkt4bJDvUYIs+P/OUQIXL3DVFtLb476WnvdsWScLKEEa2
MlZiDIL+ZppYBchefCpsDCiRJ56sCvypOscOH1hwt78g2nQLB92DapSSh9PdAi8uHHRhsSMWOhM7
YuWNkxOG58ItEmR9/tTsaNFLywNVEYYm/v5NslsJHNIXlB7YIdE0RsUg05OQX+jHSPEGw1GYcyjQ
jZmFCjeLUj9QKt0Me/ADiQn6KzHXdGfFd8l6Cs4bCLp5hc25i3UID1g1hD5FQOG+LPWStfGZiTkh
YlVCyARc3izWC+qZjVgcNEChn/1apWuZfafGUM1+/f41tPA/Xu3aEoyAbWnsATbHNOiCV4gyh/kZ
U9J3rbQsrEszFe291tW4LyLJZeCJcLUchRwqK1uhg31hd9PofJqoMjYfLVC0kzUByx3sct0Okpxl
4IkbeVo6sxycYnM0XSvmv7yHUn9uBYuPj+2ptg78mEK6AV5JFizUgToWBDFMrMWu1kgtO4Ptbdlj
WBkWkU2u0D0zxP4bmKrDbv9LaQM4YsF7IhuGaqBEVEW7fScQD6UOypgiu80jttIgQIt5cjQnKr6A
ivXIXkBUIL9pKXL5541tB7a5bavKWl0IfQi2pPDDkkROobUOLPf1r3rAdv7KN6IxAVytC+idhr53
dbiTt660BIELUIvg5p7sOiW/dHs5FkGFAmMei8wdoeaBJMAMdNKmUctijKo0D+fv/2D8J1Vo8J29
Yzxn2kkARgSiPoSx1L97NwiCbp7Z9RNmsQgbBKqNBjYTnT8zdr2GPgTEU1S1InH7bSz9yu0DH0i6
hEILhNPVF3156mx65lzj2ZSXbK4Vz6wAaSG7lZWWDEb0fI+oiiKIf51OT0TY+Rt/YLZCM0sVsh6m
RknWY+GLEXrN0iqpI1AnghogvgsHCNojiBOywZZ7b0d8IMWFDXAR5MUFpL2/P4vxakJCqgbY8z04
XHMsZxH+/cA4T1nunJTKkf2a5yEWfV5cYSWkUXmiwuGFghyxUd2SNk0KsJDvbhTDOoK1qLe3YlVe
yokMULybQNUY5dcWuUo2T5OZSRuNury3EowTNt7SS1iK1Fcdh7rS7cxmGZAKJV5FOCMLypa8SisH
hG2ZyZ6/W2NBeB1eastQd5CsxYGKfbvawthIs5f+6bEGCktrSnknzLMin49NM0072JIOROLyFwTp
A7hqthCMKe6CzoNBl7g8TEA6IIVwsM99xD3l10SxvD7K3218CNGFQPzqAs38KTHtE2m1jxYXhpoI
EUYykG7eT7DavAxKyqfWp9lVp6da1jLIKpFioUEeEOighJKdHgQ5R65iYMKxccTx7QKA/GwoSRkh
xPiPqXecR27IyMllR4Mo310e0PrTAG/DvdqZurQqIDi08ZrarnH9Nz2R4IAQ/VhWB2tUJvN6/eSt
PdP06QxR6znKejAgmBJYpD/tDsG1apIu1Gvv3Tqrvdte9uvicKZFSv3ERfVGHTzog0YUWDFTfYuU
XdbYoG3DvGx/QW1/L7mGZWMvt9aSFhAsEPn71m5nb3B42RNLo5EB2BVbUWHYOU5dKPrCzirqazCk
iWQut/OsMAgOVxhJ7R49Vn6grSaCmcZyKOkezNLTj/Uu5jlYiXIe2eKyKcRT8EllMi1V7MBOE3hR
2VRNG6xpsDZaDfDztYlOaf1lW5jxFX1l2pACKFJdHnogaOBhAUGCXD7rubNhZ/sFxF9QBP4OygMx
HVuU7EK0nCJvBBh9SoOspy1U0xj1MlTfgdXxmvMrU96XL6Im/nbkjp/zFDC2USmeG+FeEmsxIPZb
CLladI1VVElWkpDwrESV7vIcl2F8bTHKM2/GQK84/ueyr7qzRSmTyDFpcKUMNag4JWewaqbTEazU
msANB7zoDXXcCwebvfu5aeinUUw+INdtuz17enWHhUUwTlVBss9gHWOtnVjjpWmqXr/O919Oh8aT
l5+EC4l0YE4KIQhhQd+Z5svXZsdhiBDge5Ok3YU5gEjQNrxtT1QTnU0QXrLLG7/SceJ1V7X3mWOF
FhhFR3S8o1rhqLqaU12mzAo9HQyaoZMSCwK1KZ03/n6JWaB8YaU/xj5V5yBNt1y9D4okY/XErmAT
zEljs1wqGxsFYYlA2UIRNN3mwtMMPGaVhdbUXWY8yoUFbA8J5M2Zod8ps3gt0dqjoGjpHkhZqTve
olXYWLeIIIoubxeKQqXqYCC4PSN4irMc4WeBRkv+AvJl/nLCJ9S2JXh6KpxyQOyjLyehhQGLZagF
i0IWijr03RAiZf6QmYRp0gWytlBpRTUmnphW7IbiMRIPZmPNLWG+p9xQilw9mRFf1ELkCo679YeA
ZkEiz7My0qlKOZyuS1atSKmH2LvgTbQZsU6CGcgIn40LBdJ9msOfEHf2Uue9I3z7GhT1lsREAiEh
y6ZnLL+AGWIJaGNBkQHZ9rcALaG0MfvvYa8jDpSO75o8wqNjLGT0IfHMD3V2fao/U3F4k/hPBwQX
YnHpoL7Mnws1glED3i2UH0Wjfd9QQV+eEVDPw5WMQvImgM7BRmeasf4ZSNMdYA8Q56LJPGH+7zU1
V00Sdgv9FDKF+GzrHhFtCCU8ga8GpAXMV3WR7FK1zzUbxLpeHQ2w1BOLcQ9YUovUJaL6vP8IdcT2
8JHAGSespHwyBncVK/r3CRPBJiUvHqKTooZZVcieukL5zL2WExFBzSwPkNDQZNZ3XobEPGpftXWy
hZbNEWc8zK6HxisA6uU96ypO48OzYcEjMu6BBRtEV+2DRA5lbwHxr5rgW40xgvJtCdZ/LCzlsF1o
Q2N865rdvJRu30noKX4YBV734gFWdnGWnGpSVy55FpFtyW/mpn0yk8LOYyK6UybOqzAXh3JD52LJ
09Ev3a3gAQjyrrdlPAGDlZTI8tqw1aONAHuCGHiobRJIQSTUGsJHW6zS4nCxH8q02YR8Mo+zsXQC
bj1WFuOjPfzhH3G9FZRcFCRDRTbsxlKL781MPUKTVpg+gSMKNJSxx3geKLjofA3wSo9hDKaxOZRC
4aeD2nzG2JB5UzTF/eTcPFIwmA4Un3k5ywV5/ghYk8nJhc7NyOU+W8xjDcob0kWRIsKjprhgc8IL
SG90DFBfenz8MlJEA9+c1xES3UQVOazIKNBCC/SqQ2tWStSCAxRvVKzub1gNZiwiNscmITPY+0cz
w+SOqFAmExNU7mZ5yF8VIQGHpNzuE8mANrvmU5TLmFEmS5kT/JWSZF5Lv9kUrv9x7xHu6n9bqoBy
ZRRkgzufXtYL+zUilWh1XGq4goKlXnSUbR4QEK1Sb8jowgz2f1SBFFgGhl9/WBmKn8EtS1GR5dYk
Lbs0tnr4avLE4BnA5ePT1CNqie9HttQHDGTg78c0ezWOjD37iJzAC0F6Z4FbHuheTEDzRTQxLmba
wRaYOAy/1fSQyB0cQUKV686lZCn2v9zwLNMqemTZqgqbnwtY95dOSXkpP3srhEDBBpWq07vHIfKQ
nBBTqYRW4MDzhP/AOBeotljO2kXIGfe4Nn9bIIMViHZ8OouPdQdqiRH0+niU5V3R26bzde57dksG
wxBV2sY2DQTCsKwbDB8IZ8UsZgNRggLcyBIxt7AWE9NcvORwOy0oNKcGadYhmkSRQdjyHiBBLPgm
KaHzX2pkBbJ0tFajaLbP3VDZKzQROiB1aE24aLNt6L5ixwWYCLtecbJeTSMk9pPZvo8lDz4IIAeW
AtjUg/PYlfaTAjpbQYNL4SP7hG1y83E3OISFiaRZzKdFB90/dxa39IwQvFwCub9muGkhqClJUKsJ
QVIvIDsMLhf6eu4IXpUdKi0nU6obrbCSDwsdIq+rylVDMkBOISFzHEmoP4IUT3IVJeg21KUoRNHf
GRkz1cft3vB7ATz9F69Gv0jv333rQyaznpK4KSq3TsmEkc0SMzRPhH4pMdDlS6+j5J1iupss9lOD
2MMEAb4Aym1a2g7kOh+fe3TNjrhjDHmBn4OG3DQxpC2Z76IO2vwjiGXxuXmAg+iMCQcDR2hZT0hW
cHmlSuHdutWxgDXZcIOLA7DOnTogVGqhyK+PbmqQZVOqIJtkhu7uQUOD/MLS63tM7socJDigqC6Z
/JpCOfvnzFmmA3omYHvoSeznYovgcfSFus5p0DVupulzjiZTxEN4pMkezIAED0ERlr2h1Rc56X9S
FgyqxdBOB0jdt4cFCdNUkBibZh27cwhwvDBypuvgNVcmkM4ri02/W41lvCpSIzamvVk5RO9NK5sM
ky29jOAGVYbknLmvL3Ccn7vvPeKwfLjxBUq84BkSoO5zJUqfUZkNJvTuvZ8Sb4vD1leTl0cQD+9V
BPe/ij3gz0H2OWJPKmXwD/11UZ56DGO45iTKUsBhXQ/8/dXsiyWdpeyiYsGDOSgH1qwutwbdj4Ro
a62jtUNIgfLbAIe4tnJJMOKzEHkbujoA+3hukLZSPuCm4Oj8zcKIgsNv8bx1DzNwHkoiGOdXv1z7
YXeP7W+QdHqYo0v4kApPjcaRr9spULNQnRICLMLYPo0W2TnCzQta/DOO95NvZlPL4D86L0EE4Zr3
TmzjMRyKo3iVU9vO1/l73XIJag1K0gKZZta7fCa5SH3gjlW77ygQ8AFuEY+27YU7/2HC1z23SRKQ
U5TiOXbxU9J/ZQMOjXCrAdokeA2pb8vZLrt5kXF4SpDn6Ercaml8pZMLacbxexsJrAgXDm4Drlv5
NE/VDRBwZtboTi8FVi/K6nMsdRbdP9khs8qSahW31ndH97OhUOyL92vvTRS1Oe5Nhc14x0u1bl64
5y1YfXxXXWwC0NfOXj/bPq0te3OrCqZd/Wr1htCOusUUzrl0UeQdrMHbPWZfmR8nk3z270E0xret
us/ENoVLqUGTEarVWHaVG0ZgBPN/vI3ftVoRWujWGWi5GqTYli6mHLAfM2J59gQMKZdex8ExeYl7
RJDOjDfLOH22JESA0axXtbt1SPhUoSyWLltc3n+ID3Wi/+8wQa/XIJjayFWPekN4D1gfltjU95K5
qB1k7/YvsWXjo1XU8Qp68mYwYhNmDN6H3KX5CiHXv0ySWlEP2O5uCMY0fZlTITXLuKqAEUWOXMXM
V03+QOc/dZ3cx1ahyldL0Vf4aB0EOmGMgsZtDL7nUGP/wCkaJz+EsplLVegFZ0DZ+W91pyvg/CaM
p3euZgEmorR6umVmrEhkNvFiym+uiMMIPKbgH5D32qtwiwUAPkCAPYr9WPwIfL+rpXvMSLIh9p3V
iF0jdDYe7qoZO9zpe8lf1VwK10C1Gz9EmKWGH3LAb7QfvD62Y7UYkD+REqK7hWXz60wL4jtY7ce7
wnpL24bh3OeEe877ebNrwCVvn0bp73447ynNCXoojVWa4iZJMkwUcE0npDp3mQiEeHnGG2vvs+CK
tLAs3RzCidbSFq27iiCbCNYFgA+uYQOaDfwhQTJ0Td8Mij/87QsCm5EkfXfAXKmEAqfEn6Mnrs0X
B0S01uI+nbk60OUUSObdhF8btMcTTHg3etRqdcac6h/RdvNCwayVV5qYGkXV7DyoOx25OQO8o0dI
gZJ7s0Sg7MkV/US9VWygdK6k1At2Q280Lh3tZeBV8UWI7g4iJ813NU3Gj9u1Ce3LcWWd/KVcRKEV
OBjVdcWnQTvOXTis9vyGcvRVf/R4Nd4OEm+9plrCZczRQ74pdf0MuBdtVpkU5v52St6P18dj+7p6
CGMhLHp85U7pamYsVhdA117i/7swoqV/cg4m2j/2HIxerKOfM42xdFHUgaJe3Mxic6znhIXeghmj
Lqmvt64tYblEh537NzYcT079lBqRa8MyajYoIkRNu4e/b4KbAewFqy7A1AB9HBhXgGEdQ2sRYmkJ
EOR/fTdef1BwUbPJ4Jcu/6m2if38SKkMIDzKo63omv49JJtcLua6Es9yVGH55ZD99EBBqoCHBJVz
xZGnjaSXfnNkB22nClIlBt6/1doJyxGlEf6ZMckZHTNm6G0GKH18YoQkQ2LG0MejcusKBi44VM7i
z/PWDWqE8Y3eQdqV3ylZOtr5mPoIcsPYX2MH+2xL6vLmGwSrdIKlvN4yHYXZfMJlxlKg9KfDAwDZ
52RM2XClIvGbhwgOmGEq8QdCJa1iZxMLEVFfQ//v+xVZnJbasr1LnKTABzEF2/VVGRaQtSczBisG
/ABLqHb7VFXYKvv6Mv8mBS5r2wjCBpggxuMtP2Vba/CSNStsHk/0SSYZT9H9QITw/gjLuIIG3odO
lqIX5AbYc05pqqtF0hIbVG5Pumdib9ecVM0WQV2bwKA9BrpiODs7q/uYrZIJhjH7CCHtkNPs6fdV
wRER3xbTK1VW5EkvZSeNQifiNYXbynpLtNvQ1rsswDVanHeJ8jk6NOuUsPVHyfprxeuWx9OBbca8
Inu7CRm8OH9BDJ0KERLABZedc+x5wNHFpTxVK7zl7ly+RpUfooYzpWPBt7sd7czbEjdCVjvN1OFR
1gqJdEHFvNg9ad+WTPrK+w0dJbfkdVuO0zAZAwA4AyrExaPxbYz/p0Og+3y9giqHhs0bY/5I8hNA
SNnTqHrsvIFcmQn4m4hZrdZObiw0617+9jEG4lAdltJtMj/ox2ka89bL+QNsLA89KAr9/4QMARg8
ZRYmivwNHLm3puR1SPor1kjD9wP/8Et8VIYRutPASEHl1HfPTT3utEBTmugIqMTSNCCNA7lUQxCC
+YNpTR078pcplBERTRYEe9wa5VK0ROcWrp+JusX5HgV8Q4maHO6DGiDTwc4EFaLOT8awt+PfknYP
V4E0l0Wwxlc8/1BxIhGzp0ir60j/bfwNIHMU2CqWb5F+LvnoL8WRix1NbpS6QdIu0hO8ccEBIeW1
kmdowuSCsl288QrRoeAUVblJrt5uA7NkxwZQHpHjABPECOOuHbiXbgkEpbcKouOovhQxew0yAhGL
L7q9wBBQAoYfjTTE11P1/Q/+kvRfjYN7W2AEuUMkr4VL++adap94amf/OoskUADeJ2U2P7DKUubQ
gKPursnNLvqufKYjtOHGVvVFTat2+EFH12EqPHMiMXsAuJadFvVziUkocWCTePv0z0Ew39YFfzsh
0O4/fp5kYX7ybPplqsR4XTJiXS0IiFqdgKHEVNSuEfIv9irBISzbLAvnSwl7TY56Aom4TR1CEtac
V8E5zFX40gPIJgdu/67WjfQaTk7E6oIS9/DFoK20tmdTo6PUiAKa1q5fUt+Hsh+IXmVU4nFD8E52
ieF+ksGVdDvKURSIKyeu78oUB9TTi0Hldv9jq3mYfFPEk7Lhe04kSQwXGWLQg0MRjlNRArKbIw7d
PYsZHbvWWArvkhJglyeyODoL1lgS5VHvq1POMtybwn5M1D35RDJz30hjB+DQ5XyrRAEUbw5/O9jS
vxPW/YoTuSSQOr6GuKJyyh9wimMjbp/KYLs1PKQW4kdmRzmV0Y/vbbXKi/okpcuK1bXauxDHZ5lR
GjB4WFNhqaIU2dPzAI9160IyLd4+wwCXWe33tQKWUwX6SVT7JctG5c4Afd1jzPXVQD065MyjGRCI
6iQj1QGT6qLB5zgmLEB4SshpBh2BMHV/YjlZIjq8TH94O7amzthfjqpMh/gjNtU7lSZGrMhN2AaU
OwQTTHuYYBXGsSC7hOyV2V7NBTQx4/k+NHNekcWeCYtKkDc1B+FKh4ZrUQ5hj86ejvln/lcJK1JI
WGizbmMDmVf+FOrv0cS+xInC48lNy+gaG/FlfrPgIVwwyH/7GdB6cAel0hgcanZ8UN1HlKEAFICs
dpoAOGh3saJfAEwVe2w+b3IQKesQM08fYu96tATtikt+hqo5oZpBrr4TG7NER4OHfPoPmmMPlwbi
8yemteMff4FYBFnE5dnUKwMOareqkHVki7VCtIS59No83zr4bhEEAFpbwpffLCuAYsKS6hpHLk/U
TvQ8SrbRLElCMbCfL6EVdTfibp3rOPfAcwv6YsBREZKJarHtYUW71Ckbu6iP2W/kGHLjH1nTFiNs
62OKGswBaDzYPAUvzaPP4LFM8jTH4r+2GGDqDJjCwvcEXweY06/OcQxemvEHqfkA9BNs8B+AkAiO
B+QiYjl+R2XIIXIXdbCTdsa/0kGifzL5RTfIP9Kh4GzSIHZBr40uJjd2LwrUnSe1uzKyM8dXOzEX
8hILDYxaW4cs5tikW2F0mlywnffbIz37jdd9gnbruNVPKhWlCN9MeAf8t8gagiu6V2BzsbZp9FqM
jg/JUa1M/NHm+x458xV1IfPN/oDdMO9R56U91zYuo/1/ffWQpnyeHVLZH3DvQuZMcr4v2/2xb6rI
bz7QraP4t1p1GLmsJKP43xKuh1ND/WvQKdA69OCaxr39QOiHKb1R+WwiJ9Bav/FkwAjmnBSV/2jE
fhuzwYYTvD6J7hLl7wymEyVwTYZoTeOUtFMVjDdBXi/1TqQsKIpnikQ54Hj6WO6bZZXf0ZgtIBEf
8uMd+tHeL92xxh0eGacfDYbLOc8paIGCBbtan/whbMZmJFbyb8GE5JNhqFaywIcFYLksJ5SIfBj9
K0LKufHjwabYbPdS6et0+umbog5VeS153+CazBW3vFycF9OvzN8DhZL38qqOgrYpQFQN376LM8WQ
hB4QBfEHYbd8xAZ14FsQmbGTxwaPyYXEfJ0+MhsUhhzhUCfGb04HPcGjpXEkJLRIo8eNBjNWHzCs
5S2xtPzAruKdW6cN6D6KTKlRnOhXtaanyoCS55UaXIjnHlzD8ZuRXt+DZWaRP2nUxBauuqep84YE
WVsO/yln+TsriSrYkOrkpSKeOAE8zEQEEVubgSqO0DYCamHoZB6y/LKJv7auk2TKxJJOOd88bEjk
uhhrPyJC6Q2FDa1JxdbxUfdSoazvhhmDGyF+kDsmMZoM/DHz6O/g30bdUc3c0ilzV0oiwHyBTZ8x
ThAGbDybw+hCkRLBNiKVxs94SKK+cIlcA/pdSkg07PIrYzvTYU4ai+kqciHNc+yi0X8jN06D6LB1
EY0EYtB/3R01SqFYYeQH7cFFFsd/KIStuKaRVj0QPVHpriAkn0ivWV+zhJ7i/PJiPPiNe/GraYKF
s+syoBSZdJH++QBVhDFXkQru7zN+JOhuTQ0AuM77KrZ2pUSk1eGVNamFkWKxR/m7WOnxDJGZ1B+m
949q3G4tWaG9Op9zJvSoHdXVKau9vxgt7CaaGWnA3VAufb3Xo+ZZOPNvenEa6BLJwVP+UJ2LcsaS
kKKL2DbcH1vQt8vhSYgAJxLrAETsdLhDopy+3I9SUP/P79S+NrdANMrcQuEF4HEfgw2OzcQTClJ7
zS2RU8/Je6BJVPQ9Z442SGEBCRqn1kQwxn3AIiW9qVH/dc6jmfeQ3l0WLkhgb+wYaFEpi0BThlRG
vh6JaRtQFlal8al4+2gNpV/uTUdDAIwVqo8oI2AwsU09jw5mh/d4jnLEjQRTtyGxuSSxYniANqz0
l6MAmOc5SCAYgGzqoTNZ+tue9dfkIaGL9z6hbIqByJBWocj+we+Zwd71oebyH3vsClbgcjsZ5VBm
5HK1SkQVuMp/fT81ZmnzbaTxSj8UHQAbOfbyAR88IyyzWfdtlKRlmoiMmVNCEeJtYtNAmZf5CXMg
QFshXO792JFLIvigO2W71g0JcF8lg2+FOQsD8AU/GgGOqqx0qL1ZFaP0AD5xNLKnoIfquWdFm8oI
qcKf2/z+WoKSyo2ho3ptPakNuhvHXpoVEym5C1o4ZqN/T+7F5SCleWhToy4bJHwV4rtNLcrDr2hj
jO588J3cSNlvG6P2VyQrO8T9lrc2gARexV0+lFQpaiOcD1pVvn0q7XzsG7sPUqZnnc0mJGCvX5aI
YcjU1mAZS9gDoXOU2Q8w/kNNceBF9WLfbHgX8GAgakq7kLET+QZxa8HsG4i+lizLgSqumL6ZLm5n
kIx4Pxt5gPWmZp/451ieuQDSZmbgJz8yBYBzLijvROH1TnWi5PfSemxvEiobXauvctPNRRoVOlIA
3JDeftLeDmI7JXqlmUXgFpHjcVPsIupqX20P9+3BtyJ7eKHvqRKxXiHIzCXbq3J6jPBrXCiRM3NI
YAZ3IQArA5OjjOP3YGrXxpSu/DaFT3aQBrKL5ZyOaNVe17Cc+0o99BZLLznIjLgAQ1AqLHmav+cO
jVREJqy684Nf2bzvG5ARZRQJf6yF8fBUvR1P8H9B/6s+u2xAbAMr6Mh8RWB0zTQoF/lMq6vgUR2i
FFAoKChyjKboywiPvWO4F3qoOCh4dA35nMLJ8OT0YJcCGZ+Os1yw6bF2x1BmPf4vltrB7/0qNUGz
cuZfLf4Ap9hQ2nNhqHR2VqptD4XgVxU74E4a5vMZA0N/4oz8R///VGDmTURzrqnTMAoORSw0NmQs
WDdvrSCVmNApPgKYKJxgvgR3PSF/na7xAxM8YScq6T+eVOB0SVvKyhWQrrlXeYCF5UMwFdux/bA/
AQGMxM3sF5k5BDi0rTWPjKC0+WPdaqsT+dn+xMsrMyMnpkg1C9AfCCMQ8q9J0K5DbHE5fPbhK7XU
qcAt6cD8Yld/h/NWoVgsDqiX2+1C7+0fQV9jZ+qgmq15IYfSV5yE/l63abq9WSB7VfzdkMENfF4U
Ozth824LzMXP7au+DaQ6VrGpIPOhx71OHkCo0u3+0LCPAa0qvGHS2vxwtVZfsNZtGIEvvjvguPyJ
IVg4ZJGgHGEFnBZ7jTF+2sV/k3DmrQNkwi6UMK4WVXVbd+1Jgze4bmNTXT+qNndmPKlENvxerEEn
7hnikOuxZsfLsEinZlbs23NPzqU4nORJhSr4YUTXkTRYE0TFXvHwY4xwDoD+P4xRJqjacIYqlbBr
L0XU+KqbvyYG7qiqT8dIYZ6e3yiKjfGvZlYCpfdQwBtEpjcUXKrWXzVuJPzBqMrIQZNFsG13kYuW
2BX0z/nLRCtUNLKC4Q/Uk62zhs8uKMuU7MHetinIJkQS7sjYJiamyEU03EXAPBiIljEqp6DKwD7R
oTOQJFDtjt7rgdKZxgDztyZmCdpa9rse317q4KrtEE7mYRSiEeJSd3p7igJwurIEeLc0IjO7+yr3
8ORan82J+HLamvj9tGLezBXY5xvDlor+N5eEK1ua+EkZxFeUAoOIwWd/jm+QWrMJ5ixars+Nwi1+
U+JKNA1Aq+vdrY+9TacxQ2TDRD2mWDpw9oVOCMIF9wr3KJwSWQypDRUM7yTBafa1cSpmyQ0U4Zsh
5dyWcv7Uic/TzT0BIdooeekHQ0sZpedGg8VCHt9QDs8rKdygVT3TpyuLC9bsdPgBO4lqM7nomR5X
10CCYIc444o8Yy/3Z4fhSojhQfE5iX3UMsMxPvBgpCDD2P5voS+YAuT+JtSP3l5ErJFkKePtTl6G
SJ/WDFgzXAtsS09Ife21M7hFAPIFLRo7kRkPP4COwDSpdYmHF1B8eSIedy4NIkJ4/Z4v1kwjmnm9
I7CZ9eUDJ/tO+iVo6cxLhv24w06kTz7zDdpDCuhKGwuOul5++mNOog/h66bu22ap50FUqcIZxVrz
tSelevgLHt5TUEqPgMIqnP7lswM4lvT1tTOk4suMd4/eQZcFFif1ie9Znj1JRUicLaVLoHow8Rt2
ZMNNr3vrTRygrqVz+Ex/1sEZMpV0IrOgzFqZf5pIUzyIMGNo2MkY84EpR29VZR7HbUYJN92mRfNR
2Depy3mD68uK+UvDWWdyQ78q8hchLde3ECCAo2/CHZ6qpvxs2KZAFXWqWCnd770GR6jyjFiEgyu4
OJ7Ml7oHTa8ssgiagOBCDIbBGwNbHJqHFmcByX6sll+YAGkAYU4jI2Ar3QevKj8HOEAJTTdL2wPe
f42E7vLTsMSLCeFHML0Xoq/1Ezc9jV0zaHlXx8RfA4UtDXzUCr03rjOpjSus70WJqYYpxhPQUaeo
AZE2tWOMEMYum2Od/72IVqZzR9mlwC7DfUtZi+lXGzTWWC4cFjZoNxCY+43NyCUjVnN1oQDSTRO6
W2W7n5fv8m5MzdeG/yt8sxb2DVExCsmZ9+iT5ChIglaJnixt8hXVGlHi/zoN32Cq1WPfSx3AECEo
bbQktlweKaUwDhva/3cwu2uFRPykAv1q2W+hPCTjVBAuRqv2Y4hcvrge4cwH4wQsgMC6KjpgwLEP
qw2MqjXRITn96Hk5x9mne0nbTcKK9WnV16I7IDSCUXBtJkffnt2+voMP47cQWxt5o+m5VuAqc3n4
wbLhW8UaqweRf3kGGwVrsrxZTFXbGnRqMXU/oYvTbrZ9rpKTVQ/xiALQggJ97se17us2RRrDYkSt
DAHoiPDKoMB8oegwDA9jCA0gVmM4NHNKY+Gb84NMYTH2gzBmd7Hw9hsyXEReY+d1in5QbVD3XssB
1Dj0/aQM3d1t/RaqyDz+9tQIxj/AfZ0QWJGZrBB63Kp9EgNtPflEO+k0q3/6QS0Vw4yq7Uk6GxzO
zbfvbYzzVrBSXdJKMlVlvZvjTIR7Jy5Nzn6i5j3L9WqOCP/vBoArnXw2T9eSc30RX8Jhr8zHdQfY
WG/QQsu8TWAHjWJxtdIbsvrSFVX3VrAmAlvH7C65fdqO/M0yUtEZpI24Btm2zXgSgo8Gv5RgvW0f
B6Ih1jFcfCFKhyMmkOAQZwhn/BLud/7ERHEda29y1SZ18Mv85QnLyBh3CNE/1GkEz4+4HoqNFZke
0HIFoyVdl5KCowl0ohyciaIWAXZ4dkeB/RTP/vc/qX8vyCFl6rcTEz/mVXSKftmir1VVbOKl4wdn
zhs929bbSefMeq/FCEa6EudDiSAePHuuYXpN4jSZtYCaL8s3IXxOrwCUyZya/dvtT177V2wk38Jb
fzlx/CvkhjiJvy05T6GsIPkZIKHAM87/UyeOaqqy/m3tcCVtb3f/jHEKg8EBp+IL3cZfLzhPJJli
qGako6g265Lv8d5UcYvJPNF9StEkP+J7II2QOWXWmTV3NEZaQDUipjyvnvX3ZNTFfrbnFhlJOB/L
OS8huAVJPx5vXNP4O80DVvBn/ov75e6pSf2JeWCRCU8lSUvA65qK3+Ho9F1XHudMdMq1nu2Vbczg
dFb/cdu1kQg448H4vHH8lQaT9BMNtn7PrkypmGwHggDqI+GQnpln8VbjDBzhQ3JuwIy4cLUOu1Zy
/VR/Gr/A1auOJxUH/mHacoD34k22rIWUIWQ69qYqkzzyDQDBC3ahajliPxzC3A9oqWC17XAwSdqF
sa38cCX7SK83S8qFBUMKOI1SA+5AWpiEinTf4TuAz+ntlArIOJwOoo5ymFZfIkoG+eBaJCmE9dAU
cn3+nMpDRbbUROirwGj5s6S4Go0tdyx0/+vlq7qsJNvnBbT+7jsT1SEWffqnN4AnlZoq1DFOWhtT
kxmV0+UgM6Vv7EMRRkgwEi1W3oiN7ncCaDK7yJ5eipwvoWY1IXgrw7pjKx5HELnty4yaP0pMyqvQ
urwJgIL2KNSPpDqIdU27msimqjQH1LWqWg1yxtDW99k0Q44Zd8c2PrLK64gIbRSRUZfyIuEXv0FH
CmE58bPR4cfFJhssnxhGCQ9x721dhNIACL/tOqX5mirhDksk6Z1l+KgfdGdh5ijTjqLkVpJa3Snv
a34Kavrmv1r6DUulzCa4OleH4adHTg/IXlrfPE5jzXbZF2qlKq8YLN+BW6DKLvAQymfjYWf8p9gr
0b8HjH2mdtcI1FyStWYR19Zq4h3XXXdLKOPAk/wB/B7eaPeI96/z9s1FafLYiw02T4cHF1N0SVw6
/9LXgZsFuXsrqtkXGZkTXb/V6RjN1tDerY7OoQA4RHuz9hSZeGH2AmUVJhmzBDCIAgtv9hQltDcj
oFrwgzlqiF9eR9emTYlaiBR9YxvSlz0DEpLSmP3X8bzPCBVd1xOhYKjk/rU4VZUogVkFd1CeKjZE
ugKu3F6L/lgJZ7EalG4Q2hGTkLtXoK4Xm2B0Ef6tiynfYvHydMPxsI2ecGIYeM+WUi6ddaSgcBG+
kpVm9jADvWAVI5EYiPlfnjZLZzcXTHw3BGHtKTIJEg3NCpnGNUlaZNpIDo4iJNWZcMwo88nF9cGH
shLfyjH4OuWDB9oPZiKEMKMjroqaFLoXfa+J+Tv0zVuaal2dTAMtfQrnU0MjNjy2t+9V4bFISqJ9
vwieEj7MtP/jQm7WwoeA0kj8AGuqzM393hHzktnMjKROqCofx4vtO4oYYHvR7KKRJErTJ6v1o8yX
SrvGG2vADNXXLt+NaJJ5uDo84CnYGtOmahJ/ZW9ggqKhmDLFZcUnI8rjpgWMfQtCreGWzL+jzann
1LO6xWlNwlv5c7GsTUMZxnFERSgU3/T+F/GG30YSSVifx7LbOfFx0vMN6EFmTAtxV//r1Kcw/zUY
qzyQNbK10XONwLYvkHi5KoNb8LSTCFEhhg/WacyA5JR6Zzyklmur80kHILNI0xm5cQMSRpfzr58g
F9oq5xm11uG2LWldisDezRjTTz+BOnH52iij1oA7WpMiwi6WIstR0nNgLaT//xLRayr91wUzPnUC
+qt95bF3798RJcMFjR8BWCwAHWXYuDJiSH471+HoYiezrRt5+m4XskGtwjB+bq7yRaOaYsYX+kQ1
hLtjEG1rgAbFZ34GhO/2MrLYnL9MgYqyElxtKkb9ZwpdHFREqRV8SGj0vlCyuDklzY864+ivfIXM
6BZtxNDrVaIwT+5N+Iw2U520ddRt5GuguFHfP8z5YEkn17+RFGiGBxq65kALwphUI9xFlASsD1+V
+sgny4Q4BFPO4N/IfPuxviNV8iFC/VAZ22oybqQafwFBdzjRZZs36t5PL+cunPLC6UKU2HHmDBD8
7tt/UAyvAQqN5iED4dMbuRQ7sIBXdfYM7oujNMvChQRh9WC+aQv0pTVbbQndm35NRaaCa5OY0YsT
NuW7nilGwbWG++9ydcLiDxNlnI5ygUIpcpAEWRi/ZAXRX0ZXUIyJdwsSWkPpsd70NJD9fMttWJ1r
Y1axylj+BNG6XeSTGzdg16oIKm+xmO1Bpxc+37mjlCXB7Ea2Pp/6hbs/WEo3Mopo4mFqXTD5JiZ9
wP+U9TeIIJKZiObCbTbNbRQZN3kzJfJotQfRPOMi0EhFZizfclHgsyTygeR2NNH1Wex2ZWvONJcO
2xuSd5gI35dQ7I6crUzriLVsxlx+RjmPwzb3zd9IYpHHMHO1XXZ8pzrs5zcxagI6+tFs2efjVPNM
vUf1FWLzRx+qkuGfqsT9Mw8DkAQxTf7mMYAG6CeEc0uIu03+h/yVza/uAT2IrZjeEKWLk3cuzifl
i6Zxnyd9A5ylO8TSY3e4Ib0scaaABG7fvF+5utwACXd+piz6X4Y6qo0Z6vtCB3W1L5s7hT+lLNX/
nx6aOxiXfPdGg9KQxB+FenSegW1qEcHgQX+4/srChJZ/uUjceO0sDnRol1qkiqNck9uzPx237kRF
DBoQUEggw2E2SpONbue6wX6izW8MObskbF3TRDtqFZGBO6PGVLL6SLX3vsTAu/IKVGR6S6T4aXPl
sGtmmtHfyrB0ndkKDqPFXn6AkjZDbmdWZx0SlfhWu01nKB7cv3oVLTrhb3HBKA37tO0Jayi2edSa
g6dVCTmo1LbHdIwx+dHW8AScVy1VntWjZYgBQ0q9lAQIWJ/Icg8MxJSyIeOu1NCBk+40M4wanOLI
o1v0ZOM666sU1CPwKUQeluSzpS3eDSA+8Jx7rdbedyj27ZJUKSMFp6bjYISXgOEHPbwO8NNzMwXU
5GdXOSm02jUrjrMGxn9l6uUBewC0edyfNo9NTZX3p/LPc4ZxANAVLes6ezkdcHCOSUZVfpt0XVVX
VCLOnzsWDQ2N2Z+ht7RDVd3zU1KMdz2Fybrl3vSk0AD3sRS3UanUWRqQEnBcbVwAdTOLc3EzjZY4
hTFlQKhCS/HoYbIyUU+E6+0+6brVZUWLd/v+skRhutlEpcGxHAGeo2kFU/wrPPAwczw8mu/Rz2uq
FcJb7klleDu7yxRfek46vGmp0SKitx6bOSOwS/VTDo52Qu2uuzDDEiYh2Ow73LhH83X8N63FLYLz
kLXzh1AAiLSwqKt8sCV/FUeMZlh0Qf+KK32p12paP6whZ8baFZkEjMq1D5FAl4Pgp6DJIqOtK+p8
ocebF4iDLj7Mu1UZPa5tV/om7GNei+bEyudVJiyDpl9KFpNFUKxrpHnxgm46oF9iKIwZc2an6HFo
3/7Yc799sgXmm8rX6euD8d2r77SFgcpSlinvVMxQY9NiOPRTzATkLd0Omu8arNcV0I5p6724Ceeg
OgjAugz3eF0CWktQvMXbSPt5IWOCaazZzJTAz8cZ02ryosCu9tKiGTfJvVzEnLS5mkxMecE7grTw
U+XW1b7heUs2tkGi8Pzwc28xQ0mR6GlnWBftyhc0vpom5OtpJH/kWlqY9NuF8fLRytj/M3TKFRLt
GWIwejVGHzB1eaGUfEZxlNspfsZM/6O5gUt1pUdqgmyRihcJOyf7yavZrQH8+vcfxzp30C2fX4SR
AXAENeUB+1PsPtOsiEKOhPDqRacVxw49Av4YjrFegt4mQAGsUG/rE0yhwwITRhFWom4YdaOswCHu
9kxmOqN0Dv3kxrfZeA4D1zwVUAu4zTWYYC/k9TDabIHqPYZgvYkFMnyELz0V8bw0chMKoJj5ZDpP
sQoPcwC6JtJj8HiMVoaoULOxqx7+QpQCOMzCD//eze10VItnVFUlTZ47jFYq5IE0U8cZcdCz+8SK
ysVEdojR48qigY2AbRRyREL2pI6cAg1dJP7+ktEShykJknwG7Uwf4/2Sp944Y+1ux0owcf1tEyOf
0F/YksBB+xzERuZaZC1pTchFVX6KAYjlDv2Zbz6+b7PTGwmDT6Eeih0sF0G/Nh2+nZQqRwte1cJP
ncGEAxAD9BAOKyi+wvl8P0EYdYEou250OyvPW7bQmpVGmn+d6Mo6KOCx3u/UyTxAmhSCQJL6viPp
Nb5qw78+Y9COnM1e5kfB+R0PC0GfeWQU2E+faECRvIYBGmlOqW0kCpUjMLa2U2OvzpihSsVMWDxD
mk0BD/iCxDB+FNvEoWnYG/VzFuHQ3j+UdUXPlk9tFT5DuJQzF0h2tBBTls+W98jhgJ4Pe+IpEhtG
bdoqCb61vTl/8hJA50KbC6/qVBD0MeCtmNYMHYPpARYRd5vjIWU/JtGeO2StOszVBbxqyglidfyV
QvnBGmlbepVfxtxd4v4yprm/RVYJnxSbN8JKsN1ygY0xEA45yk5/wM4Y/GM/Gymd3yJ4thfl3j8K
3vSP2py1P9FPj8XhW/X6iNzPmxjtd9saR6kFlYe1BHKPP3qU8u/s7Ol8ZQOia5icXLYjx1Or/xEr
ezofiWWONdrkZd/zD+QQG6lQ0ahlQGDWuPHbJlzvOVMkUPT726H1OwYGIG953ge5N0vX1IqEYYIM
vGtj10zr85S+Vqg1DsVAqPbRZ9YtAECFbjVs+tYNyVsKl+awXH1qTuWdvAXAxSmZY1LptAj3DubH
wyU4CGOEkifBP8z1zgf8tHbrJoYtFqh1F3CfgaHAqPNGcswOeiiuuK4XJ66i7ff7wz+dg6xjM0NU
qDi/Nhb41RXuqI1Y8ahQLH1HIQOM7u0JI5OWXeSN2FsMigq/DcgRnWGwP0mwRzouKrGg9Xsvb4sE
iVYpRoWFx3GrTxRyVwOiDh8HG0nJ56F8GB4ru4o5jEumpVhU+nmTOWxElJgP/aj/wGO7ZReB0xGm
XJBwB7UH0h/No+SDLZisY+a6K95fdV5VM8TPWE2aCcO9f9y8euIvhZto27+b27qpJ/3G7/2t0U7Q
775On5tN+qxt/nVaIx+Bgllf7J55vGKdI7Z/MOXHY1gZE2oEXexXgK0+JJfEn1RVzuPcO3k5Kcw3
dlUVPUy3jtEFrojriUmK3CmeAy4r4lL8fClZejLpnh5oT41w/NkPKdTODQWM6ULDYsu/hyDm+dWw
rkcK+OdrNvsW3a1gX23Pw81TFaoz0EUjdNIT5WRfEFL8Uft0K8PUVyZW30nn0+TN0qn/G+6YEbxn
tA0xgE0QY5ypAbbvL5KYWgIDLtN9pm7QE2Wgxf9dAtTh97PA7EREoxhoPMacz61+iA/k8meTO2xZ
gSwL5kT7rRaoB0iBZMjbZoVzWV496t3k+nUEZOwMfV3fQ7NGNVsmI07+908GC0wFKhArDgO3scL9
80Ae5/oI5B+6LzvE0FOFr0zmAoSeKtgk2e6LHLEA9zOsqehKiLE4IEXgpWj2SOJ0eRoW3iT+QQfu
/IR8g4BHzykxqwyTYUrLJyPYqy6C5F/ytE/qrbQEBoEOJzHUv3gF9dN2xaNRa6YKfMxI1GFGOoV5
YjBcgbkk+WZJwmJYcBP/OaGl/W7qv1cqCEL5sRq6X+DmeQ8ixm9w34XWNM/NeixiYqlfr5Ox0XwJ
DKZ8jZYZexuhPdFE9v6cl/C81nltcJ7i4GSIJoiLnaV/eoTTa9QciMRdZDCuIFDDitbF6cgfZAgM
VIiCLpJ/88DBFarsX/o9PFdt0bnqct/9KW8y98ktUrbuCRb12gZXosfjpJydYHcI25RUvgJ56EjO
FRplxQv/KRq0h1lxXk9JH/YDLNrh00F9HMIlPwGGco5EkU1nYqakUxkxrSRxmlhX8nvwzmdAj85V
W2iCmXG4N5gW/tlwE5BxWGUjaaa5oCGsgV1R49lFw6rj/wvhNbuokz5dem9XD27uK6froIk/Do6P
dsJfb0U29mLzeIPh+KAvKpNyOFmzzLzHKMiG9na73U+HpQ0FXrPiEou7Gp9YtojBiMbhmOPrnM4j
4eEfRhZEbYRmjbximx1rb70v8WvTBlGEy/WWlYcH3lzITe9H/kqfNVKgdSthk6AmnhJJ9XZB4R+6
DF5ZHnEsxEeJG3qP2m8lIg2yIBQ2ApCr5xMwiuhV99sh5oNgV6k5MLQFoQ/vfa/px/jqbjN4GYnz
rxZQypSov3CQBRGy8sCnMHBNjdypHqdZi3T5ij2YsmN5D96P5OjxznckbkD5Y+nI7JzzaMuLPbg0
sH67EqGGgLSUR2S/Ti/LX9yT7rryL8fwloyLH1f0AmtFG5zNSU52TUqrSoJmmw1+Q5Yeo+e4G0N2
39HL+RDs9L8zHg/cxxVrxLosdCfmhhXbPcBTWIbQqx2HlWei56SIAam7iBmH6ft3Pyt++jLbfRgq
i1G49tP7CEgIISfFwrXcw6PwQU1J649ryT8Ukm5qd7izvBLJxH92EosOdt5h79NBBSxOvN9uXk5y
sUdwVVzcNFhMWPGQxL+9XggPuf0WEDgUb6ceeYlagXwn8P1klCmG5fwGNJzId7UWEDYD8x7BWgzL
n6+g46CqElRXYYc5ZgCjJfjWIt4i/FNhKhSf2dVJDzs1eguAMWoqOc0sToUoxpVKyrKDe/9U19vY
J/LspyCcehfMPC9ZkQVatvXidkhl4OdCs82YamW41YBiN92o3DHOhrSp+TtBp11y2IBPerE5WNF9
gOcpxDjnogQo0FC/bdIw3EsroT9GBXxsA6q4uFr9toxspYL6ELoqs8shYq+4WKDW1fwOfWOrUEOT
voF1IsgrtcUQciVYRgWuOvkbGoPfX3CHQwU7vqv28rwj3kCHjnu6qmLkf0YwhckOvKYsZnUr7rWb
VdEpXM51s5Cqp8Sl07K40Vl1WgJZc+mjh9hRNAC2zCNThwVfDFnX++OXvEr9YyXqjkS0z9oWjwv2
eR+qupKSZczSSpmea5gHqWeEp3cSuuLy29zbTccICGuYgLk17eK2e9NBkH5Pqz7fnhV8KdcmP6nY
mZxopQQnfycjjGiIfxI4a3aIsgMmkoU+fOXyXVz7qna49rLdyAUNx6H8o81Dmpjs511OKXBXmykR
EnWx2M8MVYvesCGEqG+FLrjJImfEYDTcu/Inh/QCPvkyCwJ7l+rvCNz2H4ky3m4U0YXzgSXLw+oQ
sS7AN/Iq5bGBUoMssXrsbCn5wqPFY6g3EcJFir1bjt+K8J1CMThRBMOc23NtLDuNgiyNMxtTE8su
QnOJeivFr3bazXNAQTTxwWiurxSOH3cIWpFzQ0xSrwg61Kuuis+LYb8Od7tNSocBgd6MRaU/grLX
8wCnWn1EAufnONa+I4WWfGcFjSccJq49hKa46NyDe4pTKpG95Jvt9l2KkUhkS59IbZ8S0EkJtJgL
Zj7Q4nydDilp1GwHjEuIvTVYhEAssJ98te0k0vXvNa+ZBq5E+KAVdsFZCWbJAjsbl/p8rKgkQiER
mbG9n/R1tUYY+cnvr/eK1KE7uxqi7lpUyVtbJ3ApaQBCYesvqE0SkPGAbQLDHOZMPsQnOUwbfU74
E6sp6KaC6GOJRxNrRexDc9c+fdZ2+/RRqCJEhBYnevzY81fW0MGph7LPcx5S6HH2vf31YPgDeeov
wJTNlJv/PT9AmXiQQORD9kFp/3UXj3hSnzTk2K+raFyTmcb/N7xwIHeGOuGykdnM5LV+kiYu9Opd
723fZjdyPITAod8a8scT7y4xpZRR+enOlAuhkbDdxZG4ZV7BUtbSpKzmv1bufDr0IJ2xaq/tSR5S
XHAuImB5p0IfFmIKX4WUOooytA+uBUyu1mwdT5PP56rGIsKcVlKNqNxbjSJdorQHengr9j5RMqSQ
YTpvh6EHDMP5MGaJXgP+Q80hEio+zVjqowRojKE9xs97vy9MNPCkLtRi79Gwt4AcomcEjvHXBv4I
sFTSud8xf3RGuhW3qGyv3sbVh6gGr2cKcWpRy21m9xJlS9v9yPlks8ffl2rloGr3PQoBm3Yl09V6
KBd+7HJBUz2aMmIP+U1Qc5GixGLo1A5q2TGYzQNjOC+MPgoHEQTCc4NVsUdcQCw7itL6Tzk66MzW
7Rh6QWISO1Iu6avHh2bRN01yOFTd9DDdTCyWQ+qsVeDdROB6cbkooAxbuFFgjTor8flwwz+xAGc5
4hI/3mM7gzq7ald2xQm0H08aKJEIkV67uTljFTUQSWKaU6fPRgKp5Z86Fs9Kwe5A8KcT2Dcu2z72
BymIRF3UBeMmsnLGccmUIiSTbhNftjDhBYn+zxb/Y3C2FQbPequ0QnxAKea78g7R+Z+On7vvFyMG
+5+XiyUPu4TOPwu0YBbOWzdtb88Os0FLHtkmKvrx6RyNNdKKS2OrlFU0GP0viH8Dv8lMC05DMXPY
Mj+hNNtkoW51QFyOAI3XsAusgWn8LETkYXPDJosSzkHd9aEhTJ8Unf0oT/3fvlg/oy8ZGT52WauO
fwdnMdj4cCy+xo6uj8ubCPhfQiuyVuKl6yfwqYI+kUz/zzEnyehrntzKDJjGEQVaaPRWrYNxysgM
vrvSAUqoJV/Qp7DsopIgaTT7RJeKMbWzcfqjXlYLTaB8CnAkrTJkRW2DtgHQt1Zfansl/gmbqFtl
LbayVkJoagjxTvaQBytXyiiFAqA3AytAZpEBhQmwsRr5dWh5Nf5EUib4rzUzRbgUOyGsWieY54Sm
i+KIOs207S5j4HsOe2nXrfIA2CSnv9CHOYtiF70x8Y2y1MZJMBacJjhUL4Qw0WC0pXqiJXgjqzgy
U5TISjNwq/GkXRkrDbaAro0td/wYxYyC/+qyfuB3xpXQ0VMP+lr05Ogtk10QFh67olcdrIT9w9Jf
038VSA5X0IYnxshV50Y9xzKtxPOOeo6LHW36Gm23cJlZ3PXBwbfcrRXa0jfUhJW7+U0LViogxSpZ
rjI9qG2OdOTIKIz29wHlUiAWVv4lMR5im6O8P/anahael7s1gJ5nvqjHKy16a4NbKRvldJiAi1+m
himYH+zpi8zQhldjy9knnnm2BaazGDK9YVXBIk81+EhPWQnYI3/2r85zukxI+Dh1quB2qB6fH7dv
GV5Qrp4gOO1HT/ts3MbMx1HpanXm5pfeNsD2d77sLLCihznahkH7k3qv4h25LZhAx+HVH944abed
Gagu+gCqaKplASYSXEG/sfWue9C09gNo7ycJc4CUimZu+QOShDl/cgSfbQYjWReOPRRpm0V9Xnvy
Cm4adLmYftUx3V76pC7jytNnqGyipYypN0MpwxgJkyO/m1BvP2PZBvapw8nDW438ovYx6x8KDEPN
DWyeBpZBqMSmrKrdyFni/sDpJn4U+SxHkFLph9r2PGl8lrYj/MQy6SOKldKiyjGkspqWzL8C+IBT
mPN4+ldK63ZJ9zaTnEOx17SBs6O5GdG06nphOWRZucMpb7HbB/sB5Z3trzisfwMj09LjdKTZRi8+
tQFr7DDdxBPEHmkN6KiPmMzggUXDnztPu0kBB1GTFqbFFs5VtkvnScb6I8U12Li2sLxA/D18IJpb
6WBJp/TIFef6CKrCo/AccDgfDpYd2t7jG8xgH7x7eR4NIxesN77KKfJ5QLZEuEEcMGXt5LZ5ihSB
nqV/63NyUJy/2tcrEzZYLjHFqE/N10DBn/KTK5jWhgJh4++z2FBBZQM+W5Cf8m1hUpYaIrJac2F+
tlMwXe5K9PvNfWteob4iDJKXrABg0o18II7X4O22yRyyEq1G9GQAGWTWsMCcyiBXM9d8/o1r3mOc
IeQugAIXXrRoLdpAHZO6LOuKxkfO+ClSy3KNczrO6OfuixAd42hFeNKJ9m25XZjb0V+WJ0MH7yKb
vIDbitOXdTkVF703nsM5xJC4IDMKH5IaS9zrlaLMyzQ0qfECirBIz03CAPvQh+Lqq0/FBZRIWcM8
7a8DRUFQolsYGfImFlXfDPqPK7xQ5GyJTyJuaTL5uaJxyAXaytfNKvcYmVIYAbqLkIR/pQ6plVVk
eLVFxTJsVdX/sRBHxZTgCT9f7EKW03RNwZssPgjassaF1wTGsrC6WdPA8o+gq4yAO0/ghmyu+vMV
a4mrvnHX294i7AAR/RQHWjP3+LafJBm/bohyhOCvjePftybSi/7PGqVbfFCj02ltG7XBUVMfQn/J
YQAoWjvKXs2dSGCPUR0ev2ngEinxGpHWpkrwGl+mcpRZVfwax4akeTMHXhZy8TlCxRfLxYD9MtAY
BMn5JmB696aQ5syq2RTooV3qmVa0HF9okEk4rvFiU5trZSlVcNP45Y2EizzmfaVJTS6pFJ+A2Ol5
f3VpTVIMsHaaHkNyMkgqdd0qUbDdK6/KOH/uSY8CgfyoEZT7ujG3gDimufo5WSYlObAXVsNrTINA
QcEMSmJT1lOT/9gqhenMw4jr5wXEYnVHtOwRWv1P29s2tA0VJ9zWiAxvRfhIUYyMDPyk2L0WY/0t
BZAnoMaL5zuoxEmz62OAXgu3IF1b378ytjXjFTagoeZYD/nX9mlhA3Z6OQUb6nBP8lEpA9eylyaY
9OeTn1lkaLxF2lKg+YmoMoUdR9aBArVqKN14lbKC+Uuz59O22lSitueR4YHhGzGwu9FBJ5jdnhck
w19lxg+E0V3X6r73vx2alIPvFYQ88TFbm+Q+nCysWWf0f3tP33S8FhHuAfIAPFBjmy0yr/biaR4r
Y6szhlNjIf/gPJU/dpNsHCQH+alMJ6YgzKZKsb6q3d4RpeH74Tq/Be2XQhI6T6yvDRC691YqjgR2
xsLNvVNXnLmOTmWkIpBBLOocuXy0wggKn3tUWQK4axQey21i8Wy+vZYBaK9AlDaxC6FNIQ9fhG0A
3/3Rl3A0pu+W6hrtWXlYZ+YiGfvjhVaJy+sFbSOuNPS+MWJb8EgBEUVJL41jLYpklpNUYk82kNW/
EgyFgSj4xxPh/AIdCKuyjpweEtBkq7gC0fI1vgdB3bh+F+iXpGz+/jZA+l8lDYX6ZgsHdCA4vbK6
yq9s3RCNx2TJi33iiURYLJ5RzjqGj+jqn6bCxdpfDgF1p3CSk/y3o60tErMZbKSslsJh2sRhudzM
aVUDTYHdmb+W0gthgcn56Y1CLKu7XKaS5gDev7XuI7992J2PFH1r5E3k32cvxkG/quyY2aJCyMwT
54TWkL93trYgW5nRS7Gb/HwW9gXWj4Whvxc4g1ZmLca+IJowXpxipSlbjcPO7EP9eDQDHAt4c++V
dYVNzKfPIatG+G50rn5CJGKm4EQmKnXf0uhFberlFNr6l6PL4ITrpJnamJKQxIQ/ireoXUk8kBrq
qHzmg9a3nAOaG4W72Qvm8LzY8BsLc52ZGmH2/Ql3Ru4+azpP6s4KWY2uPD0+QGGi6Fs/LLHjN+Cb
fvFAFkPqBXrM51yknbNpSKnR5CiYuNNigoNnP+B5pVJSlX3j2VGGBidAdv2Bk26ApGQSJLykxhu0
fpysiJQMmm4RJrWafsZV706WEred7jSmxILFdKjC+1XaFuqualxUkWEbix2r5MvzDn0BG9K/UTK4
ugOVZzCfK9WbcZGTrTH9kYtmMuiFjbbJZDbU3lPSNya1ovMDMgUn73YWN3yP/JTz4QzpvDggYNy5
hb9rQL3dRzPTTeHCWz0UxxGxTcOxhJu8SNxquF9YI0CSVGlpvhI4NAtDQh1uwZlgp60ZFnhurn/G
aJxTixmhQ0AoyrM/7+WuU21L0ovHWyrhHNDJM6O9zRYxjlQKat44+zRJysbMq5GtrdeLszwX/TLc
+DZglcVRT/FczolcV8CrRa3Lijzal0aVSRj4wdi38X3hCaunnvU1481XimdtAA7IYBdLCL8Rt9yD
D7iQwD4SneXy4v6UIbvxISZESpV2fV7AP6CuVxyfxWH2gKrgIcbXjIJMyNRTd7LQS5HdG/oi1IzA
t/ZolFb1WivFB19uJ9z8T3IfWpXpXxDw9ZcUFBjY7wkNlQJ6vAX62AZ2omkZoX6eeDjhmFCJW2RC
I7Vq0TQHz572ho6YFs1t6Qp5v/M2xD+LpA4CJa/htPMMFdEHm3qzEgA+47FLoi6e2sK+qoZsgTk7
YpiYoAiXYA/3XGbbv4NIHyQB8NdZQqGCZjagaoMjNNF3dkQoxOOPw4GYaOY1mPO8swpuFBNnid06
SfPPihMDxOYGoFtdr+e0y10/fw7fbLHPMVSFM/aaQeFNxDUF94XqQHNavbGHHfROQWC/Rrz8w3qw
doJvHRupEmVBAgvpeMkVzLpF2z46+cyVLw9NUIywYF3bJOFR8F8k82B5imOQIey4TNh2HO1drQsH
KIWaEsk2PFOOj7xgJQojdJLBF184QIIa4LpXLAVCJpRe19CCXrhF130DyObRBCqTqpVT857nUUZs
BtuvFpp5v9/AhWZd11VpviSjWTSDh6f+DYRCv8wRKZ9Gker/9NDOYrIihbTaToGCTFFJPYV7JFDk
tAz1/1zh9A5BjQVMw8qV+uoHbkPkyAwQ42qWBE7BIIb+aMCCcXa55rfn3RBREW7xnPT8WEwBssEt
H7TIVWxHNEiZD4HqBDpOV5TuQMVwR0cnZLPZoYz3t+ceXlKEVCIKP1HiXVfPDROV0WUeKxaY2fM9
/bFvYh2q4nc2MlvdCF+WDowOx3SE8+BDSU8a5oe8sExESlDyeDRjYOSZfZfF/emqzuC34gCX5Cln
9NuaedokV7s8u2vqgpyIeaKGr0ifkA4qtIP7s/Lsclsbrwif3DCakTmIWSY0kYx/xbnNtpUV63Hv
Gyd4Yf5Cl9OsmwSYPeM9mIvK6x/jnp2J1qFy5nhKIMisuscOw90R2te7vzZCQqe0uYDGOQI+6gAM
9e7f/yQOIPQFBlVhF43q57b6cc06eehJQK5l5O66SmBvnfdhYNyrYOqaLNttjGf5BshzZMh1jOIq
utg1TyYW/0vHoDwKzPTLuLtNstWlkVk6/CTzYg1rPCiW0Fz6Tt1hkaY1Ud+9TRNc7NkdTsl3t6XB
7BSv9v8AXks4yurL58ox7x9M+GVcTyrFWjkaH/IOsJCqdEanoT3N38YTmkzag0exwhMB/H3Ow+B+
nNXpSc8Tt3ZoZcFEP6Ll3cfrhUUQY8PvywuFB/MtON0nHkEZgxHWK04x9/7o5DZE18mubzY4NZBK
hZz07Y4z2IoolO0l2CTsgyLrswSnPiROw1f8kPx7an7Oqr6jZMfkL3ySZBbdjOfNZZdN/YKS8py1
NMLlgMuVh4IUBgrGk+qXsjj7EPmMvDtqsJ/HfdwdW+WdF0z9ondeMIkbkEgX2xkFjP/ldAD/NCC7
NWPRGgr3MiToySVyuDHoT8op4RwayAs8url7jvc9ZIaneJEJQAv/T33hhxgg2+DcZ3WUKne+YKuS
VH0fDB5K+6tAIr4XmT53J4VTLBo9BQ0vQwd7eG3BN3BvBxNEbrXHha7F/dTQwp1YfcHcLgS/KoW1
GBzOnsTDglkgzpKoed/ZXehGRHGZR67jFVZqIfifT4sDoQEkcotA5kPahIke68XVNdemrihflXTl
TWfeUz/rRX0OTn54a+CWhUkw9atXIgohYHVNxcsKpugryXe0agv+Gkkn1UQ8/tAREHbU5W/jHiw1
kjv4IQgGCLh7ypf76yc5ct/qRUMHDGbFIBSxVJ/Mrmrcdr7Rr7UnyiLyDgVpwr7v2OxNzhG43tM+
E0f1RzFjyaEC9kZVlkCiNJkernXMFrc+G5Tf8xcoqdFS2pB+i4ugR9FKdCG95uEMxDpAyuVAjVWx
G5Z1MoelDYvU+n5G4FOjFHmmK9aoMN3VUfZsB2u30wu9JWHkmuQBEWLhcre/xuDQPtFpoeTdvxUa
bMVW1WpTcihUc1CwpW7TjI7cY+UMYVUftr8WK2RrLZVy0N7rmSRhN5JdTxEx1XmGAm2UHYJYqlGG
FusaMhnYwotIc6/YuxvOysNhsuyU+J87yovOyNqn5r8WwRsCqnnIuzD6zQGYP1xoIu5Cy321ax//
nyoUpsNm37RH82dzbeqnJmOcQp4omWzU+BM/9B5pDFsYKDVmShIQIwMKCEAicnpY1BBz35Hs3mr3
+cBOuUgGd8kZfWQn94Tp+0Qb+bNYl0P3IZwzrS1+Id8PFg3d2ET3h/2udobsGcnT8kPa55PoE1Ym
76I1piEYRRUr6xvBxl9BhuVgUN4s/iYFZxh4vH/+Yy3HiUaEVCfitk0ntyaTxOUXlrCPpUIvSEGr
ynRzZ1Ui7UWOMkeXxDXVdl4SGLH0ZEDMR/nNDR4q2yLm4wutnx4dJl1sS1dyaqolkGEyGynZejwv
bqCBgTiFt+OK6cWlqoTk4Sdqw4qsg+gh7i3KxgE8rqmngkbaoLPbqTlCP2wPxsg4KmKIKjezmMPM
0tAypc/Nm+XC3LG8HpA73vONdosaSut6MP7cxzcPcscOAIcicETFJpb8J/c9aJKTE3i96tYKLsjt
eFvqhxNBV3zOtRWWbwUiUeftLbIBQhpAMrguIw17W7u1xNaOaiTaalfsCHoNTer55sEt2w5ZKx7r
VzlvF7FeRB9x9021JeevaRjkVmKtGsMUQxil+JrU7GW1orfEIPYqU0ru1vlrOfix0eS/e44z04Bh
lflzJdIoOD5EqVugsukgzaQlFrDfE622xHsor3Xrx7HkkdeKz+sg/3qiYyAHIjE7C5gOIawv5nVy
ryqPcy2jqDFejFnuTR9cUI8AxbBbbZtwnD/NBrV/D7yjMc2UJ5XUJnzRF74YUJstqdZtOfjSEyrU
+PNrwg9IR1bxeUTxe7PYgT1y/hi8qmzhmWhEbc6K1iZ6HQsvRwpJrw2ny9RyA6ZEIFROAEA66Xek
QNdNkfbzE3CPyGjWYfIHqdWa4OI2QaYXt4XpiXKfsLyxo0G0cAYT9HxSndfKv2BFe04mh6yEqKl8
ohTKAcJH7fzRM1Qs9+e/ecTOyXmO+SuO758fgFclCl291ECgA5pKZ5PYGG1d3EkvDf7hUgLAG0O+
bgrXDUfCn+R+5yQlyPPxyiwEn0giTjlN9m8hDytU0m++MW5eI6m4KaLUkuyTPPhzz2mqOUMDb1ke
zj1PTHAz2NPi1azXGi4GOW6HELicieFYNwKrIyI8YC/P3BoBQ2A0c4qqOyt8MXsIhDqhjW0XfRvy
XMDWmK0JnaL8V3mPO4HoVKLfdsZaxtlYy0XX8ReUGYLE5Z6ARnlbObNGtA4SixAgyRTK+fbcq2z8
2liQK4lTzKF9Jz/K1qeNGoKsyhk6M7aAqqxm10cVBzcbHRMTD7iooDAZOa0pvM3tx2188xoDVL8b
2h5LYci5weelzHKUBs7CrD6N9XjRZPiewbVbF9uDAbkMdxbbZof0qEqwvcG1iriNdzmPOCqpBl7d
SKx/t+K6vmnuD6As3DLfSPSVRH6SvRssjWZ79B6S9f5HxlKwnBr9CFVXWSQMe8rNYwDO2Mp5vu0g
szFA0fKlw1ImtrACdOTNNp8q5AnDNuoWKJksEYMEWoaq3R3p8yug55E0R+mcB+LwRDFwBVDjneqx
1rpeL9iYI4nG5ZqWYS07w2GQSQSAe1nm1z5s1cO7M1uykr9iye1gCbipjjf8Y3Y1cZUN7A9s/FM0
pKLP18kvZgBywu6QOQ0zAFLDeY4I0o5vnnltX2Etppnl3iGGhFqBm+RLvDPQRIjsJNY1Uz/ICyPl
Xm35WMY4Ew0krCB3VIbu3d123oOnKOML06Lu6kL9l0IM880/pWRbf/x8Pz/sJRDAa+geUfytkBTd
vWfhDoZgN/POgkhPQc9Q4LtNojLc0DzVwQHiF+4t7rwZ4Qf/Zrt5hlxCahPUagAF7u/oh4IrE71a
wBGafOkRcyp5m869OFLAHYVbFGAx5MHA/m8u/SzMx0fnBoi1mCDiUjnt/G7+ygWAyzRZLUcZbVJP
dzuwY+1yO+sDMrqsbpb+vJrnoY0wTDBs3tPY2nR70aFabULaUgc1B+sDz8qvcD5GejMqFYHgV0V0
qJVnr5qBAEl8GoRtfiExuUmkA+DilzLnqNTakTSih8JQuWALsd+o4Ed5oJpG8hQP5vZCtSGoc+jo
EcHvO0itb9AjAZlvK8PhCu2II9GtXGql+9YpdyP2Vjh5mIEJbfvhYwYa9grEVVlSLxuDDhBGQQhj
22oGrdIH4nafHFUFx52/MeNZVSuY4Za3NVhzjvZfHz3JaBDxLpedKPajt+UPhTC+aA+cO9+Gf2z+
5L888bcaIs/J8ckkv2vaIwJVyHxY+ZJaw6g6yRBtHotBbINMEn8/FmH8M2ssDfwTDLx1XgupZgCJ
k4yCDtgtRcG1Z59E1DY1YG6cJToJoL7i1q1I7sJwtBFKE8ADBPT20KFd6yBIBz1h7EqoM8I4Ctgl
rVFmiAOF19L6kf8VjC7DoGINgOdrFd/tvmK9Ze//0X3tSj8IxuHGgytJ87JrprRhcr+O978ebt4I
02/VLXfCocJFmaVDu7yHYT1gR04ymmTgL37WybcAwaZNQkdylAqV2Lv1Wu0yOxGuEt/662EReo/w
eEXFX0jQLtsAsAgBPO0bnLmhfuxfZQbUASpK0+86CUYP3JwKkKju958yk3KqRCB2AzdCr8LFThiR
p9/q5XwKeNX+fH1MuunvtKW4XaXeciZSxmqTYNCH0T7I7MY1Dzv28Hdo8ZKAglzpNQyFctJEG2rh
q2VBD1W4Flk7koFnjS/viEGxxJ7EBGbu+SyE5OyMuS/dLzS4zwP1y27vsUXqwibNqbpH1OO4vwga
sjxIsy6m7uoQp8BOlP13Xqc1QgLrjKIBmGhsM4gso6gTZq+EfZ0q74CgaN5Tex9chkwGDwVYS9N3
4EXFox+yW5EtJzFoTtfDLLAG3bDk72///OWxwWhBQQykGkkFEX9b/6yWqyzjN8BEo7xuoxyAeiIE
gfh7U1GV4PMr5Fl9LdgXBpZOf8Snqu4dFDGzsFWif/XxZcbyYYrvI0tsFUy7mMWKri8yyUZCBMbI
svTkRTDBxP33DazCv+ybernSbTbEgkrYWTOhmyhiTkQdZiX8cTLlqYoKCCKB4CLfhU3KGMNKK1cR
/y3bIt5ncNrkThInP9p69PlPx7/vyzVvhd0jWHnJ3zmnTPCdnJaknf/TW0OKcNSBujzSN+FN83eD
ftp6VkzfnV3aHMqTRLfVXFSKIEo5WCADhX/6k4FmPKzN7JVFjXRqiIEH4hRgM8o3Cj1XfQSJ3JXg
//OnzXB8WCreiQ7ggIeUWh+3qY7UUoPJ/mpJyRGX3huHjaAU9eX9ks3SW/CqpYDxE5LhhqaiKA+D
Ui3UJl7fMXF2Ki2qblnqODrsifIsEqNj8rjVZAY8AP0ZKAqSE1UK3+QPDpiFp5yi2/GPEIbWXGGe
OfAIC4MUKESqneNSjajVonYqgKBYeyteGFbVcDNm7A/rg8qkviurr/oTcCHNQxf2ekc1G0ZQpVy8
Kf2b4xeemKQcDym1VmfIZ3axVkExM3NAi5JXpYoPCTJMxUSsqbhspAGWd9pmseKTT1VURDllaJCq
W4HLupn0YUbZwthgnITuSOoSc9+WAlYDonXzz/kmScb95+jzOLkRtcJKXPGtI4v+Y+Jtlti5YlHl
OoRh0WnTczxL9JrMJdxU63YZBho7DtgieWKcRIb7aaRuDyPSDuQXIPQQDe3/sBkzuHlLKzH5o6mC
OD3fieuA4nhUiQmWlSYvfQHcQDMUJZYYYkoFJUDjU07t4uxMawuWk+oCKcY3zNVotRxSORQwSSeX
gG58Vy7uGphgrYmd3ncwGYIki6vEvJ0eBCyndbFCuoXAyIxYMv0kZz2O1INQzdVE8iT+Im1y2Zxp
rR24Iwa2HCHs+qlWpRYIXoSHYtSKwrd+NYQBJctmKS6Qs7XPYsUJdrrDcPGlF5NZIQSw3wbN/DDL
u4G8VFZDU0FCcVaKhloQ/aUgWppUS50U3pm4xSO1re0PcArkLxfMsh8i8MsfX9B3+FkwJ9sLuJwP
A3C8ojnNICB8SPl2BJ1TdeyQf5WrXzhtwmb90sGc06sGf2+wdqL7VVtuWpKRqLrxswJjEfXxWG7A
lX4pUELaFmoMx7n96nHdrsYP+HxmowpH8ZnTedevboZksnJJJp9fkQZhLzKPBxF+6u8embCVBfVj
P1FYYavVPZ0NqEmPXgli5KAxTWNDIjKLo6po4kYCC+aexdRVLm1CEe83YuP/3UIpigiXnaeHTD+3
iXrdMHbu5bEs3MfLI8LDDfFly8Qbra1/TkjqzRUN0/JHp/rqdTQpIB6Qtt0Xt22D95p1fwpXdUgO
ZBttPiFQgXM25vqq4TREkpkhM46lH0WZoWzxOlfH0KvLeAlwETfr0B79/OXl1GJGauoKrA3xd0mu
dCn/zoMM5LIGBBR9QrGn3u+y3zGJkWgZKjXg/IYwbnYamo3L0GDk2oPH21H28u6EClNE9oD20IPP
qyKii70WS4DDtd91gcEeZFoiXEijZDjtl/dMMtCgs2busQsmFYrfyFwJnmLmlGwMc3SQ8vFyUVKF
rzWIJwrJT2ZjoYaqJtuQgHkm7ZS8mA2T3lm/2LLpdHgq7PtbGOXCpfb3loz/54lIa8VWWMO1v4Yx
GuZ7XCPfNtmuxjVHb9mtXFOxyI8fBpZe4q/LCe+gkB6EciamdAIu0+J/foZwutJdFXRTNRPb2R+W
4+zwUgMTMMqSCnNW2iJ7ptZWwHAt0KpEZngVUV/KbHd/GzcE8FXHwn058NAtWuVXB/OPkyaFKPXl
XxwaKFyYvhuCvJB9ZmK25i/LU2KXU+uHkNGCvC0PDVCjiRrQOBGejF8k2R/UjHQkrtLP6AuE+0AE
GrgR1LC4dvIQjC2nE8ibmki1nojV0/p3iH8KnAMVus5QirehGQ2TZSNLVdoqn+FifCyCsE7lnrKL
D/TE7FecXCSIbqL+7Sw+HuHAXiibQfyH8ZerGgJTxalAkztC8QljeT/2H/FXYD0SZAL1F/e/xnah
/mmIlkhCONwkn32SQWYOqNLwhpk9J2j279/cXi07xOlydUm2V5pmeX2WW3qmGyzuG0rxECBBMmwI
XhOmkZFgz5HijaYH9Azp93OdN3sFvSE8kPi78Lq7pFqwPCQLTwDpJrMJ+4LLHgD1mvRG3PIuV4fS
9Hnil8N54pCi4MyYxka52x6vde0yZfxVYpOxBsjK02n+3JMmDA6vAxIqihFJAOD7QkfbLFGTEuIM
EOpZQCNsTfAF4KgXmt/uzhjKhSfZC6PTSyr0yMNPsz/1phVRCLQMV4yv+WtJYs468/fjOmYJawxF
ZpYO+aaKMeH0BDkihnGaEajVJdvUPNl6MfG6JBc/rMsPTmRNcDSLOZHiZ3J+fz7qp6J+o1APEipB
sZjYBSBba2ZPkOPQedg8eVNmEre+JIqT9NwcIC39WvvWYB4WSunPytjfHtImPbqFIleOsdd/zQYn
Le/7j6I1UY927rKbgyVhcgakmfOxY/NdrKcA5k4hMvQJSkj2bACLW8HxGNAc7MigAJOnyztxuanW
TB/Ceq7C0qH9Yn63gIrlZrjfmCTWgP1THwR/7THxm5rCGDzJ5E+akJOTI/57Lxn5V51I4oMGPMYF
0P0GBhRy2cAhaUcCB8DP2z3aoxOpxx9bXbwa+Aw2rAtm6Cx9bRhx7D9LjlGS4rpFWXCCsutlh8Hw
oWWzliUd0x2Oza0xC7eH5GuLBIGaEndpKwbGdzsZNapHotofpaMhMl7hQSCQarUoYG6BSdtT3O2e
tzz+u6BIpo8RL2Kgl7cflJcDrNPzL+6a6YQNcGeW+F9L/iKMI9VGLUtA6hmanxqLJD3TBhRgjBPm
1uzQArInCd2T3znZRlwoULkAfyPV2/qX6i5rRzhcqNBiaoVpoLaFFmYxB4DM2GYhlFp+T+p8pzfn
GSO1SY4vMDDlTmLLZNbXy4FeU5jpKQd+x0eTgvqr1DkchhYnomm41l+XFmy+RtDFmKWMDJsmuojU
3QaurYA2/cLqQbutVLfIIbfpCNRGDv0LDKmt6TVOCtJARTeo9qB/D4UACoqMElHdzJxWpSawHnBd
bwqRf8wJHDSgfK1VhRnoz6C2zxx8RX5RlLfkyqJRRLRdxuWOuD9/BFFFuliH3ZqECAKVWg2FjAkU
FGY0d/qpPcBF5g+ic2swISHyQCysR0ljIJaa4Ht6GoQKy8pRwjO3Pbv9/yRyBAorZrWWv5UpUKF6
eJ/QmerxLwQrc3881kj29xkDervpYfXjro9YyOs68poGVlCibeCxOfrW86UyOz88kd2zYGJvEOtV
DzkGqoqA9dmJhq5L5/qlcMRorXb/Hu9uvBVqVmkdDCClq8iboj8+qX2WXPfZI8YhhifPCdFdRWl4
OS4i7WvYOCV4NoSrWvXLPB9yFfJ94oB4jcjyhRWoyUK8gSuwjOALz6yUZHg+48+K5kfXkv2kjApR
R6nhsTBX4ulAUfgkFfB/BNPCekf9rJYcCRw8EKp56uX1fzcl/9R0wmJpXhvavoLjusKSU9+00cFv
WBFgJ6KByNZJdCpKN3NOTyYAuKZpNvQMNN1gqbykv3Ex7uR926A2KIbPG3OIjTHD3Xk76NcXzRGz
1UjGkjBAbjQE3DKpF1N8nYT6XtypiG83NZf1YFormufjXP9hDKjJwOJI4ZL2gqc01bhlTVXSXYRg
gHYm5eCbr25hM/PHC9rVd0h4hjlW4DxFS2oZVZPWWdFGo9PHGOfJ/QB3XTybOK9wcC52rB88xC/y
UovIAqmeT8Lh4YbddCXDVeXTAOYeVKcQVo3QfUFzKlmD5ngYuZWYoXO63qUGJ15bquyqPZu7159Q
OIeOQA4ztikeCFcpB94hyiZJbOaf/BXZV6VZjMopmF+mF9Omd70gp/BHlRq7h7yBN8+cVwXRklt8
xL9s5MvyF8IKRPLXvFMEE4kpdZSW1LL/5PFds7dBbQ7HxoqhmtkdavYU2zX86/8gSX0sCEztM0A6
DzWm660TdGcxFZC0ZW30u4EnXFrrNbK1Uu8vyCu561XtQc8UB5ublmAeEx/B2OQMtNkA3tFhVkXI
B4NxAQ+XKub483VmCjf5tMyD5mwGurRTOaTCfLa/fWUFQEf7SPdYVT7mir9rD7rN5jzNuItQkKQN
hbmwPrXcRQDff+qoL4tsQOtjVSWG4n3mop8Fe0/h+xilw5cDycFww6o40VLv+JoyeYmwx3NKQcik
pRJK64/hcXeqAqDF1jm/+4MGiv74fFInezNdPSnbMd8RPWDmBIHZy5yYUTDb1nxXoPcc1h8ZWsjB
ct6d2rd6W39NheCHSkY+GUJXLsx9tRJieB8wju+QBDTMJwDURfQB2sqXN7t+fe/0+blAjtDBrtBS
5OqST3V6PN+RQg238pblTPf0jmfuxUcydp+b7jwCMAl7mER2KsHWOWiNxrpKBIRvgIzMixtQQCJX
bXSjZvN5GyGX+EmVsSod9v1tdBsmywOssDUsoBwl+qzlLkwlhSuCHmzgBG7ZWm5NGl9YYEKLlvd2
KY09OeGSCQ8fsFv6t56JKy78WYU8+qwedRhImRIU72vK6wPIh+KBz7uPlqUny8DIypjbfZYQcJgA
yfgUFvz+dHFqrYlhMDyH2d+Zk5oBCgBanef/SwNmatZEQ2Dt6yyJB0W45ZPTLRJDBfmWUEU2JvXG
pFLrXXyTLPr61MLpRZfOibsFZ48YL4S8cGAAN2SYO113FkwfLDoRUM8UGJgB2IWzZldP9XOZOjwI
7v6LugTcFxOekThpzaaQDXk4nCheZH0Qy7XkA8FhgETAhZV8w018tbPOuy6MWEmJPV7rB4q662br
UtL7/S/4+Jo/CUrlVLkJ5hoA2ma9BQOhEl4VgtcRy7PLq8yBuvlFrVPD+4DkP+uy/kSSZrZY3OWb
XwKyNYcT1oe7LZaIhhZ40Tbj0raTDHV8zme1mN1h2RHueAYiwv1Z3Bph7VelTfmyJsJvJkHPOLtH
X20O9P+kEKxDGS2VyZjQv4Bp2xg+967Ue3CCZlJEPbsraShOJE7tDVQsnr6suGk2wajgBTCQTGzX
UYS0p4Em7+IcWvKxvUd0YbtaFnk08eB4eVA8TCETfu5BOP2z9szxbTF3tTWSSbpp/DZ2vj8O5+nD
uUP6zONKnC+VrW47+N6sKGnR1nP6ajbh8PF8PE9bGweUJfkeZz+8kNuWq/0zsduXtdu5ov3uwUD2
U+3lC95veqI58QzFoBnPVCCjTh5jyj5YDjQhtCb7l4CnAE77/4fKgd8G71I0qzbTXaVYnn6Sf4IB
EjRWMAKnUuHtiP+4uAHNCXMrCkTGUPwcerG/BTHmkPuwUositip1VtlVCdNGqxnVKWYt+dOCtczU
6qVgoOKDTuP+13Yrcv+nk6RvNHaBeNESd1cr5bLU1mtAVI4kYMFXml4pF2EVTtbDhGmuVmVdnoZt
DyIcCUySNA7bJ2HfBNvpQk/g8nIjzn16RBku+E5xFlXHMUZKdx8s1tji2sxco4cNBM0i+yXjNK+z
g+dIxMoYU9VQ4o5a9GNNOJ/xFLkhVW+M2/O9I4FsTg4IOutAhRyErQ49SVuAONikoA3tvfzc1mdS
K7WWxstUlyK/SuJISiywaeOzRSvsRQpSTknMx+xToRqzx9U29fdoNj+5X8ZHPMUy+OC32AV6xM4H
YwSaQo3xnqSuj/E1c+CeLk9P1QOz7QyuwZI+NCrbvWiaLKNPPLcmADWwln2Wc0+jcgt1ekfwaEcj
7dh7HkOxgXcwQbJgYzR+7vUm2sqwlZnYc1dssp3fA9IAMFh4pia8tZUoJOWwAMCN52CWUcUs/aci
BEOVc9UYUeD1uyeMvq6DRlOo4HtZcA6zHd/qH5yTGVxlVKBhfER/6nWqjDeclnVOIHiXoZHB+7DB
VSdq5I0zRAY3pf6z3IM3Bs5XKkPczU5wUGRUEWFr+O1qSBNAQWke7kx2darEdaTD0PoTFOWlPkiw
FtyUDLSkRQLQHxEYVrIVdWBL7V2OVFgY/AWdNJJK8ytNDJ8+W6RbPtndvXoV7Vwp4H+208XjfvLf
6bLRhwFzxDwWbxn4K+NJ678aZWPIOkopydPeVGZqEjBOPZXKjbI2BGQtbhFzfGGCpgEwDKuA2Ly+
6Hv6RIIstB5l4xzvWLZcy9uL6w2+Im4vnRo7zXAokreEMTM75Zwu2ccc0GfhzkQ1VGgGWR//p9pE
18Deb7qEe0KXFqIvL6aRLMxc+FGUaSz2CuA1u1IxyccZuDCGuHpJtomnyu6JgedKt+lz4qitWjUX
IXORTSnHq+rQ2IWLXOoOqrYlzLvOQmi73u218Z07y/0rewmjnrvHDsHuX628pHs4ttbMlImoAONF
LQxJJa/Ciwr9t/po0LFmYnPu3YZaTHZgKLm45G+NvX1xlUEfuYtLlCg6wOWgXwQ8et2X8qrKtgOR
+u9CnxcG0JfWQkMzKQ4QDNdHyQl//DRmMX0ektMs8hZiuA/jWaGOnSxAsG7H+9HZcSo8HkPvJ+WW
0c6v5G5pNdBQo0aocvtwOnAv/QT7jocl3BgoSQ6OdpPK0HZqVYL+JOHBETe9HPFe0bQxKuLF09/J
v9GvTAZDNCs0KX6e/QH7byAAoMcjU3TUKt0/+sMW4+2h/fNMGvYeJJKZlH84zDRqmfT59Xrjdj88
IhIJbtYs4cZUTy7zVWN4o8HtiIwj5PD4SNf67oEIyfkTfWyncF1nQI7mRfDeSc6HQNgKyGZes/tc
AQHyB2oRbmsOTk+S/Vk+49xtRySooN4swKL1HarjpQQ4EJ7k+v/hRE0HN85jurGhWCt0fGxVNYiV
v3WSHBpic9BUXBwUn9C45Pyb2lbeHODJGoslDiUME68bVWhOEI7KO0uNz4LGK4M5dZrPzzYSMlWe
/e5gKMR+sy77KBneDNTu7WLxlmpkI9/GaofGK1+HOP8bQrRllPewbEsMbRoIrf4emqjxMLZbwO0F
gz/jD8WIt+oiAXfeHWv1/q2jafmD+dvOtJaLe62GGptfyghtbuPuOwJ5uLak9pF7muQBdIT2zBDg
n7pMdjHu9y9cwtKgvKJhjgHMp/gbe3qXVxOfVHhFhPrUqCO8J9OhurT5dRwK+18cs+oe9vsJmuU0
xcw6B3igzVoj6m+SXWUwJ8/sBYcassDpbfMFvWYkhMreFJ9sU/oJkpZLzVFBghwc5r0K2QTJPgfy
+7dysA8mSC/MRghAmnXk6GETWV9fKHsGdaQdzVcczjgeEqUmO9HWB3570iAki+UpRplRWJE2vm+N
ojXYj/GNgJgkEVh0j7gJ4MYNSf0XT9U+1LCTJTEVqrMwKSXX82V4TQL3zI8bVxyxwRzmheb/StIx
QBB9/shWhLRnsz9k344MrkzxsblWc5AEe43RBwMpWr1N4FGCUyZhBBfpoe+mbG960Dlo144T8uX5
u2YJu7B+MqlPk6PFBtLzPYuf6t3fSkgZ/BGdcIrJ+plG+Pj3InJUoss1zqbC4pgotJdWfDFmZDYC
PL2zxH1jIHi0QsDc69ncNlF/VPEYPclsGsShjUPcShWjrMX/Rucvij/MvBcPn7S+E13PXOM66LVT
eXy3XceZG078Usu1rDy0fca8DWibCWkAejLCPi3Z+N8QxP37I+fOo5jk3+0GVqVRrkU+prSEH4ip
qOO09iXooth6KLuXDfiQiMhC2SgsszEs7hIVaSA0/HykvLmb1H/4+l0zhr3SnUjqShtx2CTKDR+2
3zxiuUlRBzd8YtQ+F4fOefINwGPVf+EUbzvUcihPMv5Es+8VDz0WAXesAaMolKccDW5ZroFLcbQT
Dwd35aF3aejEh43ASHPFA56KH+ZyhiqsuW/FXFzE+rdhsEoRARgbGMNFVuVBkQShXC9WdsQI4Pdy
AogRnekZUpy9dYM15RKEJVMNnp0+QNuTPXMELZZ10fArdBIal5ABthspODrDodAqN6zqPrW9t8yK
l2I3PJOUUzty0CF1xkrtfR9Bc0klpGJrq66/i5M5O/tZkQyhuIiS+4gIWwb73MhsfSL0NsDZ/e1l
4JSO/Os+WHcKbVzMIXPCD/wW42OyHlOsRGq2rrMUyQOxpldeeXPb06Bw4Rf/2D/BzL7vKW4tMn5b
FpkSEnbVkapjpdG78sHmoZao+vB81ijFFOlIRAVszO/jzkN/jdio7w0r6fyxElkqzHTTssbOp7As
FUmrWhU959YKlRmykfB7o1Eruun8gVZSt26yWxF8pgRrXNz/RzFItl/MXqTLrc+kAaEpFPScfPJD
rS872J8thatBrxVAaB1hryTacgsVmmAU6qubsZshhJRgqoVVHJOlu4T7tBkOEHuERACsdeBbLJZE
pKZArY/cRZ9mmWAX/FKxTfKw9iyF8JwyEtTSDjpT/QJK9Q7TR0L+SXtXFU1dT0yif57nq7Q8c+02
nIWyOI1MIdlJe6hMqQRaFN7iV/Wi+BhuRVEoGSC+OlKOoexZxGYQT9aDIH4WttNfv83aaqOWaECM
5N6iZx18wnaiVPpy0MKWsx1UaXq+EJAsKyD2g1cCfoyLxW4899QaOW0Pc4hnL8pfpRTBiyJJc6JE
mVgOYnAG+wpb8Mw9E52zgZ/RrPRbxrSAuqMH6S2MWAackI7FQ0ROpwKO3dfa4Is3Bka9y7ZYhJx9
a3PejauSC0vxIi+8YmrefmdUzl2lDq2OqSN20kkKVbAt+Vpi41oydWfXG+Z3kbid4+UDty0Ajv3i
3mPZ/9qohPRRQ5SIkUUA/HkEej01OMI7t974pQFfN2gKHwF2P8Ac5aTc4kQq51VuLmJNpTxB4DCr
WS9JaokFgfRmLIAsN1NT4MgyRA2IFvi5XCxIUBjVT7usdC5Oo5tUQQvs20NKK8+F4843G1wUR6N6
0VrtyzIFbrXCDhNhx4OEdoukxT6ZDk1thSyFGXsOCwLx14zA/0/vBo+WHBSlMQP75IxWoX+onKXJ
nFyBAS4q0eTRbgkCvPAb/sSAHrM0kwcyZXlUJRfn5S3Cw+UjoBLPAknG/Ze8Xpyhk5WxpuriOSwP
vAE6KKL8li2fGCLklR2tN6UxZoBrflmiYJkfPc6S+SIJkVFi+JXfpg7NBXk85idmjAvH/ToRR99/
iXyT32ebxCJXsaqgdHPsRdFk7zkNezxpSfKctuoUMOu4Vfg5qsV3QVJU/PH8wvyxv0dBpk21w0iU
JTO8VJnvie4DVwG5qFZjfTRIu1X5ImeOFYv1KMhOgTfJhLAEJiXIGpzbm+VfpoITvKwCrs2wZDAS
L3rJthfodXO5CvYGvpNrAFJW58V3bB1TDaEOWammxiZgGJuR7QIAp0+QauxeMzvFqURH6/R5mxRc
bKnZzCS3n/rrW8BY+JnGenl0cLr2xEwfu8mIPcjeC24OKsUuprN5KhP8VIZ1ezU/qniL6zH+amm6
Y1SZXmMzs3iJV3XCL9HGAICPt8n0rS9YhxcFQnNTHw12bKOC+O3YyyaMwgplU3YOxyTBrn68Su6d
t6gwvHh2Z3O+watW56d0owDFghrQq/7fS2hfX48hJODDX+KiOWDrTn059JYGjivtdCoiPF5HTvgw
zFp1sTr+UQCX/+8/ru6nizbH5nF8pu8OT27nNK+AgeOoKxnPswpXb2/EILGWNo8dJOlrJBV2w8/L
M6NA4GtwgVPyppPlrbdC5vYcm1rGK+FfPFCzr+XQ+OxCdZH44dJJMwnYSPp7Dmuj07qakYn1kPPi
ayEuU3KUKvDgCUaSL+DUFfXojkA/ygJuQmmfMF7aYCZQrBgiGY5QMesk/QunurQT5Q/9Aj0FqI1f
/Ph2nxLXpuggXvmVgTbFGmkcfO2swpkTMvgE36xw5x+2F/6gaq8TFKLpDd4bjV4gIcyBDzgb02+k
aRNjBgi42kuT3NRok2sLjYpuiKEz2IgH5lgNmaiiHAI3Vhb2KIq3ze4iRH24UZSUGSCoRIB8bGPs
qX5POhL/1uz0SuD8SKLwzS6oGzF8dvZc9HKfVo8NxZhWDEdmppzrnQmm3SaiRJUPIQsL9B+z0TEk
dYoOFgfmT0QIYuP0XeV+liJxLq4axfOWS5kqKcJXqmToswBcSn4DdHIyTdLC2FAm7mImJCEe8nW4
S7nCb0K4desH8ft+or6YAJvupiJkrsSXyT6GggBiPSNRa9MQ0kj0zzL+P3oUNk38IOGvrpznBjtk
JVuuEXocNn/ooIq7lk+zrhqHkzeCJSYGzjbqUau9RLF8C/WFIL2dRVn1p5CT5f2KH/mIZvcFt96W
IwGM+6/+wAgE7ty8MdGhquiW5VfWh7RJJc/80085ev6kk26Yd1W0yp2EKiPO8HXwPS0848EdP/ia
w73ony04KZN/xOX7NeLcEmchzQeTf49u9TOF5o2Cp1PZjwyPSgy8v01IX3r3qiKbUjHmeO6O4fcJ
+lpVJgmAqcOB+0x9WHifX7iOhCsVQvWqwS6BF+o14aNENlvg4iB3EEJmvcuErYkPmxdxYAh3FrAX
/nPlpcTTNkTXJtuAv9cCQJcRv7wMjQy/Uuxgz3wP4WOs+SqMMRRLfV6iHf8YjwxOh4FZR3yzhBZv
2/Hc8sXTOSvOuoU5IIuJO7KzbDcTdfr66G2BN+6Q4TnsDB341EZdoxgQccNsaYqAGd++m7Q1XF0a
NyyzykM3JY640kw97Di8/EP5fuPn1q/AmlYqezt4vtCzyUlThwYXbY7acEta6kxDRDAUXGeQRN2K
Z1LgOWr1nqeiu1Wx5Nx+fftE4vq2AqwurEbB8BagnUR9GT0HVpQIIRSySCyQC0zei9LYgshiNex3
afv2dwJ0JkqkYw8CXHMQhCtfci9pN77gpJ3YTbltqqman4K47Npa4w1CL3yeAWHxoMUJROnGiYSs
w1DOu+A8JvjGOYp0skdz+SKNPcikFA31gL9kw7DLLn7GwhLQahZs7sq5KehTk1ZsMqBhvGWfOKN6
3+mbPay8ig1C6Cy4XJ/Ed6Q67rH060qSTF6pdBQrtkfyLwNk1dKsG1ZQWdTqBAqbZd3HZ6448RR7
aaJwCl4IVHPL8tXnm5mEZkqim4+oqiJtxaJ+/uNSN+791QIfiT5EqSCUEOCGJvKzKP1hJKIxFW7u
cX73VREs0lHnMlY+fwS6s2g3d29XY/sLTKMEQl3z6Ywg1CuiG5zVPQ797M3fgGazS3i/Ng42tvuQ
WjoKPjo6uKaZYYmf9oPoX09NnW5hC+SgEaxbS3SqB9wcdJsBYgDnWJvJyqJm6Rg45v5m+0kdgcF5
s7liQxOxhaCzXu1qfxWd8lyRVGwkT9hrix3qV38zSelmPKwQ7CJcHvwK5M/EHMI4Az39xVA1CXn+
yXBpcHR7Jwj3NQvsEGHwZqbmd2W3Y+s1ZFMBhQSEfDXMfvhBzi2AX3u/d21jLd2CQfsP5bOhnIWd
wzNvNYGxpeHfbzKF1SCdbZ5SXPl6PI92DHFSVhy1vGU6o5KvoqifswEFAbehBlCOdwbqxPkLgh/v
qckkX8Ii6gS/NrNj7O7x8YFFOE1ZRCVXgpiwQyQXml8GZfVgI/sa1YC/HhwMQFQXp4yHF97ZefUA
gn76avxKL2oEY0wOmXPFsA6yAvvSE44CDBYL9j+VljALrfVvyU/3R1m3f5V75Y+zb6seYWvUodnI
uMfCRpZAYFI+gQZ+1wcM7V5ucrcVYXPmZGZFatJJ7uWMhMvSuUS5loB2rH18N4aSoo5znbgCOpvE
H9me6a90z3TqPI7/iZbY2v5iITfLTWXoyL1cJrLv6nmw4DtKA7ngIYLfKN0MrOy+a0LH+x96TEFf
Ns7kHSh4OMoUeIMYR/RqHHOMq5c6qGERnzwBFpCOo6BgefrWTunMxHldNFlUNoHFFicObZmGHdn8
mnVcgLDuwJXNdHOtvOXTR3S5/ZLQBbW2EEf49tNGn9KBXoRS458VDhXn/4/HMA1wBR3otu60jsI5
09OezWlK3H6/JD7RDYCONNugIIZx/kpRtH9MBW/XB3dZyRYTT695LUG4AnutmSaDdXH6/qNfKlbj
27JX/4hnphc9fMoOiEX03cK6d72Y8K45dEMAgaOcMO+YWJe+qP/3df0KxmfVkyTMyjDblwe/WnyK
0LG0yzFDPeki8XqudfsD0LY37V77yXPauS8S2GE/kIi2/YinSCEPihfEDxGxLPluhADXrZs3iuQJ
P6/NcNfAPKrlfSQ/p702b3KVECXIKzBsM205xdi7hZxcSrnoja/YejICFjoBRWh70D2YcAq9d/jr
OgFFLfRkeJoHbCGRE9dPwcZPUqxXlGs0WjefeqImNywNlZfLiAAmcvJjGgMi4QjNo+XUKqjbup5P
NRQvRAKH+NWwvCQptw3OMF5qaiYSC83F0JAXbmDEACGOOuEFownm+YhOz2fFK/Zprx3B4Xb+9u9W
gKpIissCXgmCpengjDVf77x6+/1XwbUb/kflmXOXZXIE8PHRAcGcsTE1iq8uVN72NhuRDEQ2KtMa
riG2QbFOd1Ag8xVQFyq1Slh3QLZ3zDv+SDVfTOaPNKAG7fio+TCy8XpGchLtllslk4kBKWQh+RBY
uq3BA5G/JC9eiqbEQtstHLzTfqkkapy4dRK3N2lQaAefwqZsu3oe6G774vufIxnpfc4AhYgmenBg
8emXnobxQTbTH5m5dTp1bwhyhN8YFgnlE/RMj975kt5lkJfN0zhQK7+AXsdD121POmNhPqfjcDBm
Rs8JSBqKGUrmTMRYoTbzM4G6QuW6fMFpmOkrNudXKCoN7kPk8eXs+C6QCe95ACJ9mH3KB4Qw6e0b
XMx9CtAeyWVzf662CaqPFnqiZ2WXxCQefvrkx39ceR7xGWuAH5Tz1M3wiIDhlYP2cCM551rjzWEN
wa81i0u+icN/4Cf0cxeRnvIEMfyRjQ8dRviUjgDDidXY3u172VK4PEtufNIeU5WwglR666xxt/ie
9S3lKHXAvn8KlpE1UE8iNy0Qnaggq6gDNW3oh5EHomrgBMIM4L9+y4YxHje9yjfy7Kr6TmV1dNiM
fNT01k2Zkiiv5MNLU/xUkGI+4R/ze076U+Xdb69kAoByw41SSml1qQeVH8a1BJ/4kF0zS8NI4zYc
Qk7gv62aWc1Nz+Hn0bdDSoFenrLfn5FwkGCw3DbhAO54m33CAoR1xVeMwLMVH0pd3sxOjAbn/0X8
wEV5sSwpM0CqR5lRixlQ7qbBMeksZR8vBL9UvCJ2trWD5wu77rJwXFwhSBImZ4DfoqR7+y/k1cpZ
2MZ3n7aoXVu9J5wt2G7x0uPShbyyZ2JNeteW7+jVPCNGNDTQzasCNwG1eymspPLE6BdOfQgs2BWb
clp9wgZY8Rc2ZP3rAh1bR6Q5c6OW//NsLMzH9d3GQPhvZ8OY+5MOtQNNluOast11P1cPAaOO2Mvt
2Kd5AisVJS7NvW1CYdftGkmvN45bQT2i+rG3XNU5iwOjVu8NbGxGMl+rUJe8QiqMtqxtJWICRYnm
m8n9qHRa/l4Vmv0/jeuayd1IimZlV+BGODg6xAE4VgDaisAK8Ygu5YzKUer7nuByrmqDS+Y1o0ft
+4p9b1MDzzN4w4rx3ZO4YFUUFlOTT9ICSnpliUUsl5kqJD5FsbJS3RBdedcy7VRRejfrTE784RPR
oX1FzIHXcxYkuO/XVHC3yMNb4tOr8bfXP2SXJA5Y6yJ2KVTadjTHFv2ywSG2cIXcRW3Pg75f8Peo
Wi7jup/vGB2TycJk3aMyjL/FJ7UP1LURADqNlRYocDx+yMsIA1rjDhDDmDn6YfcyH1gEJC7Q3qnh
DxcsIyz9+RYrQgtD4bBuuaan3ki6qo1VbbiIO5DYrQHptLZlgbjcyD1b63Q3d0u/0Yym0nUj/68o
XZ2xzEKrg/N2N7aqVhmNqP63WQesJCQEtsg5hu4zr+N9JxRsAJcmya1CrfqjfpXICVMxciWOuqss
elut6TcucdlLO2sstMA0ncScslIXyp5YpFLPfwtKEwrhzq1+oH2gy+joXYRjonPLuF6yw/Mk8lT8
L8La+OVqN8XDWzgIhDijFj9Mj9Y5N/BWI7uYy6cJEhtyhSjZAomBkX+8/hCG+ffcqfTDi5I9MWEU
h4E5n+pn1Vl+YHu3TuxQczxVtEaN24cNHL7Iksnry0TPtu+l4nf1uy3Dc3OYW0e7RErtu+GBEMbM
mqW8ONw3RY45OID9rpumXO9eHvc49Ytp/9xTbfIZBSCrlLkMEJ4gbAwEy6cjIvlY6w5Gcy24FVG7
Qx+d9of8F+gNN3rKseEmQU/h5MlzR/qJdwUTADnaAtp7PLdHm3J6TbxP1YbFJtSuqb1PlO4MmIq0
hNnsBweNO74vgRvJkIFqPJUtRFDIFB4+U5e/EdLm1zVrQ9HM9u6C/Ea/mpUy4nsTWhTxPO4PFvt8
qkOtQh2fE5hIw8ZeClntHqnqQ7LHhf2dqpTK9NLiTB8kMA8Gq2pH8ZnFPGxh3f2+igtsQJFUkLVo
9RGqwG97u7VsB2kTFwHAlytdLejISUO0GSa1sfTIyuINtVlEXFyxVSxGWiPXoNpZ32vOOsBuQV6I
ow7y/PhAiPVrh+LbViiPbxlwIB22XJDE9xy7tYA0YEnXOh+JyilNZDE76LlxiddukZvF378/E/Cg
/nTL62Xp9EE5nLfzCSpy0ddGeHq5AMiv6eoB6LZGzAysSb1UzRjf0OzmF+b/JJ5e/UEJVLY5JGTh
tVRGmg3DwOI62Nr4ZGOSdpQSXbFNmH/TugCyeaJLYSyH0jNmO1Ih+9K0ft4XnK2Yn6jqjaeBXAER
GGBF99Uwnn+iWrWgFbXI6GfrIbSO6bmBOr1fKwnxHMrHInotAkS16Y8NBUBQGoDyUR8jk6sCB4ID
RrmGE0aXDwy6bQdHcjsZg8jZEYlCtKFazCAQOu/xmzs8aSicCpHmFw1n7nZ32SxvHFdnnxoXekTL
wq8sGnToV9ysVGe1TfwIsY3JKY4a4k2DjH/EZIX6c71EKKHlA9J9+SlZXvUWupmDiBmjtTizUCSj
/bO5oJWnjCnveE/EfX9xFN8dYv92LWs7PeczU0yFV4fUEaLR2KiAYYdvC2q/fBkRpa/gFEcFnrX6
NtD9CP+Wu9qFl942A5r+wJJU8y5Xw+TW12sKYWh1omyGQYIpZc1WU8vojFN9f4y/HI1AXRIKZSh/
UtrOhaF/NahAIjvRIhpvzlR0C+bVrVEJz+9fMNlmF50bIZbFK1vYaE4wof2X8SNXh7Du0OBKsQWH
akgt08TipckcnehaYDNG5Cp02b6yt1H0UQiyzTDuRjxx/sUCyJ5ivjfgca+HmiGxPPKCyaHW+cVE
GrJn07Zgjq0PXDrs4cyBVG+Nv77Vwu3tLbJXAUxsKUZgPaCwgvj1HjtmEAu7CICGKFdo7Ga9fNBp
aHpN0FENQdHDCukqNNl3aJ6r2ESsjXY5qtClhG+tQWjA6QoU2NK76CRHDUHND7mCKNPHEBq5Tluj
8ln44eNC+bjgrVDJqubVexo0ffGY7tcROivffMcRS50ig2NQAOxknsnYGsg4gjut4p/KB6+z20Ks
9Ph6RyyUcTuxGkLiBgWSPAj14m7NVollvx1I/FT3UUeJotyLXbiMEKNmMYSJ4LtrQULcLAZUI2zb
wl3n7JKL/sFUtKj7lgBdsuBBPpQ4Z0I5ZZhowyYdz6tZS8hZzPnTd51L2Ds5oTesnVpOH/MY0Q8x
shQ9UO6j4lGiqhcyRHaF5aITj+j+V5jmhLr5YrAeq04TIClYg48LMcpdS1w88QntMx+nUqiffSX9
NyVJp3E0UmHgf6l8hMrh2rh025YkWTm5skQBaWg6spmpvlYsY35gPaZ7xYymbSBPpaLWIOfCbACd
5/UxtqkMHDPgEt6zk7xknWF+8UmyQO02+m/ryTPZQKXaK0iKG6n/i2sunComIB6x4We4Yb7FHAoF
/wCrLQDKY6ZzCj53FI9n3/vT3mHCXV4/SWiccS4t4gP3mp673YKo4lj22wYyz9rFgNFXQHdpYGId
di9b71LzsDY/MHyKbb+S8AeXHwTzAQA2AJmRzBKz16QLO80AX5m4AUjkgk/Anh09vjK/t9VcVSzC
QgmVqHJ/1iDryKdFwut42ezaDdB9drLyaNFNXQKOpklEKNQSxP3YLmL7CyaY2eF560LUtGe+/IOJ
m/Gn9sMXreinVpAya3ew02Io/07Qvbp6CLyVAkZd4QtEZ0prSEuNMK3d13yV3ZF1MgesB/pUb7qJ
QMxutJDtOjcKvzNpNwNSFCwTqxV80nH2S+ChMQiBh7TWQVdGId76muRgXi016hBPmizvhvQ2Ljn5
M0stxan1yVwRPJgDQrhYadYcvwiAaaSouIwTWw+Hnj1P/XwTl7JN/+bAZZNx79lQIwSy+vmXgMJ5
bj/a5BsKMEFXzQO8mrLRK2QASCqpEngm5NqUtnfcflGIYM2HS+qBCHqIPt7UhZDy3vXclfYKksBs
MdnV9yp62sZj3NxykKelolGvgpccTsu4WVfROWpVDnQXOLmhI2k1xXd59IaDHUS6X8u4f+tDTgQt
Vta9A+kim0hy/fZuMSP5zJj64neOQ5A3WlhjjWGMmviwBASL++modRdwdPN190ltC0pimVOrNtoL
GwzwHi3gOQ93cGDElY+miOanrofIl42BgYmVGDZIMmEs3Wjo/swYnbptY8l7plNoZxzoaST+eZ/N
CEIQ7E8pj58TTVPZ8suTznMP+dK9jzitAAgRjDshZpPc9e8nE4GSTaQFGsByLLIZK68e1QUwucHo
QyHFEHNWm5hMz3hNtWGueUb1po8vLKTl3ioFoSATEIPxHRqG7vBSm8qHkmotB5A+sNu5j6tcZS9t
4bWnyyD3Ra7lc189d2FuVIA4LHHfRrAOmsE2HmM5gX6Ai74U8afV/+7BogD3mH6+MS7sMCDMgcH7
5WnQbL6cbsBb1cAeMb2Qc8QYenxpoP++h7bC5sdRpgmBz9+APu1Xv9JkD8+Zf/p2DDXljcFs9QCQ
RR5ju8nhRM1ZgFLZR0esUyAWgF5lxJnsBilix+nvW/h5alv3IJ/n8KVrhh5lgyiOpYCfGbVcp5sv
1tgEBbAPwJVORsOipsAF8PTYVs2GIafRdx/YTavoq3Oke8WMcI1PimTo+hR9WE6UIiiaAV1ofagY
FUZHxyQ7V2WpFddTFloFhX5NGrbtWEjLojZKotxSSRHkn06XjdtblZI+4dqmwfJdcfOVqluDY4cr
vta+2pxsfqjH3GJ8mAT4jWvbh/VTGNhp9UAB6oUA+kB5d9kHvfpgkzm7udvjUvsZzjzwamhgqsJI
7FCjm9+NEZmGqKBioMo57s4ymHTguRU6BbFmbyIW9q3HNoPQ0kOmtGwWMNphgLj4XWkpLGPDJ9JE
48Uvb2M0A3y+W33pmUqSd6Pmpt6aX58j+YbrSUV32rr3YdaVBGHCzZ9bTfutWX/wtp+p+jzR+juQ
OWyyx0cd0Y0M76PSC5I0Hk1tlTid22SLj32jfpkXWF5dTAjoo9oOkkvGd+qP6MBiwJa5XuvEJ7pB
otHS5lqZ735Pts0CWDcDqZyBNBYlR+a0NmQiSQQgg42SVXNtLYeFo/s7HwsSQlH+5TyYBtjbdGM6
MVseRK0bSoZrAU6+u6kS28XvWBdhA+x6DXK3SoLsdfMp2s9sbPITxRzYpr6KPthJsL7g3R8o6aAk
TwlCsAzF2EbTAjPeYXGLNB52YHQeB/K5rRT9jKCsvNYIVgdXeQDnSllwpqC8ZiHwOTJJbLNbWpsz
htkLdU8Z78oUgCLYr1ME9DAWgJoBJE5OoDt09K/4ggRnExEclGlUNqhqR/NMztn0YNELlvZNByXb
XRQfDAiubBJdOkTu1NWfMYoAoy3xAN1z1v6A0y8XbX368bu9DkvcZvt2pfrnWCgIfSWxkv1NmIWC
g8uudGxkTopfn6T/7+E4BW6cLgbAK8BrpywfshG0s6+bsoOVol9XR7hclqqbvDOnw9bXGvQv50ZW
uQLdCTP5lY20iPF9e3uAEanufbdXEh78vJTzln71VppkMH7bPvqYZ3QYPhpHEFG5ih8x/2Nt+0Ub
cDAmhItp9QANLHGYPELby3FbcYIAe9yODAY70ZSPD0ashmtMFAjxYlzuzPK09RXA6bZpyE4TUcEb
FllK/M5fXws4WvKVQ+ijPH4rwFWHgX7+MDBoaTRnG4hEE7NtxKFGaLjLxQweuw5ojorxzWg633iZ
Kzia7oIR1CkaYp33uV06aVbj/MWqquxhiQ6xhh8jbLT6rpDRFYcutD+39YqDHtbfX5I9fpAQ/ika
90QyxRfWUyllzYZK6IdXkbEaWxR3JmtQ7SEVSgYGULG3tflFLR1CbUbRhqcOIVnwW+hsGMKjMuVB
3txp1aM7QuJdK5kbpxDnIPRUOzYelTWAQYX/7V2WkBYO06IVmGfRJPGLDkMA9aeMiHcOeKoyVTO6
U3GOqgQGRtBt2PZ2OfgWPXODH6xtFHCFObN7vzLfo50TncrYkTQ4gZYx+PBUHaBFuM3O2EQHDubB
qIYoC+Qv/4hmaibky9I9oF+zLGQJ9/1PU7AHnIqvpuwqft3AVSZ+sCjlLVVqGbYmqzii7239HgAL
7HmbSFgtTbhUhOsehZB4r90JvF5bPvs/iMHUgTR06FMnyEEzrCxzPIEjQ/pTJ76aWNV7qvmuEY8c
Pwcd1BFnduyoZfDlC0cvXttHGI5ECCWzQ03ta24OWZyW0yMcvQtj5PxCcaTpyiaDStIFUWsvtQPU
VHa84hIa0SlEMlAgYlRaf5R6wvRypJInLQpTBsISV/MIeg0kJdEP3L/+B01BwYKu1GNGKVE0Gm/n
DRxIJOxgkBTMETucWfPO17vRFhUodf+/ZQa8Ob7Y4qAKfJ013TkVynFnYN9cvgYf/ZScrHiXiI/9
G96Ij1uKa9DESQeDZE/h9dcuTxJGylkP+aydmAIf7FkfIZuQRfrT+HLf/eRcvbL84xhf4pDFtHtV
2Ig70/oyUXGA6lAO3MmhhZQsrTlvmvWibzxIj5grukwqS/LGfQ1Lc+dsniM1Ewb0kxMqmEI9uZ4k
FQjhqYPRVVNcMXEVvVBbvr/+cZHDKaumID9XE4jAd1LKRIgd85Ab3OWJBqJqGaHePCH/9bhQSWN3
9fggVKoooGQfEJdhHWBqsUnI9k7Y4DfdbB4fw7MqyEKZcmN7KyUQhHO7NbnKPbI2c4Rg53t8ztzE
Tr9zl6FhtmYSW/yCC0wVtJwip3adMfZhP0IpRHC769JBFJ/9x2oB21hG/waZNJ49V5wFBA3XIPav
GdzgF/Bl/5JhtekXN1h/REpu8/L/b1Wdnjj/yDB0x1UmV7EPXj47pJbOxtfiglQUQxbIMwtZ22QU
y+8ZL7CG4n6GmHCmcYCWap4ZMoyuMEQcn51P4ucc4N+yWdHYdrbpsYXupNSKHIKuUgz7qwPEp+yT
uEZJtfiBEjGAzbDcj81K1ZiYVx5kcQs+9djSMFEiP7mOjkBURChs5rKkW4++U8OSmEvXfy2O3fMh
RIcuogdf4E2OP8LTF72RaHhX1uK7TnUMN3swFAmea1LF67IiJaoQZjIilOjPf4UU+fGRHKNEskvZ
qdkN3xp/aSEy9gA6eGiXpCOaibE+JXrrwYgXyE74Tv/3O7RuO2yd1DcEuzaLYlKyw0Oh9v0Q7BfT
0t/DV7i3wkBDjrSkAUTK9E6YNVlJceqWbpyU2E7hYEWSUlbV5+0ODKpiIBKbTvD8emCRESZeY3+w
9fDmAATn9h05KPFWmTbt0KvHaXu9AHmZfV4GhPw0MHsbgcqFoPgToLSpPTcKbnIUdFJHx3UkDNYK
k+BCAQIF5QhT2tLiu3mjtZstt7xlt2kCcP4Cc9M/+6NLiMTYQL7yAaF8OYJE/k1+ibmro/C46/eI
8rU4yWqKa7Be13Kvwn93RN8QP39OymJIXLQ/bNDgBlAxQSrFwMuGroHjibc84jHeGvJMB8v/0aB7
MMJQpbyCNg6+IOW/aseNnGoyFfBEtE8MdbJ2etyfNp1QLRcF8D5idWa/y8k03iFYjKHfGWVHWyo1
qBG2eVTBfxm40I8DgFGw3ZmAGEeFio6dgZIO2mQrFmadkWvxa7oL7A58EECTaaB5qDyv//odhV0T
TpvJ0+3lxVd8mfRPBmTiNknPCF7y7YwiMKcqQOvSGnZR2x8c276xU5+Qxl2KaiJR4Xw6NA74E0gH
gP+HjCC/b1PtBnoZOThU4dIEr7E8uMmmKezGZsZhaPXUWXH0nVXLRQYsUTtipIpgAEcqQ0o3VqSC
TfUurP69R1tbVIckxFjXEvPesBTKPsO9B6mYh7X57VqbstSy/6VOyUb/Edy7ud4efIPQQ8EQ1q68
JQsVlMrPfeBMRYAQQmNWVEqvM7xlDU1DUxaUzu0t9wKNHWmUGpNJptRbL+4edsYjC3b9frFy/Rdb
o1IRUu1fVddlk1KSw+xib2Mead9gh0eRDW13cX8KR10y+/Jz1pQSCh9USJW3Mer5fDTm2ht+x5IT
33Pnp9xZjV4rz4numdCLYv7beNULb/nosaVYYKdOVMJg/ECRfhe9xQ3ZSwXTBK0KvSzWJhOYAmtv
h1kk0WeiSpTKPQUGiuPbKhMjMoGULuHlLY1livrZAqDkKaHgzyKtXInZbYIEcFa+5m8Kh6rENDJq
Y8QwkC2LjzenS+HVL5stzgTmrVuCr2/8gS9AYVaLKQYypVSqPt0ZoNCYHVq4qUvXb/F6w3Y4M1h9
dZrUJ9gvg0/vbv4Du177VfwAHH+qX+EFCM8CoBODvKJ6H4UW/mfkIyKN2KIxlOpXxnJU7+NxMeko
79nW9X2mKjHaymRDN/U8xEVZlQGdakouMjRcjVu6Aeq7d8J3z75I6e9DJJVMiTIIQui00iVfi96z
8hNNWbaPHbGobSGNn/rdXiw1Xv2odagEmYDLG431BfPnWcClVJf9YYOMiSN8nIEB6Jt8qTpuBl+m
6jUbPgDOCs+qr3QYqSo4UhQqeVtYSWlDOEGW93+YP4NX/TbSWTCPGkod9rRMbP0mbEeWd5GAmd55
S236f/8AAJX5hFstqtez0iI9PfqoH/iMw2ZE7Fwh8+x80M+nfQS9i93SdExxOrWnWfDmgYR4bP6y
0CxJm9Nc5VHGxTuFA+3H0xA9LG6NDZj8hVpl1bgIZJ5S2ULbxIPxvUJDC80MsPzJjlahznTp217p
KQ2gsqfAOT29U83D39HK2fN/wvSeviS/B4RIA1kVSazeLD04kZMmddh+tvA67DytPUWCU15brPwa
eYuXu+29CD5WuDktUp3FCjRckPBrFuoZed+xGv8BaIwsBSaJIGrJTGT5xszWgcQrgu9mdUSwQaje
T4nAN5HaP0gRBMR8SAdRidZer9NjEaXyi7/DCu1SYe2OBgFn+nDJGDh/rrXAe+ZdqFraMGv0E/RO
lRDhErIYeOP1X85htr8E2+dHvcZng+xjtRLdQfWJRG/B7ugWAtpaMx3G7a4yXLW+0dgi1TNu9pQG
coYIZ4jThvMbfUBjYhBCe7Aje09ldpJcmtOiQlBxmQep38xdvioVhaEG+qeoPGIXg4kMRcmqjHU/
4kzYa7Ol5O/dshBzzhpqkLxnTZsLFnCjECSLE6oAtMVqYgv/ts+QTi7EnNbyVizV98d4aHJjZO+/
Jbunvls/uQmcMDfj+0i+fkGLttz3tQEUXN+X4oSok0Bta45eXkKmjxObqqcBolsr0vlpQmyJCqvO
AIY0wmCgXVetqMiB4gd3rMB6hzcl14WPbXLaDBy82uUwxp1fGp/jmDyEO/lBAM5f40pjnYqx0O6/
1QcfkLFml1sOGRw5HLHH5Ej4Uy3Vh7jCZYUY0ffGgj0DOThNLCO2LWIKZxr12B7L92/gct1I+3BS
tyX+SMpR3kfJycTfce9VPQtjrsW6lNJHEzpBa1VvSILc53ZozBWqdbWdZxpEAZjFAOZ/Fev/YoFO
bwpUd6reb+vnebarbTwrqCaYulfOF9g8uIS0DzKPfzvC2h6+Tj0cGktWnJQggvwbc/i1oKMWgmbC
Yc6SpQt8EIIqKzGTcyOzkpDPeVk1TjG1UUJmahGF4Z123q6vAzmimwWj1DDWdq9LgEeZc5ucTMsT
7Ee/oGzd001Hc2/AI7WqqF4ucNFUp+7Ubld6VJ849ViXkuyGRfG3E4tk45IpPgDWyGs/IWjfbr1S
2ddENLua5V33iPBPM8g+5raDxq7sgCbf+X3ExGq4UxaDMAzHQvVsq0VLielWV1n/M8B/RkWsU6jO
fnHWXBtB3DLoI5CMsN1sDOdTns9lTk6YxI12dDgtSM7qq3W4jG5WVTIgjiFsA0vP0yCqnOnKG5te
8e9Z2+g6ekxAzcEVrruc+jVFUBcrqY28JPeVZaIogkBrJB8nujjvXBsLEUCFAupcvcfv9HCCPkpt
dIVbCFocTjdOaDKUxPOlTxoM4BRX6RqBZN2A4eovhrE54pYkHFnU6fKP6gahQrfWcf0CrIMz4Vmz
mXiCalGMxgEQ7d29SekXSxkF72KnD83LO1NHG5LQwRrTGxcexZZpZ4jKHI3K9hLd72gtVi/FCpsA
47FiAcdPEWPoftEyCJ9t5ziQo41TEEIXqY40/sh96h0sT00W0rOUH/1ftTb4ahm+tNgro4eiCJg7
3RRhc1oin2pWPaaD85/SQy6rZkytn161ZzAHbWE2c8hbpHRt2OBHu93BBfvfhIn3swX5Uhtrwu5l
7zUMrnAlveF+u5q2WHU2gFK52U0Y9bkqC8gdzfbjnNS2bgVVAXdviFWM9N4ihoEWp1yPK7SNnUSa
UXz1OqyUDrhuwwe6dZ0fDrv5gjFxgs9I4bgv7Bk/IDiYAmX2WKrh5DWAdD95UyFrAvVdzfOYDRO6
E8+kgsDSQcbculnIAgUslpgE8nVI+L/3F2x3harIgqXdKJZ+opxuEq6I67s5CaIhyOFtUDylB3p1
EK4O9qGDsFN6H/K7dwaMWM5P0U5UEKfwgIO3q3SO848S9MpP/dZNvYbOnyqITFPtxQXi1TrAw+bD
JZQDNUIkGIkX9l5etVZOUpGn5Bpdfet+pqOKH3lksEruFAtLAxyGLD0GOEzYB26EydbPE19lCX5+
AQDesg3GiCblewyh8iiuL/cinJg8JSAJQUD3jBFoF9GtnO8JnmWBVa5+4OWTk/rwdEsyuHlBTVpt
Ep2nslyQVaZe92CRmmtILxi/kXUrTMixgIaP8HvFIt/BZ0FcDFOjxn+QciymHiOlXnImpCxOlr6M
DEwGEoIrXwmS0dDH/MkOgTMMFnHkIyaD1hwNeAy2RdmmzNikRAj6wzYE4KBMOBbfhpcWHE5v/3E0
U16zMC8B/jogSJHu9BCspXytdc2gBEx0f30j2uueBBYq0oDm32QnN2oE0u/8TXqk1SJkLDCf8ghO
8dvA5448BCJT9gPRnPji0N2XeAiHhJezJbKz4ZHHvL/yheQdXFFScN2HmOwkJLG8sQFQ6CdFAwUW
aY+6ShIJd8nZ/GiOaTDqQ3hWR7pIpiBX8ldxxcvAy15nE17sBkEcN96QWU0FqaRXakyVD75uh9w9
TFdsIAwU/20/PBmtzrU2qJCd8Euxj5dTIW4gXzxpJlZTj0BkVkuDv/pH1mtlSuenj6N6e6iurcXw
6FsofN4UCqinz9fnlVwL3KDMdVI8tW6CygPhw05GmC9YyR2VcoochOjjyt54dFk/3IsoCDrVMnWv
80kiTAXkcpPv2UrMAUVh61dKzGaJDD0dQF70zh15s98KpVtexyY9C6ts7yZntexpqgRVyUMIjvf/
PyPK8vbUxZrvbA0DgOzzWZ7Q/nlvmcx4xj2VRXp3DgiMxLmI8IaYIErjJB6dekIlKdqL09g3DUua
aP2bRzghM/ozEMnb8aFtH0IA8CjUxb7AOwNiw0nof8zQNagM3gm6telmHpN6cgY45903hr70b0U1
HzGccoCQD2gHzI3HYPglane3D8J1O2oSxs291ZLSfmWlu7uwHi/Z7hnC1kZDghkjcOjkwSNtVLXp
rl2yL+oh9mBon6Eqe65iNwE6Qj69+bViHN8AWuGtXns0xy38GdgtFCKl74NY+sUUokGQlD31kCah
6YY1rzoqzQUczPN1Z7SsQMm4AtdZOYJjNSpAlXOb3WdnIzdIPwENr0dTt2aht3zNr1xnv4fmcCy+
6cmYUvUFElxkOOwkMh7kgK9Aw7tdfon8kTHQy8Dy7gKZCWCYABEmgD3dwEzImcywHsc0n8tL0Ce2
qqR+tpkUzX7wVbCpBO3f/DeMX9UXbfUzqRNudMHh5EWRsxvRBdxD5eci4m262pVXmX6L0e+AMDxB
JiOi1DsVq/OMPuPpySi59Jxtsfs4i9o7C0kMrspYaAFmgGFebRbtaPwWbTGn/MPSvgdUQMPc0MJ8
l0xyFkoxp6HJOY3NpECKVHm/LbYSiwwY5x2bIW6YR2FU/DgjiuiNj8v8TqlOUhojnunYAU6REJyd
swaG1xW/jdPH72GiIXztmgXvFOqAMrHlcR+UszhIsoZeImDTLFSnMiJSp9pDNz3ar7H2oSumXXto
T5ihpLn8s2cI+F7dC5wzApC2kZig3D8OMAiWx0eBC1Q7zG9cZEm6HtzWMc5dQmpfOQzFKuIe+uDb
qRYaquuyKEqUUJ0oS9F++6G+XTMhQvdIHj/Osp74g/TPHV5skIpkVwCwSKlDTalhA02xFosdi91l
O+59S9vpVNxtKFNXBZUYwbKG7Rbddu5MVr77N2l5aySiriA81q8hodOZw3sxaiIopZnfYkRgx6tm
1bJsg7NAsrUt/aOarP0AQsI5JLVjrIBHnptotJXBqc2lra3KIcqqWa1cboPop+7pd0ghTNGyQgqw
7DXwrWRRpI6U0Zlm1cN1PPfxr+WAYooHfNfZ5pbfjuhvrvHuCgtKBWh+NJWPfoB77xz1++GXw+cK
ph3ZBMNs7dtTzCDJzLSYjhdftRAYTYGGHKWYpu0cNvCMopQ5XL7j8Dqt0EzuqOtd+c5/6cMchfXu
yq1c/x3PXqk0/sLGhH/rNqs+e9jKVUsv2MgE247RqnnqgWJjhL3CwKzLh9+ltuu+emiSEilEwuA8
LGUwmOVzZ6BWMnurbMmYNheov/q5J7LPpLOCtlr6EO2d2bnh/7KYfHl8aknPSD1Ep5llnjByd4wm
7Fq+ciRdhp7WM+cu0rOGvuruja+IpCh77h+Q0iBZlo8hMWj2sR5kWvmtzdrUrJrvyOgS5ETor1De
Ze5pgSJL5zDbIZPleJ1isEAyDBkuu7MnScbXwEqb5ULIe+6oKzK3NHcyQOe87w5WuHgwqaxK7dwc
EGqSGIKzgKzHHfmVPY/i910DEStyHGcn1y01oo4txkraFT8RupNgjWH4EiaOXwX9gVLH7JaMW1B+
mged6Dv59DGwzhUl1CfTL/J1YY9EBjKxxmMd6p/xPHDyaiyurM+/QtJ44e6cJwy9IBNFeZl31mTB
814aE/RB3IvRDIYJHTd5UtN+N9NGh6b7A0j32LlPtVXJDgmbtEOl3J9923buYPxSo8mmdHKU6SZU
xgtjS9qOqGsCr9BA07BOlx/TQSITV4DZ2AH/Ihe7cZalKg3gCENT0KWRHamOirAr3JdAn/RuFc2U
PLxoU1Ay4CzAHCGjtIZnD43cimnDAHQVCNddPRmfICRCIYh7E/WT26nee7Zmt2lSGubdm6wYIOk9
r9+I+NjtkfTAzoMHrPK1ZkmxWYVkr9nrjdAU3hTKD+pzqTIq2sT0ZzDgnwaIvxmYojvXBOM2foqb
IcKUoJG9xxOhG7+lNcfXHpgBSdjMQ9Z3gnsXpVI29IQrQS4GB+u7t0CggzXDlV8gBTewzibkxRyF
b5fgPe5t8lX44QSmY5ubbrJ/veWqBNYTkCLF6csETjhQLU1fbBpvyUHmmzrpTWKDrtVafJXBs3IW
FIuLyJRymDNKqFi6gYPOvp2PkHTDWrF9/EijZBrfgLQHVGix4BJ7LHx1YBFNHsLud7jEDzrEFi5v
RsPz9o05wciv+pFN+AK2ZF4PBHSRRCy3XWqzEib+rBOI88/FFkKosOMFpyY1R05U0vy7VlHkNF3j
H9SNfqQmQmb3B9NOgF1+UTxKT3T6GAoaivp7lCS4N/253r+E0PPuGJrwdLNkoa04zOKY1BGE8XyI
KuCgMIlZMKjjD0sPv6aW0vqlYUIOGO4mX60iiXfU/xOXnj5L+XQGVNMELFbjnkKiBNWSqqrNguwr
wjVX7s0yG7PNwKyL8fD3oatuBOibJpFMazjCLN57wU6pPJDnY5ImePV9jgN36PTNlophGPoWBcGf
zaPkORkyu2SHjn2eDEaobOeLmIY8/FQHQt8ZutBlwS68ND0pXohyPlgAcGlGHCJYX9CdtbUXaBFH
3F/RJ2ZAxWN+OjfvYE65/5dywwMaooirPc6cDwwgAG2Bq4oG6h58R8fu455SZ+7uNQAWco2SkA6l
5GdoWk7gmbRiBOlEyBNLYxR85xj2qnsJYp+IOdBAQbL6uzKNSBqPQv9kCPGFODZAR6grllmXq8n/
JFh3AJ0B9Jpo/F2Yf7cK+9dBdYXxk7Y7Z3HmMnZoRqTvh1TTVHgFmHkbsDdtGmfPnz062pwhhYgw
Tfggrx2o0sPK7UPTHfJJmRB7eGyiIeLLnAuzRsRCSOZQTor6YMwG2PTGSqAmXouXZa/U2lN4jkWb
bw3b4mQbobNjaYLr8eAgfwVDCVai5kFEnOcB/fwhmWTHVacPJWM9M5BrjYmzUWKdpOOJOvWiM1g4
/H/o3YkEmyIws3URdL47GDbxUDHjLWOTojy+gkpj2sFePeqRvXUG93bL/NJ2Q5YKgIS5XBV10zWA
6po5oeXYMIsMlIcmcUhU0JEUwxdVSnDh95nex7c475ry4RO2GHY0Z5RKHSbi154KbCrU2Ho0MGZr
eZn8Mz2ADMEkI605rFqaPdt2kO8w4R8pRwxFB7KkO+7PiZ3L7B1zF1MPJHCU8+Ht6EAt61v+rOOf
V+efFANVQhFzJ2QqtpvBeMtPrJTiFTTKRWxHosbtE3FME4fzWr9xoi6g0IB56UhRJKfa7H73V9BT
wNviQDyv3PmprH/oeY9QsOj0CqHKp7e0CjnNrwuJx72TJURDdFBKT2lo4oh3aeyUWxNabGbF+2zS
2MU1MXIIhFyzpA0kzE9mTpC9S2RYwhxTs+xS4MX6IIrdq2tXGVGeSlKkgYMErVnHm0g3CkqRkDYd
LBd3RMcwIfTM2+08kCdgEekQ7arzn1+KGE131yRx20FHEN1j24b+yvAGbCXDvpL+MuZN3ciox6En
i/QZHFdjEFlqgCe9KO/mcdam1bIsxccmfp3gbtkoqOR0rLt8n2Cf58pXDS4dKr2BjDGCnKXGmhIr
8ooZSXKmh05OmwU7qrrCHKkBcIMwV760Dxh3VzpM1QiUQrT8tL1+yTEv7m2yBCanjJGj3h/z8j/8
3BqMgN8gpzFxVEm1H5k7CIzBpx4xYuT1+mlrOCkw/yzF0+L9EDUK1lwglTgjPCzTGEAmRMmaI89U
3Mvf0PitFoUsfayq9iADePBCSyVH3PYWqDM5tqGA2dyApi0/ev+EYZ1Y/8mk8+fzkW3eR4qKG28u
Z1NsXyIBnNMKuks+fqvO2nhHERszCTRBkTp/9htHVEt8KPXTvqxfqx1KyBQL7f7cNTuyr8aFbVyC
kH4bA8zs8/Fs9TR2Hm+4zhbmZX1PIh0Jyn+A66SeYvqRHb1Q5nAOD01nedn56uZ3UO3tA8X5WxxT
Mrirp5O+/6IF7bZIEuEA/X1311hMZ8r79vcPt9tNobDLcGccXN1XEDTjxN3RKj7BqsvctsfHh7rX
abM1OSRvacmYul/qq9dUIrnnHnAOiRIdpMgzCMbcSJrn+w+N6jVdERdtvugTgSSo2vAqdZrvoJim
B8pqFGDZ+6NSc2pzc0Q3C05FDsGpW9HM5vfCx+wZfrYYEREIDWUlKd6X8R8hXMPWLKTWnvjYudjb
JtTvwrPbWk4bSRALYYQa9KCDb6fLiVq/qo6pZh9GfUaJ7ECBbemLdWIR3ymVKfsofC4yjU4XOqeu
heo7sWvJBQDKW37ztnDpAa5bQ1OARGh0j78W7n3QZchauoWgbdJkfQ0PpWrGGtQxbGt0+czls2HS
dNxnOv0XcdBnPEgfKBCdYiR8rW8XMr+XygjMLrvJ6M+Sus8zfuaD/LmgOia/0rb0Lf+Pr8iYauGW
cBgMQrLpr1b965fej1GZ5uOaNoQZTYqCoWXChf8X3a/HEoWkrnjWVJmS2E9ZlIakW7YV2COX3nIQ
nsruANj/OnX0CzCh5pAXq4TcRALcmRDVcbQ+uZRj4tC8ArA80YW0GXip7k+Gv+rwBLHJbfVN64n6
VOxVpzOCn4IGODnuElJJuw96BX5in38pTRde6Q9g7Ey56STtYCryWmiV8K+TcS3Q+I1pfs45/CE6
2TrurCePcvbONWrAogw7NZng8HggnRC0SDMh/QKx3BHBmWd1RrtqhnlDuUumhg37dN8phSlEJ3rp
Nlzt99QGbcPJ4x0JrRBgYIJAVHmjq1PsdHw/Ld7KCtGAShhPyT09B0lGxn0DuPM4TEjc9nK56arn
jnJthuO8lTmHT7BHu+WYfwlNfIUKD//tfl67nNnOmrVfIg4JExwphv4JrJWJU5EqIAFU47dWDbku
64dOQuou5MxjR0CxErwqmIM797MKjQ37x3YR7330exwOynDqCniTM5dM54OjShs9LV5HiZrdus98
kNsMHvka+u+YBrPappHZ7BBTL8uEhRUWVacOH3//OoeePDfU5VJx/C0vpqavFm+V7PVGZoGJa6uk
zMcx2GXr80bLxUxxRHB2MTWijNgstGyoz1cEziqfA+bsZDbO/vhC4YJkIOIWETFzi4di+73gTce6
F24ShW2pPy4cZR/FX4XuN2lctMp9cIIpOPkBgauf4suf6BFUGEHBQXDipMo5voAXETFCJobxDzwt
huJBHiQyEKl+8UeDyRLJL8XwjRu/MKjH8Gt7gAVOY8IQQManhd7X3THkyV2XtYev3jV9ZlTimyOz
lz5hYfOiP3v5MuX/iQ1FaD3qZ9Xjk75eXS/X3foqXX89ybPUF71A6B1jOztAjVNUIgDdMni3XPSA
EHpwe2K45mweRlWgiTnxEbguXWRLUQEOkfDFh8fS25mWoBYgrtGfRkaj3U/KqvmemOQp5DQI8TB+
Zoywecw/NY8srZy9i46g40gXLfWOoxEMZuRvC3N/EvTY0zjY0+c62aW4E5P+jqQDNe5X8Kz22a1R
tjGFlEpA1ilkDpAFHM9o1KZNZXb+e+YtWwbCwX7F3Ifft7Byti8GM9QVKSjEMbQy8mvRjPR/b1jR
en5syIPZGRV7EuFD+xfLc2Uf/e5Gr+I6E6vwUq792zLe9Fr6NvYgtulM76e8ZknrtfIXyjUmkIqA
6f2oX3MKY84pqiLoqrn5/FbUVGPzzJgt+zfov29zjZIt8y36ee3JOY+BMRc7AgIodVP9NmiBvbfO
lG+m0kBFoG5rpS6b1HKMKK9iZ0LxZ2aiIE+CdA4/BNdq82mJekvaLC06DcxDJ4OzxAfNwswO36jd
HBVDuME3AdtOMlsDmAogjCQOyZKtKayl8gPatshXZ0N3+S3fq3FfIbZR1GDSl/eJM98Kx5Wpkbp4
kv0pfi1ahI8XT71lyJ1busaMYaQnOUhJsjYpNOQCq0kuj60kDjSNhdK8Ya2MPn56Umr5iiuZNVxf
sF41gnCRFg10B9au0C5nY4Oi7TCqkB8KEuViqq2VKTcVVDUQCiCEfENMvnwdIEPAcCZ/fa1bJELZ
wyjWSRvEcMTFyHPkg1fel+bF99dSuC1Vq+sWwPQz5Egsj+YHEFCWnX3JQb6SfH6eA4+oJHjKN8Ud
+iU8DvYPe8JMJaKV4Z5n32zsHeDYvpw80JOgFxFlmUVCpprbQqqckfzKqSq7kBLjiX0sRUQLmEjz
bkEwth43s/ZH2rPyrgKyAuBhdWrBAjgBm0fQ8MMAn/eMoABxgI+WepIpn8d8XL/08Rl0pgXPq0E8
4TGjNUzKrjYJdEpvtqspPk96qJru1c47NrhWlv6eBjARhjsEMMreVewD71uZ4xZZ49F1TxT/HXI/
SKkc1PpUw9WPkza1GpBa0z5gJTxThkaZ/pcw8AZQLE270aj4hNx+v1W98CbjKYKW7XgeLfORb0Vf
YZEjTrtc32vomrN3lEY9gNPuKfSF2H/S6LBzqt7d8WvYUsYDdB/qdEpZMqwXVo41HhrE+gp1Ez2E
SIld9FzV6sdepCuz9JRto1qnm1P6r42b668e2HAU0ZzlR8c1YEMOxH67r4e6IZoV5wxTuBHY3i5f
FOsfFPqWh5HhFfO/Nhs8lGrVIyfShYJ4KH0tnuR2gi/upZmVHf59wIyuUjw+Ey8HgLQLL3bddSU0
aBzdsXjHavB1E7qu2P+ITHrcPGFozO/3KsFOBX7oKXra4uXVU64jfX9uHmCCsOXwQT/GvJkESkM/
71fdN3EwfamOvTHD45vabKsRN7oa7140yA2h9EnhaQzzMCocsIkhEvafLvWdCFvSh9zOcxislLck
zGHzYB7+VLtlS9JbUHmGcFsIxqqUibUk1Zo7oWHYjN5N4LZg7LA6Ci8ZJT1P9gae5e13pKCssHxN
MRqld3KViVL8osQdv59h6/q7iKu+pH2u0R73W7TSb+k/vci94zh8jPkAerwHwTno7IsNkHFxYGg/
6jah5tQTtLsR1QFqSbqHzTySMhFc84LJMFZ5zxYpzFoySlYWM60dWWm4Aq4o7RejQr5INzLosM+j
/rIzQ9gvJ5nxFzoK/9X5TzsSwUSJY1oSdvXBo40wLRAmQFoM8edjZcP7k6U+24Dy1G9M7YPE3hyL
hXZ7NeF6cvEc0m1rz5p63BDADf0PPGln9KkTInhIXA+uYpzctCoiHJkF/BW5kzuKpf4CX5GMGMM3
nAKcA4/4TejeOaIGq/3XBHXNVIw6d6ewz7isyLy1M/gilXRcaQycV2gSiaP0z4lUEatpm5F8kxTH
bM98HrNfH1JxM12Z5o0WoNgrk/s6rBViBYyQVRV2Tj5feUojJFfbmQYO6qElRlTBVaplSL3VCt9e
Z2ufLdX1WnUjQozs1B5uC+lDzlrv+8BJ+OxEt7v9VWSlq20U+1HhIpGXO4ixpeVwhIyRKESI9sRQ
4Ssb/uf9lrwxEv+5dMaSV3cAZXZD8RsB1CCrftueXsVXN/S4SanpPhKTgYY5H3iQ6pWJPiHnqfMG
55EaxKeWzXdKMQVhNKZ9u1fO6/rhuXcc+pdO0aMRFYqogFlpP20znMzApTjHOhe9bZNL+3W/+Wik
411fj1zBX4Wlnmam7qmg/BD1Adj3j1qw1KmojuxPtITTZwAD4PDGcbXJD29c6arYEUaYPy3EK/VY
Hms0Yz1uZO259Da+qnDBBnWkWBM8hOcA1JG57E07zrnXI45+he0ZOL39OM/LfoN3nEBI7KamYpIZ
Wo4eRBfW4uXqG/M7DBfz3/nB+NSdi/w+MUUBp6JzEWgH5m4aXQ8bixK4N2FrhZzO8VKhn0YV30eW
RIZsbeILV+W+USuP7Q1X2sePzToHj/okKCp9PiYOiNjNMGCvkq6jgAF+9NyDF69CnNmqijKnQzlM
9aaMKSimk1SiQ1XK5DQgC51fAwB/B5KqtGY/+w2mQZ5pYzeyL6rjVCxNQgBTLq262rvsHvhA3RwP
XsiVOZnE1hzujZEGhZ9fdBX/BOvtnCobct7uY+QLDU7sZNqXzJ1lxJfj2w/EHdhWtIfoit1th88X
2HEqCKIljSU4GkDSo5NurDKJ8tHkc6YxUBpTftUurhmQ3DS2DRMs2LrUqMhbAFmWknU3tpdtMqDU
EORs64Pa8dgz+g3H2NfurIzoiZFKgGcbgJzvvg8AUWzoy7yj0uepzWc2v0yhwqWO/RNUJ4SVeFgy
nX2KF+idGJHRc15D349o0n2lbrJ0QPvAXqbQQQHxM6PyWxmkK86+vL1GJToE+MF0jVVKJyY3t7Xf
9Jzv92TYEVLJIa/HtCTpKb8czuYPIK0UH+5h1kFkKU9pQ2J7ndcGFMT7k741loXJYNrGBI9yD9QL
H6ks65/XdSJuN8VRQO2moSih4/Gb5V4qQ7z+kzDQt1ggcbFFU4BrgA34toWScKycjcTo9/wT118h
rujbQLRXyVg8lrpyzslNLLuFyHaOBgeo8TZ3t0LuzPplzy9NbfbAUgslAwq5J5xQGqqXjjU6co6L
zXZ+pwEZTYQaioJDMkgw/R7UK5hkyG9RmCIV4vsii6qpY9FoFXlz2iXwRgrukZj1mDJFkP13/R/F
DlT4CRXN3a2jBrq/h2EkUEZNq1Us0seY4LdDWOpkTmzNKdXW86YkbJIVWVT1jnfrAlpfJq8seWKl
AUbJOetNwqsqgESkzzjWt1VS5D04e+cHe+fLX3o58stT17YNLw86YjFGod5croGJBJYr8zBJUKKZ
YwbEjSaTBTnomR2xaiACr3Kxkmpb3oOdT6F4xiA1VETfY3fo6Vw51/g70rwygCLJ7dCw+ZcriTbv
3T6EoUW/e9B8mZnFw3f3g7hGiJHulAYMocoRoh+qpY4fyZIgmUbICb68s5/LNAWTdO3rE8VQmScH
qHsCIgzVhdq1oUSlIcN2An/5PFnQOXXiG5EWwvPHUjTEqrmpiAtCo+nTut+n2zN8uRGZy2hLNnj6
idOXZMjljh6mUKDn5nZ0L1pDQeajONnPfhC3zO51Xd3gvzfGGug3qHSsh1BZpUQihJRQiMfAKO7W
V+IKv9mKDiOEJ/VcrQJQ8ulfBOHbFNYQSuUWDbJeaf6Zbi4Fd9cDZe1cx+8xkyXux6Ih8jYXuXXP
CAyvgaQ8RHTcxrxgw4Sr/hCGD17HLYmYJieb8qsNF9tIS+7PTPCoBbNO5frD49JtUUUDomCtQJQu
Y5hP2c53R6Krfqy67lZyS4p/FDd9bPR+AWr5E5xUb1oiC2fZribQbIPGHL0Ul9RTp6mZYdW1RlQ7
/K1ORsQmQbF2nen5mAlrDYNt8wZwb0ouTIS/vW0m8NonZp/ucVKDLfeeXU76REcHd6eCtzyyeK/8
emJWdPyduTANUVFIdTpkmOZE4v1H2hzK3Fkp0ZTAh/T+/wWvsGwLIygpNLBChFgilv28n3dmUUP7
ZCtr/5LDvkr82hZQs3ndJt0ocZTDp6W8xE1/OuYulzGoVDBA37VbymlWR7izE7P78N92hlWB79hi
078a34z7Dks94Nn6LWWqy+GJ2qZVaScnTgCLXs1y1uLNigBM6C+CDEA2MNR9zeyTqDgYNVWJonkg
X9uvmV7eBp6yn2icQVB7Ee4Q1n3zl4FULuBx2iXymiB8kOGWxh4Y2+lb7mVYL3kCbFhzyV8rj8Ex
9cFC41Ct13zMlcykVD+L4RBdkVIgGmjoyMLCv2pOtXljNAa1fjd2VI3k1ncY6ZxTGZG68h337Han
yiyx9lvMcnzNeeLPe5AxJb58Lt+lgYzY0kII97FQU8elrABrx2PbzJdelrxqQ+FQduLK+nP0KF+R
V3stIyLHb9SB2KBWvvXfrrHeofPkTfLa2GG16ZTZVSC+7e7V3k+IXMRtxkO1sIRNa3n6axlHR056
qGtU916LqwohzeJzZIRmKyA0UsN1Nalir+YpDMW0EzY8iLiemvLqYYA7SSx1XJ8fux5xerG2e9aU
sWpwIOEZRgAnL6Vsd4by4/+YRnOReFGRY6LTNNDRb3hQ4As+h9Ejiq0RZD8Q1iPYmgGIG0aQTzeh
JMziPWoElV36MJyto1V1oK8Tca1Vw4SueT1Oz7VylhfaWd7mh4QwWm+IcaSPeOmSoKaXPYNsT2eP
IybVEqlludP6phsSNh84tLQogS71iAk6YL13c9eOF+L8jlrkRRKVQ5MtcG+2bXhW4/7tkCUtXh6s
XDIX5w5iOcMCgfkTJlkoxud0tqFhtCLy26AdoI71qqPOZ6A25hAG6SOfA9omu63CaQDeCDqF7bVU
lmz+xZ/xLbDnani8Vev/1is3WUzDdT1B8p+xwzFuUooynfjjhOeV8XTayrfAdGLuL+uXCZeLI/mg
34pMUx4FVhj+HHYVTpQjrTPjN9dS+RNry02yC3SWAwqFls1lhqdEspfoUzpjaBnp9hU3E8rtkJqc
TDvHbEk9IOCrCm5u4+W0TSVOW9Ue/4LNhVtJhmHqOIHyzvPgAz2iU7kfhvQZIASArX1rQn6HV4Qp
/1+xDkQfXC4Dp2GNv9aPpL8+x0dmqTbvgaTIUhIkxrMpQ6bZy1W+JtU9Yo9m9Ri3mTqIEyH3gtTE
H0gOWPe/f3nayJwvPGrMio4ojJPm+uPeJoSfACX149aad90/2z1TeLO+Nu713Ct+zuyyTTJbC/kq
eVfbAYQyupS+WTs645Efyz0m16BDmJMcXYnULGM83JEEp9A1eQDmhFge0NA9B3NM4qytah4eguix
ttBDr2ndeEIeF2diKbLwzOz3KyEAVuS8gWzq1RfM33EKxNg8splUSE0JCXouMYgjX8j4V14Ge+/P
x9/tH6Om7V5hlsvrXTYvn2gUHwJ/geigsubJy9jl3V8TW6NdWNbAD/oIE1IJTRdyiSQnCbw2AvDV
+hquZjtJw5+6NN+ajl1H5/knAGycSXJIS8J9I6MZzTQbQkDaz15VNB4FATAt/oS/ZuklMzfNfYdz
YiafMxncEIsdjyvYxn5C01LUidpG8yioqhz7yZqAwCDgomNIR3gO5HWIDsUfEFL46X4UzxZ/cXMS
3brzsk2CMdH+r1AECV9AM1T3WA3akmU1VVzb9ka3KJ5QiM1Hwq2caBCzDom8xhvnMFUk94mIrgyr
2WheHSqTt+CMaYgWNOykJMkgfgrsh75ZIwLlGJVV647eUH7nrzd18tylnoYhy2Gu1DJQZmZmHqXD
0kENFhDKfrKsc4bP1jeV+U9pc5Q/bmj21OMmdGS5bCc/P/FlinPPyjGTePfAo5ZBGqlGQ0hMAHAQ
0rYQyMJIw8h5O6cWIzyKrCohprP/lU7hOPTazUczFQLxUv54KSQa2QAp8Z6JoPspj1jpqRAHl/oQ
QwXuRD5mjLh479DpmQ+Ll7Khu/Knw7hAatEEcBuUb7WiCAoEW++eEVUWdrEeGKZ9N97a98ZZ3nSi
NJhN9z5pO2uqJQEXxBxJ13QhvcdvJD8yfrHCStBscs3iT515pHZSNewxyfiSKi1Lx735klysHZzn
+7gg2Njz8SxZD3pOqK5ELihlaUr4qbFbgndgdua1w8xYn3TfPsznYuRuIl3F6NxTpzwxGcFCOn41
aQGC80XM99o5Emp3zWa3EuJWojYMvA2wbena726wUMEJ1dJMF9Bi8j8sDc0W8IYxwLEb5PGqk8+g
ygeSEBbOcTzk4HNkYBKFM3ZlfS5IpumGj2rTHPYd05Yi4YAd/2XcG2y6VokSkf79grVh3Vjge8O6
vHhYi08ypjgdUDHEy9me2q/B+1NggaB5eQkioiATZuqj3k4lbaxD07RIVHogtSlVIOt0S4uS3hc6
meIjwGHrOS6ujqu6Ah9vKT49penpQ7WSbKZjQnE+Z0NEao8p+P8MrcSJeaZkNkvWOruqzyohPU+1
mLiQaazfD9aRXxTCXjBeSajU1fKWLRd8AS+RvnHoc9reDedfQMw90+uyalQK6lGoA5oInUNnmYNu
ycFaBUdbBGifA3r+1UY/3zod/7gpbLYb4QhjfPt7cQV6kPXUqtjkibO/1DXujF8NaQ4B2ZqjGnK4
vM+14Ur69aOYK1ScYjmUwzgPvt2U/f5BrO8XovJihqC89vr/PM6BI2E/RrA7jedvTjWYjIHl7rkI
py2H8ifgvKucHINAGN3de8gnlaud5ZqKw+dLTJ+w5Ulne4n/S50djS56nH9RNXzguJrqNklh2wb4
N83PfNl4Bkoq7Bt6ToAOjbXz1VWOz6gSCC4M5fUGnGNXQQmhXO4oevXIF6OuXBBkUG+9DDB6gHgG
4973wBeIAf7UMSvUlzXQtPIWDVzU0MDgCzXFxVc+OAaphk36+yv+10KNjR4F+8goM0UWQcXp8WuK
ekWfOebvtFG6cO84CLw3VR9zRxHdHKgc/4B2EaAxsc+PiN58Detid0MglahOQ+8CcdTmG3DqnnTQ
SGgFhEjg/1QlXVw9Sxhs0GGiWLgqPnuEsmXBZ3zfV/rt95GvvYk5+fja1nAkYHlyce1QuF1kJXIM
grhptAYGawPahuGgTL0pIQiNT/5uRRfWM/D8W8/6T0wmQ3sGyZKseIXeqjP24ISfjTc/6cJaqSiI
P6J28bVqKyORDynYfu3N50VMSqMD6Ku8OHtGbOyATXMXiPdITeJXmjdzRGTXFYJOi4OmB8hAoGeO
yIN4LvjcV0FyAkpgTnnngWZFyWXTjmuFeFcCGY0GDj5pVz7V0WgotAr6Wz4bnfgFIrlIS+JS1NAq
yHK5Tb+6j4/MzqU0ml3CWpwuG1ZUcLqi3iVISl+bS5gnVBq6O0Bzc2rguFPKs1pNLyz+fr/SD7qD
IpUK67AUZi/Pbk8eTxQl9aJMTNz92FtX8yrbo+jnKI6jLzKqV9nB2El5uDa4fIc2R2d6jjwRY/vl
cGuSXmZtQYH6IyYU+8GB0Udu6vVM/jwE/kPtGU6kvKZoclzyqmKGCohkUrBwwkt74kWNpgkox8cL
KRt6S/T2ffQHyXF+V/X4jU0qF2f1KMJHhVYiccUcnmbZygSxB7hpPWmbXF5T4HC6QseeeZsqVIIF
HvDfpC+y6zlqFB7fZ56m4DtcSGluIzzKr0AmivhaqiTA2lq9eDlJ9TmDFk4fsGjSFcVMgoN+YGGL
kXGat8jyQKB7p63ZLINJi2Fi7JPB5KwmFT31CUTXEXEzWovLNVxa+FuWGMItHdKcVgh4G9HtamQY
L5MIUTgAGacU+18QiwpFsvZhUEGDKpf3J7F/zK3xM/EBA3r063tDfWyweCLA3R577r7a61dKr3ov
BbplqtlteV9Mq+KxzUlwyO5WCMnL1tIQAEsByze9T6VTDn7ElNWF60poU6yOY1tbNS0bMI7F9tFv
T0exrKQjT5cGzCDlFcsGM/eAXc4llOcdnrzoQytgdY3678gArcugOIdUb6gB7iF//BUm0Gw25BAe
pXbJZWV23O+8RRvZLywDfALuzoRXhqTCVQlZGaYbKX3h8rJqKshFTuVLtWrXezg92QmCAmNqM7R5
ziIVl6GcHSn6Uhrq/HEqscgfmlUxnQ1ZYy3Jw6NK2mHj9Ul78J4Ig2pUbhDM7pGSswcSa3CTldVu
63o45RMpXQ3SIVxxJ16iXrSDVM+npXe/zkmXLjEhzHfKuULRJPN55aE6Z6uOUwLILX7BpLCui4xu
XXprAd6vqVMUVPsdWgzc9zqq07kcrEMWRAGrqg5pZZXwri3xRD0V39XokyWrsv811Nh4QwIwIFHZ
8lgWj5N48nYTzHcIBOIOF/m3AgwNprGijwasrM2+kft+8BOVpy9X4vLuMij35sS/ORW01ffnMDuA
7OI9MKM3KEaITv6BD3lK9WXhyx3yFth5F8aROMWuJzptNKUmf3EkYI9oaAzYPV04CVRf9uQLox5h
Gh9dam+tDyZdzhMh1s/uKuOEK/LkG1F1mpDWJ3hObMc1MHAY4IXxoyBNoX5F5yOQ+XBZuKBwRANb
ArfvN0s7++q5XGYgUzpYVnMNC1IGxCmEt2tlYZYL3KkTZMNHOttBs6Z2V23k106bpMXIjWuK18cr
0gAyWqkDWS/lG3RhYc4PslPopn88LKatHMFN1lgy5tjCs4yD0o7NpnBPbtfa3YfKdY3u+2wy6Dd3
Tw8hzXJaKk4USObSCDPXTx4swNcVyJccliLOpeT8mvRVgOZXpgvj/1R1GSX09unHCtksKIAfuL7h
go2EnK1rKwKFFiWBt/xL+DgUtiMF5RcCL8LfxthdtC22q5jDPX3Sh+xXg9XddjuH1PZcyRE0R+31
sUykv7OSXoFthTmp17MosrU8aTo+y+L2lL+ybXlUlTKGJLV2LZLVTU+Ed22r3v122h8X/S30eoCu
cvXXkE5yDxsNiNtstPx73LVWPXCZEO0vjZ/vEkJY+DGoTUq1b9yxyzOluwzFgpTyBRn316vhRovE
0Aza3KVQzHXz0Ds7h7cKU1gTXOBpBUontOB5i+Sgj+pm21pSomhHoOftKGhrfQcc15nbzW4hJAmd
pTCI9U4Gzsdohn+ERR3Cl6AJVIfi4lj+bGCBVa4gmjN2j1aiY5ocYz2KjC/rd2RXLknKqNdhXqu6
vegpB+GYzp4aZ/VCkunlaWc2kxGq4yEePeXF4qVmTLlWqmZy0I0YD9OIaRwg1D30clVNPAOk/lcL
ceX/pn6XP8rronq+Xw340nPVlABwUFHm0Z+b2VoHCocmb1PDGt/NKtcyE5JB1X7I7+YgxWEspWOP
6wPKrc54MIYFigu5zL3QRK4v0dekMKBuzhAzOVgrlcHbyfvyZYnJlfVTxQ1j3BMOStBc+5QG7ktH
upZHIPxyN+6Eu99fJ1IaCF+/TQYPukBM/BQ8lY5QdJgsGYQ4KtKdoQpd4A7/qOUIypA9nwFCVwYC
jsNq2sYU644uI7npzB3gFOX9RK5FTBF4XGOLcJ0t9DJsIpTla2HfZsIMYlb/kWCIXE6dH5Srpd8z
028qPPYVyaYptWq19Hk2S2cud7Ye66/1wmn5v1oiRrA+eRAZYH4Fa2LyAb/3mHurDEwC65++Jd3C
a0w34oKECHTCX6Q6Vk4soB2g0xx4SyPZ2vl2w9w/0f8EkzSefvSSRuVxTJiI5yYETmDLvaxuJzBy
VxHpQp02GdZYr0+GMlZtfYBYinqan0OTTu+3d0/cDn5ksum4twGYEIsalK2VZVmG2/DPHQwubGGl
k2pZM95fosKK4RfSAo9JObvt8KFUjEj9iTTmj80htygttWyqZ/zVjXyLF3rWR0hEkaGyq8rLsyLp
M/u+gJp5chQxtBf3z6e9kgMfof5hpvzFeSbGbu480/9hhzLpJKsivyW8p3JbRcN9oJHAvQdOp1p1
zGHH0pwTYgQ3QdJPj22Eia4fDvMkFOhPdd0qmxx7aaDoFS0IBhkFAKJ5zu5i1OHJdWzgGcAV0Xib
h/XJicL6ReuOQVrfOeFHAuoBAztX8+qGrvXyzH8VE8SorEme5x/xA9nSgcM785eFtfjAbfxougIU
su1vnIpFRwL3KT2d9LQuY70gkOwV0UsuFBcMo3LK5KFId9phSwjcIT7C9PI6X5VYQbRd6BKUb4HJ
APRGaX1342Hbdi+Fh38IF9qXIxS75LAXfba9IBIe1xiscuUyVR9vHR948iub7s7oNhT7B04i/21B
TPAbIngh3fmHFo0XgD4y2gILwEyXgf+UmYJueg6g/rsgl9pYAnLniT4LRqjqQLPSfhbYEENoPONt
6h6oflnQO82f1YMQ/I9R+chgOcVAf1IndE4pcvKQjMr7cx9UMCmQNNbH2mDnfap7Yl/Fn4azd736
43GN+1jOZzkSoqSQAIybvWpoQa/kb8nZr8q6F+t6y+HQiOvg464JIM1NyhV5/WkVDMTmdLJ2wHom
2uUeEx6oirwj5/imLdk+9Lk2kKpNlqLeXgaIxPB/dZBs3MuEMf6W5xwW7aZ31Cscplpk8USdWx9+
+hkLUdSYru+B5Lsl+jAynecRJI8Y1xA8X//BCRu5qhOBPmAWyxYaG5ETUupQ1OsXsbPLhFX7ZBUu
KGowNtPdCJO+kH8cIR8zyLFQUscqDOtcfJZkfTxksMm1dB5Amq/9NqaSMnNCOoSc6M0N66QQL8a9
0ozFxMQEvc566G5RUX3hlaVJRK/WvXbNvbBYX1dmzERRlJHwOdCkR6XKiBYsJGqiH80873PiWHu9
BrgaLM0jqsPlWLMTMRIg6wfq7CAccgyndmkRem58saXT/tBZASuNTgWKyrpCNzbrH8vZ11FT0N/K
3S6PqSH5EPujP1RuqgSKk9TuWu9sCtwPXxqpk18WAhzyw7x7/MYYsUGMk+rf9rGdxdcGw/Nr0+VQ
AKlxFnjJlSQFd13KiH5g3CCfZ935cdbwM7DGi4Jkmb1O6Z8f+pGd87nAKBtM03GM+zFC5C9OfqfD
TktNEZRYpnBZi+MrCpcVAt+Uu2pS1TxzPmpnluwlf9SrqpkQJwaNCTgzdUnqwPz9YEe/sWSTWRkw
Xzi4VQN6ZxGPEElu67sDqrHXfUq0lCsFsAL4axNXIiB6qf6fYWAA7Rpd1di5T3B8tl5Y6P3oAT5T
cwP8BlTNI7/OAldmwLWztLlq7pWFVPdiHiYBHBEGnmD2cVH3qbBTOqEm4X84qKJnoQmjoPc3zOE2
7vRjJn75vaPyY26LKMmQGrg7mEGw5NING2C6OpsHQEOn2QNYEACCYxpmBnnsQ1XjNgTAPHAbMS0L
cWIBdyQpGhfptwA6G0ii4R1mMvFD63jLDisyDJjKsT4pj0C0Z4TOwl29DgvSX46Y7DaNj1QyN2yn
+Au0joDgRL0HRzLcfRTDaUIRzEKiz4KTeglYoa31vOE098x659NHEQV8z798iDMxD5juyJcdqdjr
+eUaeE1Q5Jcut/8btVrRYU+Oo5yiPOK/7uUVBsTpirswa20ISXBT2Ca4ApHsZksm8y4zXw18kSrT
OYE3RDNi4puJP30seFmkTZNPRaYRA/2mo7Ef0GPSZi6SV87zcHWwDP9zubC8v7CWwBct03f6WmM9
UHqcqmx4ZGQQLcP1NtWW2tJCxTlXVrayerLTDFul8EM6HFnnwzvpuqhWa84KKla7Qny07Ug99olI
SbPHiLZ21dISjei9w8mJPmu8KX4MTziBE0k3XkYrr/qjlJoQdh2v+sUHrR53ASo+tla3KW2WFXi9
IB5oAfmUJDd1VmFw32TXWEFaVe14mfPzg2cD96BEaSxD6GpRX3wSC2dfzoesml2Js3zIa40PV53/
nATKyR1XMS0BeOx/qWfmuJMvJd+bnkmPuJQREmS9m1lE3hfQs4RK7N6IUCn0XRbO4LiNuVypuQW5
ZWdgGs//KYESTZRaNNeUh1ktXkGLIFNPS91by6jGnqhsg1APvZVfUd+VMaOU++rMiSp06mdzvt+o
AoMI+z4lh44dhw0arcUAL4HssMK1cRdZLBlSgw51LrtP55e43xzR7gsZiFdHzddy4xUsBhScXBYJ
J8W22hIlPEkAdR0FCxWfyprunCzEHBw5V4js2YUkbfn/tbge8PIPUHxFG46VRAYwNdsQtqz11TTg
6H8OkUvvEqdq29tGpvMzW0kbUnx4SgNdgOpKD85UOainCLa5dZjKTz5GdEheisT3haNfoMnvZ+Sf
IXTbGlNP+kz0af96JpijCVCOy9rU3J67hvzioZFD1Wegs8najhVEHNlvLLWvgeGsB3fgndVtOVI0
m3d0MNHwzIdoTPIrCGb0HdpJjHzzZSVV2nEDGwphNW5Nbgl4WLuyLpX907PgQrLe4mtFa0AtWk+Y
gYukoQw3i35idiD4pTyNNxAWT3vxQ94vmxbXxSbDB7l5QrlwwWujyWSEW4UBdIzYDfSw5zzzMO7r
dYxy+ZlSVI/JrYe+9cOK/0SAdeA1yreK4lBZ5/F2Efs8N9p2fQugTvl03Ew2CQtPwh/f5HRE22If
107KbDZY/uZe0BFUeEmNPV4YMZvidJMkBdNM2lh56222+4/RN7ZZeELbQaZuLcOh3JLEk+2xmciN
LSBP9L7KUojIgSzqqtjlVU6X7DK7krT5yMXrBD+37S35hTg5E6IzYC6jXxhN2zIElekqW9ujX4hJ
+D57ymiqvAlIvELz64sdPfdjPDMrDXlZ1W0LAwEVNsnWxX3QdYXMtcme+F3aJMsI2rRwatzrSjn4
c+RM81CK0maCUxc0MXFYu4xYydzXaeCATWPO8ztPED7SRgElMCJEjf/5KEsXf03FRgyGVWjKoKmP
oi4MfyEH0lHDqBiWSfVdvt/ejcMTdH94sdmWbnicUhXNfHFbZi4l/SaeT0ZHwEPvGRs8Ek98pz27
40PQHG6SNlwGtspB5OM9nonIuDp6ersUTUjUtMh5GhfvRBGukif3fqz7p6jkPNBHvTT2WifAKv1z
Pry7N+t3HTX45SqsNiKWm9RWtkQ7Pgzr8MqRIDHfWE+i8nYXn5+dJ43QTk9esZuLKvcI09rBJ//s
u21kVgK0Pt83mEG//rWiWzRPG3NfltMSe7Lv2wCv9IosAOMW41qw19WUheJnCZmE75atSPS5dOju
2KrqClZ0VR2X554RwjwgijByl9+f+/az6wzJqRYYG+5R9ow9kLLANxWznTJBoEFiQC0uDPyFLDOC
29GLLlfzi6kWXZVVcCg91w1bTVJTLbNWhcoVsgb0WdjLv7n/4jql676vb6LcijQYrgVquJxN/jsi
/tAIE2w9BcitTVH8V6PeqKAGHTjkY7xgxfsvpZKS59bty6gSE2KT+zg2CHZ0pR2MFkgoMl6SOCxc
PYkDhIv4bN4dgDql+sxYChWukO+FZS5lnMjnVOKhWfB2St1WBMIABao3A58hxrOboPXlSSgihR88
WzXSVhB49Mz3HbxmqE8JDWy7YLP2SzL3V4PA3iyYfZ7V2Eqe3ZVrZV0sIFe3F4vD5T3Qb0CBpkPS
dQyvnzhVIqyAaZJqJhHIeUDwtN9+NX1FwmX5hwXXC2VEWE4hhSMr1YZuxAZnmpRCMSR6qdk5dRv8
eeWg4K/8do00RI9yREbBR4fih2500GhO/zFpLko2vL0Gqck/ouoxY6r9MAkFlMxH/cQ6cHINHD6m
sQSGw8WMtn3XoSf3zKRBJV+fRTlgRR+NyvIyAvy8hl4t2M/WV51xoVQz2qbTAuwt1RPAvlwTt0zd
6atBfmZ06jGbgPLdXEJaDzZaD+sKPfe/ZeWj7nkYA1GXmhACoH4+pVVeiEt+sEQvXmWk5EzBun/L
c6N3GnrY9yyXKf46weWIo6v6JTvenAYTa6ekftHVh8ahfKeqdEo/abxRswd57IZ2lhFjq19ePy5T
PPRZoU19aery+HvbnRwJcgBFjpNMcPSBUlTucUGcSqrpgI2406mBXlrH/JBgSz6qsPj6ZelUabbC
VonNjWnkCOCJbdTBm9MdrwgT6RBTCkC94VGfAOP7eap+HnQygBNffCWxFklndydrYt0KOmXFPeB3
oCbrf17BImHkCqAF/W20sBl5YCQ60tv4lR/Rbt4XtEzg8DKjcWfUU3ZSNA8ns91AzCjROIBOWgw2
gd0reiBlkGIVKT18O+fz4SCtjYeCdVG9pQnnJCi4GxbhPwzWLQ4dTgpqOTHrlZ8DXAqkd80ni7/B
5iCRMwM576tcJ61daW2SuWi0yjhCNC5WitMObUj3fFU39UZh9DkTAYe7bh8+dCTIV55Y0LVvDXEw
gu76Sg4daMqFHCaSmFdCGToq+0JWrhgNh2wbe/xqjbhojIt0UNdxiNtCCNnfcrNj+UvFB3cGHg2Y
Y7Ng4qeAIc1Hj3vnPl+QoJldjAM0ojkJMe/ETyd/gyP+/T4SM+zhqEIN495dcPRc9WARpnb8RVzf
RV4EE4Z3N/CQheiZnQqFZ0ZZ29wAcGlYdGpTd/AiPDkrGMUfW8MpOhcIVMF5Vq3mpsIwaIkmYbZM
/326B5qEbZ6P+0UbYH12HSnNEu4i/MnPeOsomsqQCCizCkDdejRXV3JU2CXqS83w5RFhhIyuMS4B
Rx1BEVPYxCiqSMU/OW1Z6VWUkpSCm1GIIL/3wganuxtd44VGX8SzIGvbZ2Hulg+Mgu2/ItH278jc
OI/H6CV+sZ1nZcC9t3KGrc926nmgTNHGYwSgCYXXqFjtQij/P43wcbmeZ6YEtVVNjE3pNm6bXg7k
6XchHrU+OkZKnhIV7uw8GehpoG+3i/ajwCW4TxsiW2wcuSbt/cpQsX776hHIA7TzXj1SLbO/iTY3
J6r4igPgaMHrCMOUL8iijUdRQ28au2qpkc/Gq6cL9mGNn0s2Si1+S3+1p2RRZxY/IuuNRDiBaJ9b
1UGjJcuRH92zbJtDlDEKuee0D+dxfAWDysBAVRgHQyYNtg9ZbHbGTLs18RZdZ44ggv78XOUr3BwO
PnsvMJjq4DTEvn3vE9B/sGrg7ER+FNQx1UimUkOEvNAM17QdMZVhOZlOSfrPam2mDkuQULj7gd0T
EJ0Ld2CwKT23zyXb32lZ/h0tAglj3474E6S2jr9p0HmMGtJkLYnVuxsZSWp1ZnJHOh//+fmgpG3e
/8yiwMJGc+USraxglDitPdNU0qX4TVHPs4stTkoRiZ1tuCLlQQ9p8GHHiqU7GR6xUetsEtbOuaSS
3evAQx0f5JvhBrGGzcInuMvIcYOnlWXbF0GUXfeEXaYMujemsyhjpgShUBxZZdaYUbrF2gAlk4S5
XXL2cNW0k18H0OG6X/82cG3nfDE+jsHyHpwfwXmh7PNsqLYXbjQvxXUoPvnoJ4CJV6PKFSqMKTW6
sHafhEO4CFrd+Yc5GuEjbqvSHMq9BRnfs4oDJqpOZFHu2j16lWdlT+VQFdxVT/Dil3ZCvQAGHp0g
7xxQzomU8UtIrE+u4DGdDGNjQPT/+YaiskndBd6ahIiBPnvjkqaegSaAjFK3m5bm9Y4bYFmrr7BV
RVWx1Yts5C8azU+rRtNzrAoWR4OCns6eIkF6TGsJ5sa92Cq+qwDL/8DiZ/cDznRcNnahkjl/LMEd
V6GXUCYti3MOTEQ3NY+O/UYD2797UM2o+m57VSXn/h1xG0MXmAn3G6Nq/HOGYUArrN0JqZzBbJm7
8k8m+/A1C758MFoh1Ps0/kzGnBD3eP8oSJ+b06KziK83QE13VxAP+QKjlEqZj4ol2ASaqxPTsh3r
hoVLWA25mxRAigmz2z8A4xbet7FC8MOMBX779svONw2Zs+IQ5Mc/I0xmhgQZ7KSJ6UBftYQPjD9U
koL3m97HCEBjHNTOc4dH7SyU37+/914NbWRuZNouKPueWjGCGml6a3JJpcIsNeItBYk9fDQ6O5ea
znZbgu0WT8/GL1f060LZGDe4a4LU4Wg6zOoYA+afGap5JfTAmUId/t8TufHNvMAFQTEPhrlNIRJ+
7EQQf5lvnGHaWWDentg679nxAt/5hOMr/ukDWrELEpiaI3vWi1MJIZ2F+wxzIM67Ht1EL2oFWe5G
FDw28w/vcWcOrCR2FkTngwLtkW2Y6G7eMr5sISVvuoTFL60Hti0ZRbCf0N4R0m1lXRVHbRBe6dCH
muTiWInSgXlKymDzb7d0LmiqK49hEjaF1DBPchr9zld3aBpmw707TTldhF1ATb3bBjpxrfXx+2EP
zYbSdvfkDRtdfFsxy0HenwM1IGh7hpj5dzcWWjTU9FvsMViEZLfZYrSj+54/+hIc7J0WnnWrzwwg
GZ7aNF9LO7ABkDOt956vaBzBj8sRgX63AEk4BYjN/aj9W0pPZ7w8xnUmHLAcL4azAWLSoXTfQ4Pv
Suh3f1Erh6iE9t6Yun/Pg382NynNUNUIe3TaX+wuUPfAax6r51fbu1ZnMtlc7Z6a1Vpq+Uc72I2T
4hD5ytSWhblZ2ppz1yGxrxqfpgNTdPwhD56kD+up8dngKv5qcxsodWRtFFidkkcNJ/qG1RtUB+vw
H1jfh3tHqPSPDB7LqY7+r1ZFp1RF8rCxpeQAi6qN2+JldvbIEqgJEV9hZIRhzQ3iJQXdWSns9Nsn
D9aVRjAx2n9KRNEEbOGT5bRJBdRt6YHQ4TvneakFi7zzrp2ka/xByEatj0eaCZWn3+vWGxVvhPbG
Rrg6abrVQBs6G+b4gb0cbYs+6q1QtKRfDHv1MHPeXwoHmwJlLv7hlKGuKdJ6171uVV3c1aTInuFQ
9pBdoYLsvrG00voj+sMakfIzu51PDg5VDORU6cTGOH9IecVjeUrLysBDeUg41roqZTBIr7pbCofc
4AuHC90h4oGikelpB4RNwLhowtW/CxRX7rxQYBNwXC75nvObj/BLm7gOjV/aZR4nVR9hUcl796kK
RMznpjn0OVR7hLKpWowvKEGLbFTi42EisKy/sefCaLFCeQZr3sgwWpnSAmNiBgaD8TUMLbuD1+im
05SmRrfrqU3PQkeI3oEiHLq6brAE/NNLeERSjsJlsDiM/8ocho+EYvIHNubXTNZHqmsPNokx6H9S
a20YyiIxKPu/e3XD9qxE7+j6tL7BgKuFXPR9kzjEKbf7Z6JYFLYuLnfBNSdn4MzzcbBiZ7SxCAF2
zwY4Nt8STRzVtI7b6YVeRBVPFvxf9r8o0PZW7ay5z40Nk/dIclJsirZQwxq5yj9VRF/Br2Zo7ZJF
Gg1hL9af1l7/fLmXGDOjyuKR8t/lhsw2iZ3gHcp3MTmqNQsRuOnY5MEL0xLsGHsB3s9+a4N5x3a6
mxyZP9kPNPFpttbYHiXCgeyCZGM8yu7HSq3A5gcEQZpgHi93+xwHdmBWlXTEHTiidFkMTeqrPSkC
lWKHhpBk6qfpfxxWkLSdGJqKZd1/2NuLNbOLDP5vC/IUwScU8wfrW1jc+v+28a8w5lPf3lL7rOds
3kcZtRJDj5WVD8Kdt17vjuQAK47vYWpLYvJ47Ednuwx57h70qK3oOu+2bOTzCb2xcx4Ljw+xRm7n
ZRb5K2BXCbxCDBtwHA9Np1y7/wdA2wYN+c0wiF1szwVOfUn8Oi/wVqCK3CupgIB/Nv1CbIlCcrY4
6HIAFBDVJ6ArsPqc52y8J3oGHvmmy/QilNsaLJhjvbw3oqr45Nk+DZCVEwnetwDX4OiFMZSMcajW
SgzmX80nyxmuVoxy7d0Uhd7/zCogRri3HSpxd9WoZnHpRzlg5d9Rofk4334Ae9ERtiZIB7PaAEOw
QUbS5utFNxoPk2ybGxgLOsvPT9fC4GKzz291by8Bh7saFPvi0tVeEGIekY9gNYgErOJAMRKKzsNf
P7F8oiDWIO0jxNfgq4zSZuUdExlo3RfnjqjrjRI/0Xv6YmmDrO8rieR5394vt80gaCXCcm0cuvUl
0LpdDS+X/TRBcNQECN9DigJeEzse0jW/oS6/NMAXNe9XttGlyGkzYLYEHbo6QGhqCvVNtnmsE9U7
HPRuAHD7Cdwf3K0NsRLyXijA3wy/uum+hCfXWqX/BCng2nMNJDdc+zrknvUiIGkEgqM0eadeaYDq
ukjKw2+qpJhr88QbGAzUh7Jkdg46Qxm2iYT7WTEboJVt/0usywS23Ez8i6EMKQxw2W+0Z6758+YB
xg+LEU7+P9RD/v2BQGYScKcrM8lBdOyVRs9dFMjaYARamj2I5RrQ2q9hhqzgW0u5SlnQRAqLjnUp
Vlo4v6+7vQ4KHQAy+RVCV8hEKNXXCp7Z+WeMUJbEBl2pSJeyg2BMyrIONY6IyJu7COj8hwtyowJL
cSdYAN7WPKpZiDzBpus3TjqwxMCof7P/oymn5JHW8HVwO23TBcEZJI6djS2Q2qWbDUd6ibSO1Bqz
F3KNE/+Dr8DBLML3JCQiwgMMFYAegzX6NmFm6bgYNKRNK0pVWnbIB6aN/0wuCC5tVkcJ7JoYbzQf
oAB7J5InoMFCpACNcjTrLLQav4r63hFmo+owDZjm8J79tj3c+i3txolwCWus+Hzddw3/BzC7cycr
C7GfkKcEoHeUMGw9jZUn0PqhzSwuOvJxHwgZuJkY0yqz0nhsw7aPGTtIjA2YUmNGY7f7wbr0Nqwn
yAqo9IGWr81p+Xd3MXva4ynnpRqdk7RzVqU5NEhzvkJ9RHGya3iDK7yboQ5wMfI3SgzBJd9bDjxt
y/CqTNRTovRS58884tzDTheBmVpFkQbf51Q1J8WbuBVaeBp9KkJ5/9sIBDLuVmU8D/vxV7k1bAoJ
Ywa5aCphGnvQTCZQNtvzVDzOQEPZD7GiRshmGRzrKkLZEWCmYq/8SAgqdLK1YJ0x0BpsDaKG+FtC
oEy0qVVLbgpMM8PqwBoT8A8DHXS4A0oxMtLAAwolIGXflAU0v+L8Z7T6EfZej6kZMvamTCbjTaKT
2UwawpRB3KA/HmHwYYkuNxcptH0RUXxkiY9gd5r6CZs3jKktaWgSyZQweeYCIPrAI4qjHS4zETUO
F+xrGR55nGcFRwbHqSFw+NE5vpY2k20CgNhGLEOJrRAkfIILyQ9w5LPZzt3dBZvCFjSpP6hHAcMF
cJk3phyh3tBCQq9ILU+W/QfjpZzhs2+ExTGXOqOAIWAs549zLwVKyWyoTCVZwWdjhkVgpV/iqhIR
5moG+HtwKL13F8xRoBSb4lyoc7ffq5aTVkAOIFRu7AE/Zf1LuzqOG7yKFbo+DUOYyqISQ/jPTIq6
/FibYJryeH5ld7g4CfS2U8B0Vc3wMU4Y3/wGk3z2jQtFntDUUMx9oOQkywDCM5T3zW3wleRFA8Ar
OZokS85UZEmd5f/XBw6t6a0JxjRh7Pl0c0QMIyIG3Zdg6nvZnKBAxpcP25j065M0vryyqr17o8pP
u6EYJLX7aEnegr8ZjvwUQIYMr8nYLTLqqv0rvMzw0nxQZGCg4hvvG8tkXw+N1muK2dw+4xWqogxD
xIhsEDuQcjtN3XkafA1pdxJMw3Zma5BZ0C/sb7wjZzxSOEPJEWnrKGAcjXzMwK4n6DbyZUUDqLD0
y7H41v4BAMLYSFpo9XM8AmqhNCktR1nQU7Dotx0Mhj5REhyHcEJnBdkHsfUWt+KIZPKhqjWrLV/H
NrUMBElDponIN22ekfLmC7Fx9az6qkeQO1EXVEZzCPZ9hszADztm+CzOsx3hcg15LQQ8EkJC/kJa
/kEKZ6LM/QUksNxmDcqjZGNxC/jTxzptFjnTyz1BbF/ETPnwaX5rg8tVTNp7fIFDiBLpN16q27lG
b+RWulmr29QllJ/pGmSakeQR6jmROKMSKYgHv/2+yDEmHle+gPOAaE0tZw+2zB9zGhTFLBzpCWYj
dWSDtVwpk1eCSat+NkXxjjjvhhAIasjJVN0P75dyQ5BPOCuMQF5Divwc5mMMIlifo6ezL9R53aWm
ML2NX8bU2yGgg4mgJUs6DIPIufbL1B2A9R1eMi0GaqEarwhpr/pMEjAbPmN8cxDDgkTyWzQO56nv
8J7XKRjT7oyy0qKkJSbihA1P8soRREiwoWJKP51c0ijOJOJbkIh9bqxm+rkuXDQXmpWM3Psso/n3
9/UxXLphFM4wx8eOC6vnk5iTegJ5R67r7O7aZI3xJeUMYiQGbctMWGoA3dxoYVXqyQjdg/QGiQIG
TWZ53z0kRbNJ/BpnYYyoF4RdMwFpwdhI5zMgVT0ZLoKvJAYaTD+FIGA8dAb/AhLYW8tmY0CB65qI
QAgE3G3wxdUXuNA3YcoLEwAEJuEhzt63tsyeHtBkkEy9Zu2MhLH6LqTpaAGpClD15JXWkqHK2HcF
90q6vzxwy9qQxoopoCOBNY0/5KpXQhl/+zFp854AiFM7IDeWD7DSxoi/NkAVAAjpd4zNy4lhL+i/
IIQNZp+WPk/iWun/JjFMR7Q8AIRJGuLV2hJeGwdnvYEXw0uH8HNqD60LngECpRCa55kpEk6bdrAv
/G+soaMKTp0MN00iLID+t81Uf97SlJIRARM2LC36qc9IK06t5640TUhQ0Vh1rolxOw9bG2yBczC7
ayyIu04JRtlr8XxsMetMMNNqOSLNKrU0vZ6GvmZtW33ZphpAPyoNnjcg+v7jyt4NG2f6IiR3ggc4
84TRLcDSgYw5Kzqjk4VYvDRc5xpGEysUp6S9RjOKBU/4RyVTt55xdA+Nh4XikHdepRQbF2kd+qDF
+GLXBd3z33lbahd31dhk1SQetoizqTZwrivAwoV5zqW38nPhSO7Tsk1eD+Y3dkd49jhfIoXpLgjU
tnSr3ht8RM3bjB2BkiL9Y4iYRYG7w0PXA3kajkFFLzDxL2/kshy9+5NBjibs8rnYwa5DX4nJOqgt
DQNuOz/UM1wH/vhvKYBaIJadr+PPBV2tzuMCri8GqZJ8UUQNJTZswOAv195lLmPCsIoOH5Dh7srW
D9QcG9q0Wvw5vDr33gM0hFQzoI8DxQSOVt4ex8eyYq+afGsE317754h7lBYkmhwviNIzg78uJJY2
JGwpKMRsTatZrp51LTlYoM79EsxG7u/pZURzGHRWdjouPnCG0Sr6ezrQWVBV8pAVHtbDXNzRDxht
3RSxlr+O09VbopyP0G17NtLkZf/DkqlsEleWrLe5P1nm+Qv6vxLdqXKbqTo648F7MwpKno5i6rD1
RzPl6STZhQ7VxD8blIKSseeXP1ddiJuL/c0EZJsRrj8xAOHkaSe7k3SXSwDtJLrHvFzJdv+/E/ms
FEAwMv/BWs2+bbSKKkl5lam/axaLmKP/SIejaO3CvAuE457am6CCYwKhb59V+NbMiIry01RwvdBq
D/12fEa/cjjTaiPSaOj2BKgk/IM+WzmrID7D65PB0U9KZlDhpZYYaAR9HNobv0MZ8Ufb3JgHTq76
4zPQRHG69JiBuwr6nSmIFD/XaJd7Bw0bUAZqYFj/2tqLSwgX1qGSxvLVRIkJcOBPoaz62GwQ7N+m
1lr8Be4YOdq1rVq+tRogqpMcoUvRnkwXKH/HrO1lDsVlTVNVuZAnnpq9ZrfBIF0XRERshoELSQ1v
Wn5BwLUIPKk+RLDXnrVurVg0QNhzCc/xY/G8r+LcmQ7ZPhmK69A6edOS2orpJNYdjN7afct6lXUm
xhYNhTck3a8mAstmnr5pBLPpdjEO9xuQphUkFTaImtWe+BA9JCOu+nlYPQWXVguWv0NwHCbjnGq1
H3MNQghYEmBClWT9ebxdW9+N3JPGjbeAnihTqHXSCws6QVf+qddpLYZzLRXqmMBPFysdVm63XUXm
X2XUTOkChlyyK0rHD8XHgmsq7uG2ZgBOj9O/ZK0TYS6Gmg9yNiRwocpQhiy+jMeZvVjVSjVWuDQ+
K2j0QfHZ9a8WGmbpy5vSW0aeYPlb8U5lerC52smi1tKlwUDx6i52dcbpt8dntGl3YTmJK5YIBnQr
fWY47O5WNMKhYmIDR2odsF5mx9Gi6pxVtxTLSjKeo+yqy9H+X3xK9IJM/jwgC/g1B0jSbixKfQM8
KMuaG6Y21locHZW84s10pfshINAiElirpJ4D0sac5R9OeGITonC8elyt3PR9hsRlzfdIPpJEOXLT
3JprpjI7IQdGmUIIBNkJFi++RhUOmLz0orq5VCpl2NmhMSrjjXScxFXM5dpap7WgkKff0MiUaJh7
wlGBil27UEEzxZDlsv7n3bwL3Ubta0NyoGYKFTalhtfzy87T0AFSETtfHD9jK0Hy8b+xnnkNCZiz
hVkACPSGVKLc7/kjDeSxR0LtrAGqba+eRkBNYaifELOYIU+KN29Bi7o9oTW87Yw+XXI7fvO+I1+R
y5yPdlfmRjkTFPXw+KQh1cx5/nyRKuoINWN0mgyAYVGgM/9WE07IVESCZkXVFyx4Cndpl4O3QBMV
iRgKijC7KnQza2glmXJN2WLjWOkxnSM/Y+KXNin0tBYk07RtDgK8QMibL0fDUls/bi/ReDXM1vwW
zLUttuD0DqY/z1QpA7yiqCdZA9JvMwwqx0Xgq1BFJHiCgEZYNz3mC25S6q7hkV2q/FcP4g1KtF0p
PzE4Mo023yMd1mZ0xFP2eB+/g898Z8XjzSRnQch+pUsRKDhKviZ8lIFlTtXt6/GH9+jkArVYxkoj
Ev0ZnFJEws2eykeA+VVimt5iS/J4/qQeREneumFZuLMRHqy3pdBxN24T+4UbZkWu32B6cv9rsGJL
tces/nkmgcjO1kZ9AZHhfids3VF0s6C6xOoMyJUfph3AoLzA1xHwe8oxa0sobETlz2OCsuB/tqNE
WOZp0Elvpu3tXALcMQIYuyg1DBhgCsAxuBH8RfmWADXvTL4dTwXDNQM+5jlMyWiUlCvmkekdb4vx
yo5Ai//sZquUAB4BkvL0IelN166kE+7HBGjd8q5HESVRI5RkWHC4YZL46+9scIK7T/+80Cz11Rjy
x6okUtlawEWHHFv0+YqT+KU+d6qNghWqrVf7E0Aq9xI1S8hEhVPXUwvDU91B7vHn8Rv3MASeJoOe
DXurQGgR6zO4XmiSXs7V1qlRkE8TF2bolx2afxN1BcXR3bN4NNW6JWvM4plDemF8TSxfFv+VyXAq
3WUbWkttO4j/Y9OmJKuYZ2ToKWB2hFED5UKd7MQMTqUSkE0RmP518J6Zd2JmgA4AKMo9Ds/lQY5R
i0K3ma7EGBjq7SeuZiM8vsH9+FVDxzhTvSI7CdiSLmGJjhMVE2s7y1aXEEdeaQKaPvqATIdFwOI+
OUUZX14/hDcN7yOyNLC39wGxjuOVRIuse+JL4ocaP7jO0DNGYU22Pi6rT3ODgeZEc2yojRP2boxO
ffZZp29yYyU5bTyK7IIMZpOsQujVYuvGf2mP/+ajrKJ9p/3ixz23ogfNskIj3u3qlmhA0OU04HPI
dtXP9OfSrxCwTdcj1D2lSRlpNd4aNTk1bUGkdg0Yok50b2xhYEUSboCHF9CW9iHaB+jEEAyQJ2Ll
XzF5rOw6V4SrXmu0OYZGDR/q/2dTZkDIdtR54PWDDnduP669T7//svfHd6UuQah+8bBLF8jqPVL1
5ZER342RNdg0tq8ndH403sRvLABAOgohXyMEg6IdZwshg5PPSEB7DxOrpeXXHgyJdQmScIOQOjTx
F2y5wVuYq7pKkiEokpRAmgYcfYklpZr7Z1KpUTgepmlaq3iufBaNQVk71NomNbeDO8MQdV6pUDrT
gbyXqC3DTJ2D3Jt/eL4IPi5HWe+aRo26B8geTGYkH+4nvDhsRYTGfUHWeW3o7u2HnvxwR8jF1wcr
Rt/K0YDDV1M/bwoLD2cqwkItXkNQvxe4iDRCBSzUVDnLCq0t/sexG0Tkt5zM0G6MszMoamlygkak
v9cuwUMqpjzfHcHgpECgjIK9NdoTEGHsyuDqeqyoWZw4emOk75dJRDqi50i77+Ltvo8R6FxZxCwj
X0BnfkcqomgexeTBM2vS5BiE+BFU/KoLpGmc+6j7I726gk7ZvNVh+8H8JJAnSXCxopI0QSiEGx1I
2zcc30eA3Veq4axosrmHXFZY7CztEV/rTVtxnymVQc8xLVquZM4C9G3vIOz1E7CygwwGqmDX5cY7
eHvKY5pvzr7NTCmVqDjZIQ9zGj/nZh/PZW/cKqcVgR2z/onIdab13+w51ViE+LnZZgKH5NVh0w4/
+zhgw7AyJ2O2k64Rsi+W9NchWNC6saXtjBYrsVSEWSkm6SR2/Ezchiv9hsqJnoUjkKpMDYA4Ce2t
5h8RrKcXODOHBYQQF6CGr2iSR5slTKwBnjhpar51Pc6yhq3OwrvNOxlIdwy9/EZvGJtxTgUfRX/R
z0OYinlDX+Pu5QqFuh8EX13tkiQMutDGbsknU4328pGly2d/OYAtqyNI3Sg41JxSVvQyqMWingl1
ZyQij8ZJfDIkTwUWKvTMBjZ2o2UbfE4jOGA+KyRVT8nYSx45qpfJyIewiBloeHucRpB3YP/cYu/l
tqA9dVqpK4N6dUqYWAlNnNTyUzJb4tU7XY4hoPU4w4+/EfzjvXvrah9eCXwoWrfCV6rNNELWWtiA
RaFG7xPVC9e+gfpp2iRIyPmR0nTJWOckAaW3yb84QY51gPOVMJdADDVLBOGhq1ElNS9dv8Wd3in+
w0xI8pKuUE88L5t3axqU4qc3Il1zRVHiIG2nsEVvandbisryNnDsfpHOhTwXXYWA/loJRt5nfKG8
KdNvluSPYStvubFPC73YZMgm6Q3Se3D9uxv5PNI2XvkXplLFGPAOmBhZBWEyNtSQ4HcFybqQLtwG
GlyHfegxm2UKDWcJXt2I9/RrubcLqz6EGn5soBdNRHBAs9K1y8sPM6yL5TtE85/JKzQr82gWjx/A
7gRlvRO2C6Zzm5UwRa5sitliIEziCFsbG+NG0hu+g7isnZ3od5Rx7KlbFhai53At1Roh4kwtHIur
6mx4aetrKkVDZMJ++LU0BSQEfLBefgduI50BTB0bvrxgTffCH3+0fAnpa3HZJDdIRUNa7RSL0ni0
1/9V2iLNhUF9i3I63fEFMc5AuSEZn4tNiYcA+hzg4OPC9SPISrRX6wsOwkqlRWyMwGEfVGpfUVsW
RyJDIa9dMKHL1sAH6Uo9IrtLQdc78w9CwESHpgFLsi5dM4JVMIOZMTo/jNR4r9eEB3c2Rw/6u2mw
j/tjQkrhRusHx1puftvB7mKftqE0PHVE/kmk8mPZkx0L+kD6beXxlqL+ohoOsorwvWl6PGiov+lu
Pl1I6YbhMMF/7kuZYsGmM3GMDml6ANpdqsVmD9p4yXn3HlSSgH7K2MlvauWZ17LcwJ+adlivzGVC
0iuAoWfXiQaGPm/4i2tYnEBfmMIqqY5JGCIMUp6DLCDODCoKFsc83VGlKxVTUHiLey0UzBo2I7df
XDDRkySrQh1o/1FNe1hiWmtboh83aI2YtStEw++tgFgGQ8cwSBCFKUG8FIx+7MD57PHfNW6FdpE1
9pnKw9vWunUPkdW3BSPbuF1Poqtk+uJGKLhjR3wTWv66rzr8Tdw9PUOM5YpNavytC8n7Q3TsP8pi
T/QsTYUGl4bKUMYPqEL9+VvKRZZiiYTBkjy9UVtXe9/IRBVUVJnPdMC2+65fiKAhz4GAuoy7r8bt
TJKkwni6+tBWfD+goD2xpm+a+YAywIj1tBwkREa9s2a4sfHFCshewkuDwCL/cnAIKXbx41C3/pOj
wRpWLX71luMQSoE0ISvJWYvMUd8SffVsjw+SZb8CfvC4Xpg5Tc4lbkm70H7qrLWfhcDfVwUN7H+Q
Ltp2CvzFYQe7j+2EAFP7uf0xcAd4FVcWZ1cX/ioA+0EUkQhBKnTSaS2VRjM3OzoJ33qutYuN86QX
zjvhZPQFTJsTOAbEweMc5oSf+BzlhJ0Pi9WiZqPez93gKPPfKYRHyfKFQB+M8ij4HQLv+E0C1/RK
oPlKRVFoiwEsQT2Q0VcgtN//7luYiYY0IIwj4AL1SLw50+G8UluLB1b/oMQA1zVAlPmA+VDR1L8a
TAo6zqRnRq9pVeigdHvJoC+cclM2RnLByiEkLelF/2Sr8fGKqzeEr/D1/yPqQl5g+YuEkx0X2ASr
wVZfI28RVm4HyyGdsPf86hwvlom1LXVuAHleUHdXlvEZgKQYATqSiCELJvmFrzAid4y9aRI7afeh
HpLuPJ+gwAissrm3HndtHPh6K+fafowANyzLyMGoiKj29h4sa8129lbjCDeyxfXCDfxuCjZzFQyu
hiw+rGsNWjkMPPo6O3KmA+dd3vi8W8kHz6LafWitik/4BcMVqEnuEi8T5WetuWKMqkP5HXTBtqo2
jsYjN8wAox0mZ9bV9EI/XWru4GZ1gk8Jk2ppLswTNENUQ4zESrSdxELgdGTS3r+2mpqwGLc/YWYi
teF+vuQan99WVSvEhpWLIujApdmh6PEtnRif02yYwsvqBMQPjPtaFN7scH+l/YvGhG4ZXXElWuC/
W6jk3zJb9mAKGMLB7OzMmuaxYSYSOfmulzaB45O1S6uqYQ0Fq3sC4e8VkYQY8cDSXW36BmaZoDif
dpwuScshtBoRnv0m7gd/gCa+juPWe4haecXx9ArL/G+rmXKpwcV7q/2JleYtBiUxEYsWYQoy05kg
lwCfSJcJ36qhvfq8kjF7crFLCcWolXQ+RRN3fyQhnx59MhLgiiXDC5KNpGqzSYZgoU7vdSULRj4W
L0b2rCmqFOj05mCOVhyHWHqIJO3G6AZdX1U3IGyPsG6H05OZkDOfSf1DXm5f+XcandebmREsWt0r
9HnOBG3LXqT7QZA3VE8LKBTzjrGO+p6zTYffKyiEUQ/ShFZ21JYMe0mJ3qLGguVDQn0W2iSdtBJB
8b9jOUnkkuFv5oyNNH/mAjONgePkeu1l5PVWTpnMJg0dj5L85OSFu5p7+DKm0BKYEq4XXpn2k8Ts
9wQ2lIhQ0OR67ShuiZBvRUTnvZ6uVFIueWrsllsYwGdgWNBywNUtYLFc/fRNsxhY02EYV6MrIode
4AyRBHGhIJEfCMQNU1I3056MlqT/bAzQlzbUI55Tm5M9UVnNR4meUwfgCOK4WmTVeY1N/cT9MkDs
B26RVy1cPkZHmx7E8c74bcHUD/bMUKZKRSJozACATs469hs5j4g0upUwlSgu+Br1f7s/As3Ap8ND
UH+nKi/DDDZjflrcJ6B8P4iSvguOn6TNSQ1Ck8ZBXLVsR2I4Mz0Agdkhsoo0JKMesHuSkgEEcg/o
4/S+VeAHN8TREO0RqyZ0QPjuF790YHGfMc+ynbDflYFUwsdEiuqcphHKlyk6G9uPxo/isaU8DHS6
ZEkP6alzSJIAuU5gDB4vRx3mdAdF2gS5B/lotVliaketvM1lRW9TViNLguRBeG3xc7pHf8w1OrPt
Tk9gebfCS1+BQrlOY9TWqW//tDT3zyhAdrKCRdvS9RGRj5h/mVfgV58fpUaBdiv74dSzrco59Atv
fXamFIcrjY6lebQN+HAXoJpA/Rtmc3+ei2KuyTvaxxoXDOcSHMYw7EsZ81vRD7O6XID1e/HjZleR
bsupyJAB5vQuHzX8yjw4Iqe/f6rgA5T3J3rKzRgBxRy8mE88DY3r5Bg/cbQDXRDXc9dFXWmHk/I+
GPOGOebGH7Ut8eTAjl/q5aWE/6IpQ64Y+/ZmRwe0h//M2W0C2IqaJBa98iSopuLHbecasV/mWWxJ
G+hSbZdArIu63V0202+TAGmYmZiCJDW7LjFl78y2/v1V9YTan2XGJjgd6QWBkST/tHUU1+GMP/jB
zoYmpZyT5vHk9J3zC/dRHI63y/VrMbvTFJhhB+6+ujRh48wof4pyxkiGq1TFV8mk96+8F5CFkmLJ
M8zt639/gV8jd2e3nJ3L0tuuJtwqPVYL6K1L2piNQVJ3tKXOPbPj81s0zg7INS4H/mylCi/Ojp3Y
YdsAPWBKsnvt9btOb8tvHrIYV3zumybGIXVCX+AhXJqjeW/UuAG3lbU+63/ILeU3cqthmQu4RMp3
un9+GFAT2fAM54eUzZquvInXTjJszP0UU0dxTFHZLnBDOOCuoaF40Z1XY5ZBHIwctlYfryi42f/i
Y58LQzHdUXqpfvAPQoLIBGk75011P00k3gpOPTEvNkCXA57LXYCa17RPilO2pp0jJ44/9EQBvCUG
qBF+PRlztsa0s1b0jY04EE0tHz04VeKFad6euKB/nQSTjrZTXERR+waYqjouxNOYIrS8/GtBmDBa
4d4dNIGQxrrTfO2a7ZjkL+EpvXJJ4JlwWnbLyU7e5Ae9JcHnTPg3Th1fKhgpSEySkcfYWlINs2ue
BY6VrkSwZ6uWVqk5xtmxFYX7cNtsOF11a6w3WQO/ozfTF1aprzVDxyFMa7e2C1QNT1TomKL++K6V
qkoTvkMfjpBARxjNK/CESOzImSh/tLoG034k8Rb6eaoKUvufExMJdyhNz/IjUlmWa6Q0THoCmy0O
1VeR9vc4fTBZLMi2TByie0ZXYe7h52iu0+uuUdko9KeS1xB23cJ843zw9K7S4G+9kGOjaHYp0cUu
4DC+nBQ7a0TlbPdDSjnNHp7syzqcl5yWWyvndjXqRTry1eXPY4KIy375fta+zLeQrr4BhA2kRqeQ
5LlYLHMWlvl31zwZ98jZnskkhmL9qwupxztFtGhcdAleEkCPrE6AKpIkBvTS9LwXgchTCsaJmHnF
LzeiuFW/YiZnyJqqK8HtphnnAmsm7z64z10WXifa/VkkG+SODHy7Zox4J2rb/S8nTzN1HmL+SJEw
40A2xaSlfeppROTmbviiX1i7iQoBQfK1WVvxxoj2BOZw3rwsKK8L+rdoDFYrC1Firzu3DyphU0sN
TbdFtTvz4o+Yr6pnfLOgzavpbc0PpeyCcjbESoaqla4evoPXeOxokJ5Sxcrwa0/Bg596xl+KuAqb
cSknzY2CbA1vuHpW0WollFDv/QZdNXODPxL9uxumNdu4tY0AXP7CeHeWi/IBXgZKe24BeW1SrYEB
cFfG2SraFjllUJOl+diHut6lbx4D8EtxNfYWksUrZlh2xXaqqebFWZ+pImpJ9RsnQAkoZkudBqLD
A7mwTWcc1TSh5dh3cLVEPg3V2CQPU8pNfAfCHTKOMMQtcOuibPAoSThn5oyJdtv4B8Xw0soXJslL
Fy1pqZGIVjaI7MKZRvJh3Rie04u8z7NDkH34dvqxDiQOq7xfB86VWwrkUrwwI5vfm+6teSrxfO5G
GrUj4cwwW0PqLJXIBa6eGB7DQzCb944mgH8E1TVSVnNGKpRXMfc6hcKuQibLppoGa+zTJZW6QHhk
4Z7xOP6pzs3x9AqUgNqovLgiV9/aAtPsjafbsaz+3MzjvPjdhAFqfsYr0lSC9G4X2udZkKECyGAK
MGc3nPviYHtgB6a9dv7UHuPwGaoBj86OuTrpT4QfMlzOnKo9/tZkwMBq9O7c3KKPWfgkZhMLlGDn
Mrlgs+AMU9TT9/gQo5wf8aEz3kqIXJXzf1MGu1dsn12IyY78mZJ8S8dcKzmBaAs1CcKbbuSVhEkw
aA4sygPILxkDWwrznbqG1J4G3XAET4dBrFLbZXYvI3ZNWpMW+CAbq8n1Q+0wtXwRqtg479dC/1dY
504OSgptmF/Zf+jJEcfO8T1t/F7BytEVyH3+OoDM1TbnJcjNwpkFq71HpF336VOoucEsDxV57a9M
w40Zrsn+DWSiOVv4a8G6rj624jmZzgYESnM+OTbePkpdg8kk3MVyq55/KX+OC2he4IElzHss1Q9F
0wdA3lNEIq4JhpY/GRYgcGGvLHasHC8RCmGNe724KvfY3mCjXhQE9Y06+KvWqBB6wLfpK6ui1i3K
LrbVS3u8RA/Ci9G+0gJmNaLacwfsROQmGrdj/26b5AFQcU6LxMR44Hb58Smzh1AjeI397tc5clEy
KXSZ1NKZIRh/++Jzra22x97s5VwS0VauOPGirWjowxoGrEw1aCm9F1npACM31bbvgxPZXix9qI9c
+grF9zmwmKjSHgCn9+rFMGAKAD3EQ0IReCVJcF/vlLQB9z8n9GzesmsKy6PLpTkv1a8F4Rf0t2lc
4jZxVqOxsGz5xDQwSSdJ/qEPhmPqPEsfiaDEFlE67/QIzVdLQTSAZBZKPNkrQ90kJQcUkb0jMQci
5xq37Nb90xh7wTE2QQA6thl1mXbnG1eYMYY3duKo0BLe4U64cDK3ZOB8zFQ4gxtYaCA72lER4aw1
bVEh8JGNzF1M29bYG536DvXkbRwJpEAk3pKpEaWVO2pfYJcffV7UTS6DqmkwD2uWfkMbnzFNFDs+
85wj08YrD2dHBZ4/34vMu5AnE96p6kB44ro47gnub/a+NYDcZC2yaUmFsxhDSR/PQrOQAwxuJNek
IGDpG1yFFBl8VhkrsGYhh4tgR0nPZiQf0z5zpVXu65IfFv97XIBe1jeOzBfXOToBu+vJ/G1axSQ0
mk6m3UYFG8dbwTT52L9dTredoujbOvrPXCXdS9VgatmZK3Xg/rlZ333RG8PkpzTvdkI/NoPq1no0
vSOyvO6dZrCUt3vMLMmYhUDEEkFAR71H4M4/iwWFqE5uBAFQGOt+123FbTSfpahjgZPO0rxw6XSM
Tel4ZjnGYRFHM53lidNb1fTRjEHhYceF1CLXaBJ3Z91u/XQtifLJMZyEWxg60ashzkcM8xZxvgLE
ZSmDfqX8YTFrXbKhqjX2E+SWU+DuikTVOVacQenS0TVQmvbBLX4Ib9poVsQ9rNkv0XMyC2nYs73x
7wyVhOFJLSeqAvxqfge/64oVp/C0HI1T4KFx0+nu9vDkIDuJmTqnF+bLXay22O40yM5XHJ8U5FT9
XReXjMH97uQHZ7D6elfSMImOpDGz4DCnsLCRlnSkmej6Ype9EIELda4AmaPJG2+H3g8a6IqiX2Kq
tL0gYIVg96Rkt0C50njsnWlM0Lar0qw5ogEUiSrAEXaXzUbY5s27u0+N1DuU7PDe9B96MdtgJIre
pGe24Sp9pirJQEpKadaIITE4KEJH8tcsNv50BtdbHL+1kfEHsMVjTq4Q+qUHB6S/bfLvcFrHNN4K
f5pJt9mQCGql5HDHoWAj6IVSA6YIU8U4DWNUsQLdXL2RVApsWQuy3jFH+IXyvn1gdL/Kjo7xCoo/
uczlRVU95QCbqUnq5jKO6YhPr6/2omti6SVDTb8ltniLM1vLOpiLd4FKpIdm1QzMf/LBPAorU44L
6VqWoLe2orso9SJwetErzORX+uKLkEl1xIv8nN+UzF/FjB5Ny2/PFur126hxvnGCe01duRv8s+r6
F7oJ1jxiGRpSCXM6nFxnlvdSZs3TGJM5k6JA92KdPSg5EYag6P2KqLWY5FqB2YYyaG0aAb3HZ2s8
+4ks/K0ZiAV6MwLlTwwc+3AKycQmbqQVPMKDuFkSv6MjcQ8Zh/FJa+QgBkeDsEJYapLkQz2pCWL7
rilrsCs9NYNR4TEDiN5jxvKrxdCQA54hfJcFpyEyyl5qtyDUAzHDxPohnEfETGU5AGuzBd45UEx+
yZqAkFtdsiVkiIuM72VZYgJIvKNPjYk81Nwt5kOCN+hGLvCjA75JnH3StiSaRlGlp5siJMoSKIZG
TebqCoP/y0Ti+60E8wmFW3pY68dawDVblNS1H8hNOh3nCo1V880eipkJ6oYv/FyrMJMO1LIgFTno
hbi1gzcKLOuSfwJ7sd76dCrd1jVRu3KageZtyjEAvrVilWam6nuhGSnnjC1mhJe43wDRt2M7hxpF
e1kACAktQyXtsWHBO4AWm9f3SHeAUEYIBH4korTnJZ21scCtWJCvnm/7S/fcG+SEaf8mkG1JYrpV
rJJuRsucW9AOugUjXnNTaFRdf3H9wJsRbjChoVuDZlnZ8O2Hsubq+L94+lwZaU+q0r15bL6lxpbH
hRvcc+MQxr2d0j+poFoFD/g9UvVGdrIFoAY83OmjY22EUCUe5wG1xUYDZP4Nd9FFAVTv78mHoF3x
/+nQ6uM0H8euHG2Dkmxv2/c1iWvejpSa1MfnYhu9v8k1R6hv+e5ShXOk3Z59/G1pl52OkO77PnSk
Wek7l0Y/qCfj6lub9tgGqExHjVNJB7tyIhOvEzENW9zrwiir1pH3i0CCLWrOzfKSYXF7m3s2rtRJ
qV9/bdniglU3zKvDE/F4qJyoyLsYfstOV1Vq8dnyBhhkTeK7WucwV5yZMj1UbLL6OQkFj4yhSz2q
eci8720B2LaSABcqiKzIZk6ITMWm+7AIRPt4hMm58T9iOrkNjnhnoV6pL+U2WnesOwpfrJxbW1u0
BZWnq5VxKm7zrHQh8e/Svm1X9rhyF221CpM0nwr3s1VGROPcha77FQdUZA50vLWt/cHkoQDGglkz
nw+IOBzey2iOIxCChsaWdU/u39XhhApCm1VVC1saicrmzKR6X1aNxf6Ch+6qfeCq52rIRqgF6PFO
tZOu3svABB4fNybRumQDLmq1I+ZjA/X1K9+3ubaoPllqFs65Y1YGhlkRvzeus8z3pUO7UwdAOq8x
9jihcUyjPesegPwcWUxlj9kfQ/AdFVc/Vp5am1EuZCTTPKjYKNObjXxxQKgw5MpP6kNIbZ1ux0c8
CEy34Z/DSYQ2/Yv2Y9CWupDA8KwPaJl718ovT3JjDFO3EimrY7FjrSqffnP6bwF/bfKFS1/MlVKx
yUJmy05B5nXdPy4yvRQgG/fWiEEGcyKr0GFk9LN/jxE+FybsJZ5mqnG1B9p+bec7NIP4bYEgc31q
tuvvfcvHXaL6NMHDLYfycQM25FMi1iq+RPSy7IPc6FD9BnhLhAkiFXwo4SPc5Uzh7zquE7N7HXYK
vhgQ3A2GCm3Rt2/+dZqJnnoMvfGNF3AWt7FTgV648rJcQEnkUJHhTkI4ZGXeoaAYytn4qEVxSoGj
/UdHP91Syi39ZTHoZmsnrv9mQBlOgCBtj3PiblHbHGR7SftfhDv4ocWJyHgmKB6iBp6rNiUe8CjD
n5PEWDCbYp2+ZDqd7jZOquwwQI32AwN7vA1Z5BWYVzwNx0dpxGSiKJy4vV80cqOa2ERlDfWf5vHn
U9OwabX9JEC1yDM7mtQHyodZIeISPUWhZGISrKF1nCs8um+ywWJl4W3NKGnSbVhoEMBY0rXZyRy2
r2+qcRqCweKQcnoK4DTrPTvhqJjKI8YscPY7gJpaQKYLHbP4csbnPgvKf7X256wfHbh5YYNQlj2B
V8R7SGxOsdySLZD71q2RH8e7U77EObpKJJomLM1T27SNX93LZtgdS4EO4FjH+1SCboCSAyrTVFlL
nf4jFjgaS2VyuSZfFbHXyReQzvxEmeDXnK+tvO822afAYqLv/DsVa3snBlIA7teRtx89si7lv2/2
4tZomqSiWnqq1+siQMOPbz2uGKPb42xgiHbXRts9S4hlzV3QMd6Enu1p8OMqqEN+hw+wccxoI1KJ
s4K6l52bt0aq2W1yFWzYP154tqbwMUTBnJ1Kh4qmaF2gu8iJXVVZwkP0G+RN2Dboi56QPFIxU6+N
yM24jL9FlBA00bQRFUtU2dyw6GA/tTR59x5OtJs3p9OmDwLS+6PWjYTuzjgxIZcRZs995kRQLJuy
kjqDeWXBZxX1xCRATMW4PpTDo7ib80Ojk8yEub7gSAhzJYlc05IIuuVeka4/9jy0qyfJW6l9Ex35
6gZXlYCqemhLkzBG8N2yXbApEq4AUDphanOVdwFA3EvnI9L8mBZnpPCgjhI1HnVxynl9URgSgb3e
ut8PJU/ab4VgS5A1OPdJw3iFUkqdgKQ2QHatIcC+yFDQyFFvcK+KL6kIrRJeua2tb9nj/glwsdbo
jhPwATJvVtDH0dw5Xb2qsJDPLFzMefpdvO123gCmtdxjCtWdCpDZaxjSNyC+XOZf8JoQpMDe+OCL
5lEBLhwomerw+JvXj06+nk3p8ga1uOMdoVbbcBgkCmr91SZ9zySq7SmzWaJsqIfqDCGLCDEK0KUZ
ZgKrzd3obFvBYg6H68ij1nD0+anxmYWQrqOvcySPy4NOZJa5sFuz5gNSLdVsBQQLz2O3ENKJB0N2
Sjcxr7D7X3EWOvN0FPSK/R7+IhdNZkcGmkuXzwGnQniFMmty1y7vfYanLxkWpAaJ8iG9Lyy5laMK
RAh8kyKZVmqFuWoULWXNSfzaX7sqe6d5S/FexK5Y3q5rlQHg3x4bIt+t4WtsTgpEx4fiwSyiYhOy
MFuA8Pc0ppoBqhzUXctLWdfK/YWeSVoWwEVH1X+XYuwjSUM7AA59VSr2jdecQ0kmXJVq+0HGdkUb
dXeZkB5kz9IvtbTdVni35wXaDR02v6kuiQDQQ8Bmrlqw5NTSMQ0Og3xGEgssVGdH1mTkkxP4LACi
PFKUGBrJhyYeI+l4Pg/F+qfhcxgR4D72g9hMwIXbWyfoNyEqk1HlqitWGAfxzabiHsMiSe/pLXA/
vU5O+W5/ygdCcFG18/1Gtl5URh6pJXNqv6K8Yt163nzC24d4u9C2nKHVgtvSWx+FWs2Ue/NBbODf
T0/A665cqquGGeueV4UpjI8bzABABtZXPG24ceFR4qW1MEcH55wHQoT1Quh1qkNXaqGHUMlD6pUv
vwZM+VvLE2oWSkP+RZGktRanJIEhHNwQWlElQiktWT+SKNTVWr+t7dfCWAMvsjdzUV1oQuoTC9FY
tarIh6K4swtMz/8MJCHBK2oQbIzwlSBsAo8LelQ9qi9bg0vkIndwJ2s/AnlQIEBgD2EBxkLmWlnc
3EW2IxrB/Ry08dqBSinB2he5jVVfEViBJzrvk0BLZl+X0Uj9d41Y0OxR0GhCn8lM6CEfAgTxHQSY
oyq67xXOGba4dlYbDl4SiOU9Jgt7ZmrXwQntRltM1AzOJezhkgh2mguH0nyVdtytg1YZWv0op8Mt
m/S4PDkEJ8mOYo51Wf+EhwsJ6RlQT0lMduUdaQtrf1/7vcgQGqvt4QnXSuUXd3vmu/ZD/XtNjzh/
4CvXnWjN+yolxqsQPPTpdobhtIKzDhytNCMAqVyy5phgHlEDD4vrzzqGBxOkNi3mHCSdkLh2v3Ed
1sBFjzxclL6tO2ZRI8mMrkV/rIaNRTcNRSuFf30E01DxrEvhQ9lu60ixTu5sR0cUJPBqvW4TP5Az
oDHfH/xtH0nP4PEZ5eqt2KKgr741c/+iB3a26zgYlChsZ83ocIGb1Yb2PHpbRLLaO5LOCG+wZEIF
yRWGYtVvkP82mzxfW1wNKCUPTPv/B5tbU6UZEjCCHA3E0AShIfLY8apr6rFrddy6szcM6EBf7FLu
lksFFs/p5+aOSobjzdsxrH6U6/ZNJDKRaHSUbHOizTkgSu90pvsEZpvF1rEm3scqjkBpIGXgn5vC
2FgVfGsEw6h123zSNxprzjbT0Bgw146BBcku3Qb63F3A+HgZpR9wY1zyVd+AoJQFbVN+KXwJfAc0
ZXW2kvAzsLGy+yN/zlqYbwoxyr9ft9PbcRjcm3xQxDl9+v59/Jb42VU0upcldBh0zQ1OZf16z8iP
t6LYhfQ6O0BpsRd3vxNtXy+EIsH/TdYpj5OVIwhYOrEK/NP8KHNddSbwGkT/+wIUnbUhv2Hd0Uqc
uoHbnD10t4ltl8rvLEgp13FYlc2lmJJMViU7GQiWkthffQfmicpnzwGCeeONviF1Giz7MQyDvnn6
DQNR7bneMhD/Fv4kWlfwar9KvSVdKdKGlNBLYIj9aR5Sil+AD9zNHLddg0JHrHshEh1KFyNiX20c
+94nmnWZ+eqrlfJUiqqewIdFXkyyOg4Gub3LAHTlvhJlUOSXsl4Hnxlltr0MeVWnAx5oKNdjoB+3
avr1iRInG9rI73uhBKPNGhSD87U0aEgWPwlqdfPJkwlDZJ5ZbzmYWp/PCtyaV3m6qjs0v0Z/bCdT
24AY0E+nKhe8lQOy7qf2GVII4PElrjMgTV+Fa8vWSy2FgtnY5ep2UJZ5pYR25EpS8PQuOovh9YVa
vMjcgE35tNsMaga+NOwz6IG8dICy5oV923tDI+r0KkQSb5koiMyMRc9vCteXBHcE21jCQNCUcMj5
9+dGBtcXMFHmaI8qIuqUalu0GGV8E82zI6PA1OCEn8r6Wniz+/wlFrlFOjevGa4FMYAPZDQWfCKF
SOTV5Wth5U+HW41iTwSf9v9N9KErRyQ57KWcvnv+lbASRjg4qQdgaoA4cx+ZN+1jlu7fRJq3dOGT
PFuEKGvuLuq8DXVS7R7MK775+chgOPj+K5gxPQCh+dTKrMjJcJLMKo7E9OJQeJR1+yLIcfwBfWwh
QEuDnD4L5oGnsZnqr4fBxyNhIsUn+Scl/xpy8jTe1KD38GAGWUSarJu4MXsY0JxtjtwNOzwEVLXz
LTHVrL7r48ZsNmJSxShnNoN6QcfXm9om57z4XX+hHG67j7kcJ1aFq0yb5xOtK5oL8gEwoGZ3YL+S
9bKAM8u1nA94Z2febMa4tzKY2HMVGdAijHsxd5V6KA9iuIxMsPUERPEvlFXLJj0Jv6sXY5ED9qQb
kV2wvBwKppbgoC0DXykh0dAkk2QYKBKP/F1lDWeVkTSf9jJx+YRDklkEwJuJ3uNbqxi6w5L1Bv/u
3pOdPPrTTRQX+7i5DQmEe1oOLPv0fv5dzlbLgNq21FqvUFPGepFjYW8e4EZ9tG2PuOZOKGVQJHy8
6DUdI6Q2shtn7dXyKl4wgDCz2RP6czFrm/4q0fnaxxUum6kleJIF8Uft/CcdZZ8QX/xpLhk130sC
gBXU5g7SKrLkMQl50tedB9L9MxkhAN+55IQ0ZkfihmcOxaQmjaipjbqrh5ImW6Tf8yivr6S/26rP
CoejBOiok6LZVCu4knr8hN1I9VliNI0IKoppm7cPTEwC8zLuVMz2o9OxtgTlufojY3Dg4GlFQ1pu
0HrTvwIw9ZqBpvu6GNneuxFoDnUgBJPtf/SQXF2qcJLEZcdMt6tsogzTzfTu3PpmDZ1Cu9Ow/Bh9
Ab3Zwels+zfmuidShvZXKs9Y+f1nF9NXwVRlpUN2XIY0OgPQtzl9gocUYmaFETrXRJ0lzy++kaZz
ITJNvuwM4/5CYf0EZOPcXajgzJ4OsChxsmYJkC2du8/71EdyNehvTtG1vbgxGao/Hd+xBR5RL8iW
KFOXALQeC/t5tJpm4R/WVeiC2b7ZfuQVyVlx1g7g047Y6xjgBq9NcmsimC3k1i5IG5X/oh66LiXX
sH/jdCuFkCg0mpHxo8E6E3lp+r1O2XHr+SDqTabefXar1efbYX1wnqckH+ZXtp48EPl5k+418QRy
vponm5U4sMrJz1d9RkY1u7xTZhuhxf00DOnAQrMmN9KCxBIiyFSLqBQEpy499tzLzKSinEXS4uG9
C/Aa38C8GowoCOFwqFf5zi5/KsGT3Q6b5KKaNlDFo7GSJNTt109TAKPuAb6hrikCGx8+5zE8lmiv
U1mw+3RL4n8nyXKeaU6NoXkSt6Pa5q2kRHhxyNKljwgqe0Ksp8vf3+/ewTgMXE1XZ5XsdoJA0BLS
4vt0VgUuN0bQKNJq87kOuJ9BbUBcSG85nfa7Fne1g64+n7+CuuSm/iyjuYIvOvXSAre9fhMsfdhg
oogEFi4iw/iYXICm0RAjSKU9ql+O4eC9n7bNlnxs99Vip9KE+PQG353ycCGWxSJF/vYtJbAn14L+
IX3h+vv0sy1MB6XU1yGt9EEsE4djiD9EDZUk2Oc4ei4hh2Q+vRwxIF18oyxhkdPpyxv7rmsDydVH
Cg9+tOCJeNtHaCu1Gs4gCn2fFkHR50O9BLN9A3HWY0+XrzwbXJUv34HgCBGkzHlLIsKs32DO9icP
1PclAvFWUa67Mr9FTihLwtg2ZnxFTU9fxAUBWXOnYeTxwDA9u1CvWTktlB0WdzSKrN3zGvIGtFwd
KqOOuHsdrwThlKj9WpnV3rrYnm2L7jFKMUBg6SUQyewJvOuwJVJdLEaI7sGstRR0wkV0x+iykQ0i
/8jkTMSBrTnQa0tWrlNzbvj6gWYw6vxLzYhdHdJ5cufASVYvxDCKUzJpmJ7z5qT5ug4Q3aUqLEzk
JvMGlDRmrd6gxcBqZ67bU/LRtZJNmBtIyeOIm87pQGfu6bI0D0nuFM9KS4/rNIdUxWKW/32Ee0OD
QxbFAN9obumtYxU03G5BMCnPKSlvObmNsnMpVc3BDw+/C9Xx/0NKqXozIkIUl6zfU3dbje1+MBLZ
W+ZpAqrMKbs7wIuHpCwJY/3E9ceR4KkpGt/oOsgHSKr6XCS1jzQvBWDyFolKdMnuAEC3sKKw5RNk
L6cfWXZtHnGgGFxN6+H4IAlOoDdl0xgqIxg8zEDGzKUmyUCNbDD8l7/yZQI7KzGY4ueM2h0aHkX5
zobq8DXoYwjjKKoT+FMWRdHivgA5P1wCPzm6L5JiKC2atzDQbFES+rUSqp7+/pPFrEaaeU8vB6OP
qifOXo7NB/xWUdJ7vm3VeSnVt8miZApyoFMNRKD3g09RjGxgec9cvhw/Z4gX0VH5svGdrTevzNrw
SIZYlMrwGuB0tCtGU6A9toFULGvd7wKE58aNyzt/kJTUMU6HgyolwdCGBo+p4XK8ZBqxNiikL8Xp
9e6LfIuOkpROxwPrB6G+oM/WwOWAaRrl/H3Z1g2mFD0g5Tb4eQDKJzbUBm90Vrv6FseWwj0jzw9g
R1wCyWQ3wKqE2nBiX4xjy6Ywj9o+rY607cOmeoDwiwJd2dSxO+LcAbKvs0v/6uA9v5nrMmzRGRPV
2I4WbmER60whHQ08PJ4LTlkYgT42J5qekSfn7Wq1xjG1ujJOjOa3oQipegkBJtkab9Z28ScD6DOy
IkUcShszLKg6Xjp+JeW+7jEMKij/qmu/TTeFJQz9Gs7QF0TKlqviy1DB7D2k8W2kGXfQVO4AuSok
/a0x4kkhg8NqUrc0aTgJRuD+E3/lEpBGD4A81pIj2dNHzzRec9WGMn5o8i1ne7/g6HsyLnUMlhfb
PJF0ciIqeTnWQi2IAXfAAyY/VtsJ4td/S0/3b0P9aVSPmJxsTOBzUUafeQiqml0hy5gRnBXjVJqL
NIkJDJD6ldQ8civ1Yt4PRMnNy5BCGcMt5jc58RTvaSjK7pEtUyDTEYshYCgLR3izPgDVb1d9RJt7
HR1mGWZxKaVEeVK1C9KNrm+CO4STrsq8Vb+KyYYuxLqqQn2DDBRIBEruOkEJoZg3qqpd0oDvrF0j
lRvKfjV/6o31mTwNAApgQrDn5hMhp7/WtAKJHZrNqhqdJycJxeJMZHxDMQbPXroySm5fXJBN4QpB
xFxU6vrrxArktB/vpCd0Ms/EavQfq7mo+8qYTJsX4ScnzJOmoqPVSzIuVrbembnyNffemync8C13
RIMkS4joG9toFU3TRAkRH5kLCFC3nRXsSuirtUerrCs3tthzLdgyBmc31UPC5srD6wc9rHySUzrM
ZE9SSCcjqR5RJPPAvUky1hq7WUbtqfE+vssOOUzDTPv5GTXBfsaLa9LPZ6xMNfCJSz1ojIsTfLpC
nJF31tf20puVaZzcorZoqbqKq6KJ8b1PmQDUDWvTXqi5y2JQl4DjEizQ8vUFU8+v9BZ90r43WsnJ
JKceE3L86ZGZg+AiP3lkljDOsQhrO2juNMhyHzTw1P+osdWa1zacCDVf2eDcrBryJiH4tZfe/roL
MVEh+JsL4iEyZDY7H0OHSiUwAnZPoNhhAL46zpPdt6izYuNKQjIzRo9rGRXuNJaHLLkphn9TXyMJ
T+l4MZTVwD60RZ9O1peH8Gaa+dtVNuGijLMKqkj877ikQJOQCMZooLIRfprdHaz3H6pzLWohN+jb
dCJdXXWDS3/Ea5fTMooZgYyngsE9XuoWls2U84J3VPSB0MBu5toC2kbFX7fI6qqYKuAXtOFEZ0w+
gv03r7SbMMSaA8CIyebqVvRX8ZqlQ5ALjWqaPi1AlkvIcA2t1IC1tohvCLJPJ55hyoT35mU7+MqM
iTjEOipkL33xayEefFSJv3Lo2K1HX5DTcewf3t+QDTTJFlHbN9HAFMiLeBlOQpYc1GYnRklLRalb
3lcMwdP7D2nZE57o76rrMVmzqTVThKnqv0S86GJ9u34JL4V/CdO9vwlRLLkUt1VE+A9XbmTn8ufR
5BS52C6kNcZuYIlFBMYhe0fnnDB4AbE9nZIIrYjbbb2wnrOgaKohMcoU0Vod8+gvYm1YaWZpJnwv
w/YyShvbQa9hSXBVsoVn3RkdwguidVGG0qh8ftTcIaeQTTxCQD9GLN2i+P47H9ZvVfcPVvVHpL1e
tskdfcZW44crflxG60hGjMmIOGEca06BImYY6aYxqGQUBNyL7Bk8w4UIXyVWrDa0M/gj1mzegdjw
yWoFlkmuxTx9T1A/N/Z+ePjUrMptH0tyyzCObh4DqA7CzWrPPAbAy6H3tQIvnfmIAdflZ/9Qw/4P
n1YmUzwCgYLntlP6mXxF3zqSYwzwZE+notwhuoL5/skgKRTWOjwzPdWqWDSY90R3sr+eX3yL1G7p
qPI9n7stEb3rnZUTZ4dni5w92hHWJJ9tVNZ5VXgmRNEyR/G3wOwxog+EtazdF9unsnkpGyA7WRP/
BolcmghO9y2HORz9BmaKQRR7wryBNwJMAceMz1Z5/Q2qlmRkjKPSvLQr5eCICT0qvIUc9/yblhPN
wPBJkhnUItD1Pa42z0TwotP+FkjOtimLJOpUrRUF6nCZCMrMxur+Asst+FSX8gGBHUQ/iqVjUgnh
YzuTtWtnWcpcRHwYjOzzCkjG39uBp1uM9f+SrADvpMuJmagoHUPBklBkGbWM4FpuX7MqFdtIZoW5
auj5c8F3bIKIUnmKnuu1WGJHn0JOclwa23JdAsnWwiCq2p7twc/SHgbNoTHiOz18D9lIsz6J16ex
BciQC4DNZawKUjRGoDgK44XfGoyI0xb+jEGVFL4IZlrKbbykLHHNyv/2YzB7aAK71QOa0dMwNCzQ
cwF8P6n2vzQ/17JBiGwXQ3G8A8fK0YP2Hc6Zr3UVPc+G3UMcV7xRqUOZAdM3yK7vne7gZ8uwUrAc
Jp3Tt34KpEoPvq4B5DXbKDH5SB7AIt9RaWOU1QGRFD1nwX3VdXm+N/9vBfYvv+ICv8RU4mkbpAh7
xDVaJ90MKySvJqYwIsInO7UspwbN3dO62MTuPeO9gda3I0ghTpcEsur1xhoym7bVUPtjl8hHreSR
wCMYFf8QTfIsZ32n8EgppzwiiCUG9EVNZhiTtQ91121pzsUU9B3N0SsxB+DMnDoxJbXpRiiTPXOY
o/Wm1XlYbM9RD5f6keWgAkbRhjiucwxeMyjIhp78MipSp0E9Fp0FP8Z30QdXy5C7wpfbEl4R2cec
Z+sk5LzrLO8aoI8qeNN7/XKXQ7MzxumJ7xbfbFUdYRhltEl8AJ+304SGORQKLL9J6BTfoIHVViam
oqtatiU4X22oKHn4UGSboNi/witwRW8dzd4XdjUnm49QZpPT1zYk4IOMCpdyy2BHKrWRiBP4qXMA
+oDPo3NlBdHkjJeJKvC13gHfW+/lvzwtS8zu0DwMSAAxzln8WK1daLLBAV9RADNJrmaupfXvOFDQ
jj6FK5J5y+bTsckZLILkx4oLdZVyX5+Jwo9chRPoC573qQAK7Da9LPdagJOjR4CbuJn3CfwYIykx
NCPtenKxehIiWfc4NNBD3qQ61j3Qln9ztDuBEcIIxOyXt8wcKAarkiWVxosbrOMHWCCdt6KI30TC
UvoEEQzQrEV3Rvi/C0NNcNelrIzAU7VFG/ECrD0Od3zL/KdYpiqIM0AbVcgodihRHwsUv+T3ciX3
kKzZm51rNuUM2uB1RsOFIpJUDhop0rISg412IsqwCQjWl42nfMhFv6vakC9RKKxr2vjXSn2GRxFS
VUJ6FRB8B5ENfzv5tdQM0l9oFi2BrXn444coEjC9hmPRMFnmXx8GI917FQDadDbGGjllNAKy00hM
IzXsWros7phhZi7qFslHhgQN30ahYgB+ljVsTt5a/cwP4qJ1PMD/Y+xKAuXWPio4PHbCABQx8clS
LfzzxgNWIPwMEWDM1klrwDEYg7XVk/nuMWXzQSu3/YTq1YmcIunW4n1hP+fv/JhiAQvkWutA17IG
weY/gj5Cp5cIY0TglPXnnotdtMjH/Ow2B+xS8kdyc2gjC8LMnywz2Dr6etr9lxKvVOZ/jFTdLdQ4
jcGdFzDpoBfcz3OSM9qKkd3i8EzMbQl5nlubTnLazBq5ByrgpvBS7vi7PuTyy8vIGjxns3K0VLZO
jhHiFIWFHGcO6h+yZklMVfJ8rUQSQc/S9ueqvm/efxrNt7UQYev7PsN38EzAjBClGZZEQ1/CSM1B
T2SRP9XLYYZBeHYz6WgVysGXB0RebLPxtb684QKVWwdi8ba1HXnFANJ4V/BA/Y1rFDxPioViYASZ
kehrwMi1OU3zkZOeBtmJe9CTE80Y1cx1jFrAhvsU+6I3V27F358702Tx7jJNTYtUgzcH/ke+yNt/
exX/973YxMbQiiJH1mYkE16sn1H4EEZrHr9MYSd/dWloPFuVkDY2iZYlePe/gk/OU6AIDc6BW24H
zPFuuZQ+D6vHGRRaHGZX+HHiluLgh9OfG2wGuScyPkum5r5WIPr2cFcV8szMCFgfDEOYTPWhNelo
pXwswNDvs4VmHCh3P1Y7mnD2/WeG2Lt2jxp1t41sRaikuxkCnZ+9shvomJSca2dYiWoq4C1sGkeV
tX0sTQKvbVgPkFZoAE2s4+HvSWEewk+xMb4JjBfyvxDN1CtOnLagUx6wB3ymRJNtzIWcrafIicCF
K5R9euw/FmXIV7K5hbI6Wj1K5YVr9Pf1sFgDEx8PSsZKQk+IjRkBxOBDYJ4E3R/QiquKEUrTvwjF
nFmKb1oBkhF6zyKNXOxhMyqQk8iVgzYO3/vgYYi0sLkozLCyzQrKSID+bDVXAtDQ9OLxGgRpO7Ki
ojkV8om0tsdSneNbh0Z1ZHume5VJNi9+fTRBhGIDeSOPMwT3mDwlVa9esDLptek6I3XMt5hgBgse
V5lMy+EJLoC99AypCLM2vMNCA3YmcXwXXzjhf7G5p2qnxJ7qD/LC2WrGFrBSxa2DcqOOL8Ga+tgW
PTH+BS+CHMDmfp8qNHNE3y0/fiI/yts4XIeWuWAiTrInXu1Y1hoA0GhmpauCFBpMDk+im27co8QJ
ss5VzI7rUxUe1SvYWzNZNF/+XA+m60gwB5beH9KoFNZvgyWrorywj3ylm0JTEmT4U7HKUbGwD/Iu
57Q/HH/5/CCgqzLEI3WhR5porZZDUV22vWoSGqm/YkkU8Jjo8GGcwvzMPbMV+oEYYZqJNTeiXXwJ
w1EOZxLh3KVq1TtGPjyJRsgBvGqAISbXmc61iYeaWJIbtOTtbkYXEB7K2iSUC5YmTqNjqDmvTjls
5F5kFr59p6KJIqRwZPZXZexXTaNWy8QG1FULgPlfd6FKWvPB1hzQ2a7k11p3lAg9nHlLiZAtsJ9R
XFgHua1FFQQIp/draCBCCNwyaH/seazvxzzDDtF4e8jVf8PK94y0AqhqpqU+x2PwOmYncaCvbzcF
HjKs3uqwsPmkyUNqju9mKQlJqSJnBT5x8Z9dEqXd4o6m2v1JPUmXcrGjk4I6+FRvr2Blp5EbxD0O
YS9jb45ybTmBAiqkIGdmK8EtIhqXYaWAhxa+gsya+NALut0HhhWQ1qoScaQQ48yearJxpimurcIX
TSa37oU3PQYuKQnTk+e69UAcHZ83piJ99aTT7RGZ0Xbkp5sSPuIVJf7n+EqR0hxTDbaOKBqvCC+x
RYkYs0Fl1BE2TndeNJxJLy5LPaokBYkRe3pY68SxMWyXsW6PEMmsFsVYb/F7mOQcO1dbxPi39Z9o
KBjdqeCqxhs+GvI1FjCchkyqHxRkkb4zpIthEXIGw0+kslRx+5kbyVqb2tWGzjiuVWK91a0f0JYo
VUdYG/VFEFSf2G81Tzeu5ZRbUT2w5VHDSyr8X0xdR9flXcdwL/LVJJPPgI60HyhWbMa/Ux0swpHo
dfRsjI2ZQbJ8e9BSSJSzqRFzAI9UhrZv/gMMQsi1/ReH198s/3/JfStNW30g9icknd2RUYTmz6N+
I7KiZe4vLZW/VwVX3kHyI0XZteoaHRDqbU6NvxAUcal9ZJbyR2IbGFtrk3mylrtKswm9udUcM+Gk
2KqCkGFog520e4Pru6a25Q9jchV/ZYq3B7sHiKLMq2QzXnMdj0e5QaZuALcvAt8l5qJfDdhfOgXk
6YVjHLwO2c4DzfUyQ8ikNmAC54JutkMp8LEGgudwvcGk4t+w4fQJxmdKZEM6SGfBTCM0NJabJyqF
5QyqRZwiSZFyFzXvMT0fJD8KbBn+MMniP5uuTx5DbQ9r/WuTGN+hW0Yk7jDwHGpTCdvKnj4tEdJ0
uq8et+qqmIfcsTDBj5ja0aSAunrqNzs6CziDETJIhg1m2U1hjrHVja9IGMQRnwTq2Bq1XsQC9gEL
MCG7kCIjhYnNXq7OlJqd8zjxmI6ROfA5FdJHFLYHMFrF2pV5JLoOxjyfIPmLJWWjiaK5rJj6ziRs
bBV6/HiTxBLsmeETJ33r/hapLmUIotQHNI0MiJ9rgBe967qOatTQ8+vLTLpkgMCzG8dxDNBL5643
EoGqg92mWXKfuhk49ZrJ8XfUqddzNIww9bOGkcsEWE8RIgi90B3v1r9Itd+QakXtFxqjYwkdW1s+
ZSEg5dX4X2JESKEBQRSwyF3dUW+6z56RQp0wMigzVu5ruPKZuOtX4DWxmc5NuWpiT/oSdg8jtJpY
7HquOhRXrR6xg6qOQWUvj4zsJypmO4h38CDokZPBUMFfTGcgc3frz7xv3LFB3Afj6chNiYJlPySD
65RbG1uoYbW2ZwVU3lo7Aq1arMRvPt5DIpC8I06nOySgj2m8t2NwfjAOLcnQ+kPuvtLqXabH53dN
Afr/KCr199OhOC/zcAqjRFALbIZ4MCyFcqQk/DhpIQRxqV1V4PsXNJ/+2bLleGzftfe2U1Dt6N3V
Espbs3hmKjG/AGCTU5uFuUlo0/BGqxk9WCpM+GZtXjQauKL6Y0t12YHH72FMB/naYqkRExdg5SVn
HSSUI2judQul0FKC45uZrPBhLPU2r/fShWWmo23NJQ2MFvSsnUfhFoB1++7X/iLFflBkXy5ZyI4D
eJYyVaJwUdaTFKuQUXpEIHbeh3zYeE1STweg4LU3OUW6KT3shuMCdf8jQRYsPXqfQXnJ5rwBZKay
zmuOSda1psCGkC1J4zBtl1zR1BLBJFUdk09+ZpeV8XwgPoz5NAqMDigEeGF/zDxIT6j47LRlUmX3
4yxAxUYyyQdAW4ZVfMz6G426rqcZDCM3yXevQ0eQGMRhz4T1NdG2PdKhB0+MK1qd+5+7y8NO8p0n
SWJ/kcU2q74KfqYev2iAsxh4KPpTHSmD5k65e6NBi8QSUy7K2d6sWizXvGVtYJBod7qjLmoXy9u1
eO/KEOmzhyAzPQcfTDeH79tslOG6eGC3cqL8AVyvkt1e/uoE7ezJOky3+LfOlge0Z2uxwH+4/N7q
ntqnvJmgfdux3bpCDfYG3BzHafOWznuVT5mtHk2kssQzzVgPJp26catGreY4GY+ztun3H3hLejtc
FZiX6BxHOgEKeSTe1j3H0qqgIQpqzvLVtBJRucnvnlHUuhtB+rQAjbsnrq6ONYaxV5X/WOAZM/hh
Lb42Nomb9eOpVLmqDmoCuFBZE4JHHaPdR8hbk/iuGGTv7wJr2EcXDHpxWt5THYiJUuXm7LToMTHN
nvupk0qUhXh4I/4UlX0Ghcvu8RzUpUu46vKa4D41dwbjb85JWT5FhV9iWBtb3Q7OgEPgKhtjucnq
QFnHwF18KR4JQ/5Kj8vQ6/3dYbLS9nWki48E+ButasSNNj+evrmniaFXSEeGYyor1FLKRgFmxyV3
zWQdJzd4+nlUYZ7+NfM/JSPru8U24PwpsFg2Ei3Yw1WwFUPmNHpjpX3N4LAQ0PHLIh++N+hij9g4
LZU7zEovnQFT8gduk+eMwfanbFEk2MdJVx6ABhRuPmpHhWHPiqBne98Na+616uXv2PargqvtTCqQ
Xq9sYBj+QFLY1sfVvL/ryCmgLahk3Mxh0XJ/Stj0Ib/45yNEOd3YNHNS8fRpEVv4Ovs+qNpkntRR
u+ghsTaffuIP4velj3Le9kYnez8YX1J/7ZyjZ6SvKMXb0dccrwO6OyoSMvUjyVr6D1l8TiFg05kB
+hBoqAnkk2jbHfcqwkTCZtbqDslCocCneEeT9ECtv/aIa+yEwnfyB/ifEtE1/UsE0Soy2KhtD+hl
9bqPQdoAsBMh+2lZaoF1wxFI97xebT5ykbZd9PZ7lPljP6JSC4AtYvU3GhbrM25bAuAg5CCxv+rj
v2+Rgif5/+n+j1jcj/IcUxa0KtEVBtnDAqyi2wqqGWji8tExE059yfWYzPRbLwXaOU4YeikGrYqz
UKbcL/njYguWDH7oZCnwSer+zLezEaGSAZ363HZ5We8BitVF3YkcRImEubFnRRoQnmutI1vPP9pn
7xw81Lnvy7ZWDkEgq7GbWdNZ4GBS6O+Oj4QYs/BO6SQgyCRC5VXgVRuMKIT8XSMxMKlsYw3j5Gk0
gp6ImbQhRnDOkLsbEBY3cYwTCv/jdTVqBJ8GD716t9q7fapeX0VfGWAqu64bMBeXkn3NSdcceS9x
NsLkUDOTE2RyP9avwKyUAO4yyRvuhUlWLRYcsNeRp4stx/NAz1n9Ve3qQP9Kbctr/0TF3WygESvT
Uz2L2nKrMGHTZOCO/SKekXZKNBF8dTSiNOZVrC2IkTUUGTZsEdAu3zzkCIYrn2xbd4mcy81EMVJ7
lAtzbSUOPdXil1aUYIQYE6jOSFn+WLK2d4UVIgi7UX6qLSNdo/b0xeTt5KwSfW9IBKxgDWtWUA60
73ocO3bFLKEylydhv5tv1VcjaPV53UlF3zEEKFB9RUm8a+Ld7YxWeLJVgNhVjTghkuqIxU9bP9BM
TbneR8ZgL1ARLckQmS6as+Zw3u7EwR6eAT51iFVJEkmehhtHa4MlUrk834KiRI58Yv0dEg7ajPZl
8V5O5eN7Do7vRfykCr7S8wHVnEoxqhsOuW8fvO5T0cHM9I/mM3V2QZTCY763dliv7MEvtl9dwEIk
HeH6OSO9/Q4BX49Cuh3M4b3TzZzvuVKJ0032IlRQqBErWmqQPk3kgnTqGJkvxRe6E12k45sUTNPb
GQpdmWRU09UnOBPUNHtlIFhJhiwFIA1/HYX6lxDNi1uin6a14j3vGMC5qoRg5n0b0OEGneyfZWRI
HFo7cgAX/+3X+pP1l3ENn/uBQ4GRkp0042i4KQ7BzfqcPz+lNE3iwslZxVVbRPQxUFqLPE+Z2P3R
cHBIaffPPXE7v05xDYtiY0q7xhNYGHB+kKzZKGZSAJetqnpsVTyfP1qaIjMahosHoV31EJ39VPlx
caqKiOu5u85zaEefb7Bjpp18zjiCblat2D/OsUwsLJh1DqQqpAXWNAzNbWwzxWxB1c6iRhgQVfSf
7CCYwMtajz0bX4eTFv37FmGNH/m1D3XjXOveALk2uVErrUZXaESiGLSc0o0IDBxrlEnsUMIGVOed
DscYnEx5VgxP+cs9cGG1mOHSLZcO0iQjwkrsvS3AwTJaTPIvyEPl1rwqUH0nWJJ2h41IubXzH5y4
UkfmNoBiKhcycAHjZg0VjaFpVDyQIjDDLKK0i68FS6AXEAX+5UqfgBzvY/R8bVKWNJ8puSM0x84E
auDLwb3PjG3hAcVnCRhz52yvwYHVSeMJrFQ7jc5XNWxiMq9djLkVA/h8G8CYAFAQivELUhPEPood
IoAusPsvm8F2G2pAvItAdlMJK0rmRC/VZ8QYyF36Dthh3Pj5ol1dUC7LdJZwElVL4JP7WaykX6Jb
XA7xpuhrBkD/h9O+xtPSPwz5Aa4PGZYMOvWtv5h1qne1LNkR25f4tT0UgctOjIxz+DisKxZqMD7f
aEUvkBTRO4tN8C4LJYva5ickLH5kUBdeaw58MxZfXtzzhqmJMemGnJl2VRhR7ToScUge6SWSLM+E
zYN4wfl4oQ/v+KkNmrGKbvK6Jdsz8hZusPn6Npfb1zfrDd2QsPqxnY6o0ENplAWT3TKlxVJcaxyQ
0kKrJ5FbGoD3Io+4xEmRym7hMbs0m20OQBIq0rTYoUvrxswyo4doF6LRHqlNP4nkVqlT9aSNv3js
nZBMgE1U1VTnjPhRPcS13T8aQYrb6c7e0Hx0QNe18dx7dmZsnpfEI3xiFtOUK54xs22FgJ4ESi7p
TG1mofTEk4uOQS+Xy6oz2HI08bfVHWReualHiLzk5oLD0+wV5rUqkiq9qgoU0gWw92q6f5RVi9Mj
XFfFwaZtdet7Y/S1XH4YEP5AHQFZeCzGirluUab6vVHLQbzVafcpieFmzBgCNpVX0qjPDp9vZdS+
YNYTFyoijSqdCoYpoKfN01gt1FtlAH7f5LNp925AAQ6hfstSyrPEIBCqa3eGsYU6IzvdhUXH77ja
WneIsFa/8ffdSwrXo5FMCJX/84dy92hgJtLSbg0ZWX09cPeoaAzWLVObwllYeW1VIB3puuKbT4+l
ZsGF26CQnCqeDb56hcwpCdQdsbquX5o+mUlZM9uRf3WEI5SoEj71wPYsaRuFM50e7XKnkt9Mevvu
vHAtYDswofL1HAEK3NAkBIusvlg7ldN+Atrlhk3ttF18/Awi797drukbrPgX+v3kLPdvO6K0WznO
Qefz+Ku2WM0tevFASLUmyeuWIaLdEYPJlyx5yH5gfNuX3yVWOa9azlU5YZFO33Yb7rX4Itv3kSKz
giyhHU0I4HloFJBda8eb+csDhcdO0dJgE843iYuLBWDM9RfS19jI9rZp28+rcSdXYB7z+2TwP/ir
UkD1n6yoOcEtTvkVTUCAZcGJLIi1tP3cRH9gGJih+bcFuVMB+RHMTyLO4lRaYjzN6qLozOI6dxgS
YXR2QF6s7RWsyfJAUgEp95gIaiLhstYZnkpcWxY5tsd6pxT1CgAcXzAaP40TiugNXlYE1VDZNJFo
BbZRuuoqSIircYdsI2TWjnUYM3OA49R4V0vdB7NasnOps60+zBfgCq24MaEdxi0tAMFsNzOdz/Og
BkQ2Y6fjC0ljVJ6vaGFFjDPsrmJDdfxeI1hpCJNBa85kbf1gyoXRBn6fg76Sp5krej4dmfP7yZul
Xr/4DtiMxUpQQ5101nC24XUUV/A4cZJdS5HWzTD/lKrgwaV67i7SZEaVIq8EtiAvVll6QYVsF2TR
pRchSmWmD3jWosciFL1QXJGd7FQ8JEtmGSpqkHItEJdnjqmdfTQQrNUEdaHYgB2K1Iefdzl2vTjk
jzH+lGr5YztpqhALe58+U5+sBko66fzakV8d6DuTB5NgWOWvJX70VilpBiYCTSDHjKMU8MHc3l9b
qVD4rLk2CdkiwvaA9MQN20tpVJRT9mEmcfPYKph0SWfuyWhCkIgnkV8K8LcThzlq6USuO538UpYH
avyFuxbnpNPhGZFdMzUqwHL7r7s/J2cSTtwX2Iallx4fTYsfyEe9Ee5WgJVlHCokpAm2pMrffrnM
ETjbDhc3SNzNowpUX1XKO6cYrLve581ELOYbSS2o8Skp5n0HwfYfUPRVa0XbY1W4xRlmAaeTA3Ql
fhvXknUXDgh4sHKp7buw9UY9v65OIOUYITv2r4UCFeH5U00F9qWpGDkPCCSFUz9UU2XC2nALH28g
NcD5VxFulOOparPvAO0pvLuDtKm9snOsB4wXckRv/cRv23fXpWIN5CW0Ed5D/88zHKbE3+m9tiK4
47EWXh7PxTOmhnL320FMu5ybgKlQ7AfNNDPDJzSL0XuUYeOn61HyiUPCuJFKYh7VqpEejPZ3FEpV
JoWT+XD9KvWmRcks5C7Fz3Zx6/VQVrxC3Zp4s3E7LTy61JXnNIDyu5zKE5fbLQ1uqKQGuE1ioB5W
we72a2DOo+JB2WQPXWzU0nnCeLSt4oTBtdGSw50SiNJwyhV7Vqn1EV2pmcNmH2/u5nAmBYAbysI6
lhf18LBf5NveZ9qYRel7N1l60beQR42/rPjZznw+MNKjObYqc+z/QnVTGQaCMtDpdjB2vBI95XJL
Jxodid7wq4fIZsuPzDa3j9p7olOiM8JEYLVWqn9fnBekFZjc3HG0PTJ814AugC9mTy53DgbcJnYR
2E36imkdH4q3qQ6HrBdd1mNh+WvibNG6xoWRnBPQiAFMa5Pap0ULdt+8Jj1wY/eL3mYnK3krqo3a
jbDAE3RgHecLAwTlSqXbAIurGkfuQJ0fQNQsH0HHNapobtI2Pxks1em/qa09U8oNAhw2gXVM5omJ
vIwMID9mAvlvWbmEUye5K5eNHXLU4zQGu2ntIjZ0oCaE3yvHoO6bQeumotpcIrRnMZgwv7TEGipN
QgaZCWPYJBL5bLKRMFy1ka9MO4D/cGWpYguSXrRTTFN879pZkzyWa4VFa9bnThF7kpMQTymR3B6S
K45o0+zVw0H89z4sgdfbyXZj/0VVOKN0a9SGKT0AyaQUjERgtwZ67Ns92oTNLhGXjrtCYO0N76Dg
C4SpMpXfbuFK24gFWWgnuSREiI4tz+uMaR1LsHq8Wmus17djADnRRAcAMbZd0ryfYKDml7gRhGco
HgBdAJg7qoxVhtR6J+GB+WIF1zDFWLlXFXHmGm30lANE3yt5w+ehZuz2cv3XAn/QhMWPTXrBqxOO
wbqo6ho43qX/6yfMnM0De0SXFJKfZB+y/mqDXojhleZL8fwUIN+U8nzE4iK+9HiKU1pSkW3WsWIF
10z4Gu2K9D0J4bzmxk89V/QSa2yjTzNpAY4IiAWeeywYCvM4qfZBV6iqPDoS7AIZRgZRBhthGbQZ
stNa3EUVltCH9xObYqRG/PyF4gHiYubXgU+2XT4TgZuu68rdTY0CP/kg7JYE7Wrh6jLuPQEzNLwj
dN9UUQpT4qigcgCIPBMf4WqqwHNwjza5hIVlIGW+F/ldkxCibMicuPY2jtyn+1DZBgBmxiPM11rn
Gu/wwndWY4QmA7gqfGPy+kQe+o7MC5trnW36Wd/n01/2cWNLXPaE6m6QrJ13lXxfJHk+P/B8tRCA
cVoJGtrRGWh+gdjkGYjSaB+o0sazJOnT1QiKMZnQL05rnfJL0rlv5D6ijgK8zB3Vw7cGVyMy3ekz
7MflrGudqkpMsyxABeveh8+GZQa/H3wM5luMyJE1xONR1xfNZjsKuot2HonO0jRXB/73pFE55sQr
f2Gn+S8oZ/mD1dK6HmPNp4mSvaba7FdIWJqctJB7Vx6HO5kFxSZfwj18bxkAy+UgX0mqYcnrV+5w
/msf7S6jVy2yiGg6yAmAh6f5XE12gjzaXjvLqujVSYf8BREWYHKGIhI/fFViX/NLbz21Sue3DRxB
RdNjFmLSx7QRGc1Cfral7OYayUd8U1/B6DyL9sGrWYP3WGmbKnaGzJ7jtvDhX7fIJCg5sCUo9y8D
oTgrIncFEbKz35npKKPeAIyBKhLlbW/1FpcAx5gl26epLCsdYUVS3OnRDVG0iDGWGch6q6FFThzq
3PjN51RB20Js7NQ1y1IFdz+q/vsMD6cIfpGAFjljDxwnbJU32riWgFp72p7zLVr9v/vd5fC0BpkX
3vAp2tnsfey516xAZQLT/1rNnFvNYmUfUPXTqhBQzELEJpq2UNxwjcCc6nGYdwnQP6bhBjTuWb2o
76rlVJ3jGIBcTqZxXNvSmRVWFRzeebkuQ8Phlb+Z+Lf4D4WuVTMirpTVu0UNjRKoG/92QZcRwwr+
4i2NwHRPqlJ6983wAsIXkWCo6xkyaDswSANvlXpm7OQsq/HGayHXDHG4mRCQAo3rpKLRoa/AD2Q6
0w0eC9IHmGVMgGLnzB4CLzDxGTo0p1WY2IU1/2pij+0HvNVUbT2Mvhv19D04vhoXx8/CZnj8lcOt
quXhpA35jKDaLXS7EFbVWMDiqfvVC2snKZUiODKGy4/KGxiXGxha+35/2PPAy5LKG7tBq0+IJyYX
LUoF4ah58BznLfILt4doq1GGxbH4D4nB9LDxC4E71+K4w+m/MU7X6lat2Q3S7Op1IIttTVambRyh
IEAHHumjk/n0eZ0GuMNAoiNG2QJPG7bX27ThsfiKehXk1FitFNsPQxDKTsNVpylrq25nM3TanQcC
PlU6edRLDh/rphWoHmr0m1aGQqVj1qDKu+j2E70yyZbnBN47/I+YPFwERLsbpY5O66odUyPhaxJ9
FeZX69ieEeiHht5KHe6nmQOcKYC/U49lMRcmef7oo7YdEKQfW/fycu0zkDVlXTAzRkY3X/ocVFue
H+4QtXt1eDUn8Z/Tnt1PMSh+v9g7STt1TuWInLnLhoBDgvmD/qx0IoLeG/QLeB4G7hg6xK8+YAdh
P2SEW3qHclPvHmMDKzJSIYi0t5GFOrChtZyEWizx6SYVzd1IfSYHjMUVUzRqCoVtE6M9rzLlY9RE
2m+2D/ocaTFo2/54JwrP0vE1cnexqIJ7cl9cTcXgXmbSPCz0NYhpOZNSaXqYUo9+StzljLvLQykk
OGuewwedVwZwV4cZmc/ux86POcc6nx8i+mR73T/3Xfw40q+6VIhXhMVpZh/YwIijs8ZLDBqsPPjc
p7TeJdUNfLglgEai/fu5t3/7IORdbg/7aTohXcSr0+wmoGUomawFatAgHrm3a+k4IDUy280mPXlI
ZmaZeGOPdkKtDXto8JbD9bPdjF/1qmc8Vd1Oj3zvoOpT/zJpC3NZlgLtn4NzUrrtCyJPNujnQfgf
9UkO+NapcIfSu/x62RlKPKXnkYBG+pKdKdnij837GgAjI6ft3tiZWv8QDEF8d6403AryhRSv6LNP
trCH1VN9CoKWvxr9T2WSt8YAQt+xi8OePKw2qd63GhrVTqa8J9H1F9Hqwf47yqjdiFD9E78Xh77u
Qj7BtxnnYrMZ8tW97LCO3op9ESYL5az+TSExd55bnWLWbZvmaG8q3i7gkQsB1dq+AvU7zvV21Sae
Fb7fKwWPobTb0EhrcYWGXGBwq/q+hMOdfpkV8mQ6eFsGkEzBHAvsIXQGuXMyOwDuMGsyuhj3/C4o
5K7wqnRJvv1LTlX7xr5ufSIbQecPw9EOl2NrZ1foijJFLJFO1V6l8PSSFQlC06KOIwnFby0xDiPd
+hwuArzfeGLitAdMqfGH/gzhTnKnygpP+Qdn2YjSO/TukW4+cEQoU4fb8fY7LT5WT8/P6mt4XaaL
7ej7frHkNdmNEOQQTgKZhIww7q+Vsvx3thT8byyWyzh2Pc/OGCd1W9pRZkgZJA70qF0pAsMhSvD3
08zjZCp3L9nB3k9kcCu7pFP2Vzi24cJ2ZZINJjfvQj7SOqTyqwS7cDmUsxf1sXsYBsjIzgCjhBl2
g/eNycyYBnYyulUvIpQh+QU1vGB2mOWIGSmILx3zDcDiUSAnHSJxvRCGVR5pZpo9gCJtrfKKdyLN
n9EuUS1bEZ+KYKHM8Fov24BjNi2PHd/syqQo6g3pJl1TxUPAwk+T+cgkkPc8vnorzdy/m22ShRrK
MznBtMv20gCZZpSO6WyQxike06yH1sFFUN8/FoJoM7RZ5cWYAB8M7kKG1VtpBHkZstpn+aoLSJ3d
UIE4RamVXXdsDGGswM0B7IuqTQIx0ADUB+pcq00yFi321UlV7kTw8xI6ecjAHtRoXSJQyVNlnDIb
96wMX/+ma9jiBr9OxFNo6bwbsLhfmU7OtmuMptlfSHKLWYsAd0PUeTaDGbZNXfyvvTHMnow55Q7U
oJRODN7tBtA8yBDC6cFUWORqVMD61wNO2SyP6vSaDrFPL+l8M+42MO6qtcn+5GUH37qzLCqZTzpu
4M7AAgnJNWAVGvRCnWfNUse8np1S9aAdPuhqhfEw0SXw+MIJNjRv6kEXXqoYWv6A4WfeaiEgpt0D
I2wYWFVZ6Tgnh0cFx3WqGIPMftA00e0dRUokrcZr/8gKFJbo247TiTlts8zyLRWangJfXXOcpRbe
VoJ9iHLhdjESN38CIW/67L42nNj+kCNj610GMy56K3TxovJIss5Q8wdo6dk6tw8JCxlrd1yyrtJk
SyL7E9DRV/enf0OTP+AZjG21nB0esHgbXkSQVjCGWrrgVkV4PxDPx7hNN5ntFH4bT5O2WlZIc5zh
ZqigLJpErus9rgbRRAJx2I/lX4E5i4H9KmN213PWbOYIOJJJqNu9w3OSnzVQz9ig/BE0ymUgZUzv
r5xNwFSbbo46F7LTeP+oDdg4GKwFjpBU2I92BTSCAQEZrVeTFexc4Dly4gQFWYzW1plUJZFs1m38
FQQ2bEgtTpc5UceBSi6Rtn1RQZybepnJXFq6GPw4syu9Xs7MCcJuyXBaB1OHseLyIm5WubgdA8Pu
Tz1sVyT30UkFPOobrblfw0GDmBYQaVGJ6XTob3HdVgCbQVHMYnUEpV8Tat9lSKmZ+v+53rNL4JW0
VTssodA3N/iIoAsef5HkvUPJWl9c2PXIi2mzi5rxQIabTgOtlvW5OFCW7aEDNKAgGkeYIW/bhW8P
Px4m7hHaxNdV0FBYWExk9KSGFVEUcyrJzqvVNC8t9HTcewzbWpObsnrYrWPEa/0xElkFoE+xChoO
GbYpEpu3NnVmb56PNA8OV/nO6ajURhkh4h30UaakU+c+KUx6lawPlhuuRvOfahBkzu29J9TuuKmW
OVzlEzFDa9yBLB+xgpj/p8Ck5+CKbcVHDYToAoiQQ1IfjfGU0Nxj4Fdp/g1INB6MMQ4lwSJ6SssZ
D7Jg/EulDBM1fYqhvQF6+vCjdDQeNl6ZgcLu19aSdpK6ZHdCZrY6vDWyHhxEZpyYTdMFPvRgMGRn
L8dOGhfwj/N5o5O8E8mr3UbOnsHOSgF9aGtCX3/0urg+sy9MUBTuwZ2soKXz08ZeRqaFGE04Hurj
Cgao28cHeS+lXFN6vGucOCiH4XjyWDbqSvcq/LyiPvedOz6U1wbXWoUTONWol0Rrp7GkqUtMXiwT
YIdAVuaM0Nv48Vs1JIpOL3xg7/E7jX6I/DckqPgMxbe/Lx3dxb7V6oVJOEL4fSpQ4yS5Bgs7ehrf
tABlZByHailuGvnqf2uRlE2Toe/PzxwWHj2Qvjnkzp2E849kSyVB3gfo3JydcQYDmRJRzV7bchGd
OZbtlgaGp3O2VqIzvaA2DdtksDgA52hlghITY5/N/FtbiVHA692dPNKQihbVmmk0X0TyPVor61wX
8Eq0RiQhlCteEjlK/uU2Pm1HkSnq6z9PKXcb+JP0b5J3/sHz9yKt8gEkvqf66I5NK21bfuYIHPkj
UwagxlIPGXpFf7Gu3H0fdX/RVCNaM606p2PBHu4XlPqYij0k+n3aSW8U9UWVsy3X/QL8ljGfA/3+
dBNnz6rCQwY0/5hMDoGgxLuYSrlhNsgQuh0mpnQJP+c7iFrq5Dj5Zi0JsqwXx1kFVdbZ19seoW7c
rYPoj1out+QJZ9ASl3xMS0Twxw9YWc6NhMyCpJ6dpEDzMwy7LHWG9VR3fBvSqRtgK0php/VHhBF6
RdOwJuEzjcaIHPZ89fccy1Gw7LLxvucpKVl6JVO8737ACKC4okyoAnADSqayE8XI63FwwTdvZDU/
a5b6gvv/YhwXKVFuwjXcjQNQTcfHuiF7PYQz0oz48UjFcOCsmIAc9SjF8/w0fLlZYT0rjlHh//pc
ZEmcPZW1bv7m43NwE+yETHfLwRQ+yh4FbeA6ebE0Vh8MdMH4qFLFYbeBmTSd90yvOI3FQlsma8yN
NaF6BYsaXHDwCgUEo3pk7OKmm0VQNm/c/6RgnRIS5L98aXF+U3Xx+QhiUgVtMdDZYS6tgHN8kCKl
+ciCDweLMXcfQ9nXGF4FiSAqZNp6mrbp5pBRZXpMLVRQ/rx+SW1smFnCAG8kgK9BtrNziKWy2lE4
BEboTFVwx0nxs8KFiz3QJQmT2yS2b+V9yxdwCsWGsY+ZrMNLE1qCBTD2xdSTGE7punSBZgiyn+yp
CZKke3B1AC188bzUAx4qRMYpupOlhUPMG9tnhbAjHwYSpD4ftK2mYCRZHXS5UI+mhiTo3Z+EMnl7
ZhSxnpXt4Vsw78hEh2UxisjHDeg78NxpnTTfUFHptUZnZZ+NA2EXKD0/Ay+oQ6P4q6e9mI/jCP4n
x72iHtOvElCFgeV1dEtxy+s/rEBgWUHBp5r5+yr4rtBYg4vOlJ+2ICag9nFF1sTJfKzHHQQ1WyEX
qvnKeGYgP74Kdd6zKKjZcUgZ5kPCFmHZ0dfTilQDk9kIYQ7VEVY1b3vrvJtJ1UjX0pmcIkA9FpfO
U/CCtIDTFwPlY6uoI5yrkFR9pb3fy3+5TfwFJI/WbZ7j3TbovpGJwqJb1mAXhBAAYlfljeHhefy8
lT5UdFPOv0EDj3KfroKESf61v2CEc2SeGLYpITnGPy+Q61e0FKbAS7rb0z3eV/oeCZVkho6c+TWU
vmUlHymn6oNgUPOOWX27C+dmlwsOfcwwO2wNJN39vBHzJ42S9Tkb4PpW/hMPzcVd/qQ1ywSfY8fD
eUdgw7i7uihwJAcmkKM9bfOcRy99L6KDt88xShpft5RquThKvT0Jlp/sqdl+xuU8ji6YhHGBjaOt
NDxYTY3F0UvfTTkVUYQvZTQD9V7T1FkEGZQo1HmD8eh1nNZ7G7lxqK17XztjUDAhqgeR3AXcmGc+
OUP+WsAJyu5ninM7YTYHKo3jT/PIjHGNzcy4jiFveJIzd5be85bSFhcE13eAve7eaq8zNI4myDfb
vIKbQ9096ZCbGgD3yXDPt7KieON1Ik+VgJ4krPE+2I0UAV0eTTFGh6Xt1z5nvbQcqioxrIj18nOF
xSuR4OIWr8i2iOADklymHlFkBCcG5paFpNlgyrHCcHQddW07OKjVl/hCQc3Z7D6U8J/uulChFP2g
IVZ2h78/SONHoDJuUj8qUAN87g6Od+GLaNnHipSKJolFF94UboFD0Kdn0fWJpKhYyyk6bPNIxH5N
NLFmIEa6ZREbbVXctA2+03sN6tIyUZnSuT76uEI7HTK/mH/9YipLUoTW674FAS7ii6+P8eDo8qq1
XNBQG8CxyLsViSpIaiVJx5kcaMFSRj9c/kT+PJ6SMbbGsZMFbjXxesEIP6IGKG+r0AgO0DcoTBhO
y0TZl5O7mcpfJ3Q+CpiV1jmGTHlhSmWW9ObF4T+yVew74rfDQwjZB6DeopThHuO4zUk3bgvPFg+E
yD53YCL4jPWlcr9QwCRtD16+kA8n02v5el3xoVgqdP/Drgev96Q+WB8MPXL0kJNHBfulUSqxsRnA
SdXHPNsuEKficKx5LilbR6v9+ua+B7ryIBcZ6mQHaI72chtTe9Z3TKDV6mLrckQTZhrRWDa5lWQ9
dat8s5ZXrrb7IxAnrkDyWwzkYU5GzTzUeFUgi9MMteSWdLQ6gaS24F8aIMJO0aYpMta/THRU4bq8
Z/qJ8xJxcJmYrxtHPSNfqUF/9ZTH2OryG007fxYbA3jp4PEdkQHv5oM2n0xftJk/ntB0C9yq9pyH
zqlTJxx8dUpqp8g8iw8Gr/WccqtqOCctfZ0Mem82NDJsG35etxmXxeysdKUIyVzkomk7x0De5hf4
3rFJS0axBx9WHLsVwnQ51GEdWCWwnHUQrLoLDJ8dGJS2OepWwRPvoSc4R2uhG95wS8mCtlMNFdDH
K2zynB8FBqdVi7DVEYcsviDVo6pULJOYg2zDZxc5gB7wOvmHkdA8Nz/iafzO3v+jjVvIFcw0jxPv
40ZNkAU8Cz+J2NLf6o+aWjf1E5Siw+j2PWThynEEfONucAgur2F5zFpDsagbfjVvEnQJHuYk0az7
T4sdzMRrOtJKEPRkBaKqKxZUv30Z+L0f83QlUoNO9GaWR9r+EPiE8yDNIYa1Bj+GWbfouesYbwFN
tjhntYB+RXgpOUWw9FUQF1H7gQIOWcRs/w1Z67q1F1jOW1ud9Ow9andChuAtzt614YTTdg/FTLMs
SGlV2KeS8tEuTvHA6vrt2pC+kfeUNtbeE1sFG50bYvSA83u+50RslpTFr9qOleiitio2TD0YbMug
RMT0T3/VsK5EFuThdoLjUQBxXOEXRibpS6pZnr6AdYAZdwD+QKrfud0YRYCRarrINnavR9ggbHDr
osO1zR6JieJKBuaZVrmkWh0J4+la3l25+P2exo6qydgoT+QbraKZa9XB4AkhUQIrD8QaCRfA5aNu
UDAvggP19r/pC16LV4+yMuiTYIkqxzOLaChWtZXPGFEgOd59+wwfpE9Pft2rFffTNfSMdzbKlt/g
R5E2w50tvK2cragYKmT/YVhnqny/8PPQtnf9GWc3wzgaL5LHNsTXv8TuJx0HUkvqg0zUNdH5YEWo
PjZOlRn76JgXK7cYS4FEjuFjG+zsQjvmm3gZOGcvXQVUsWvF9u4C4BKuROZ3OOQuIxfrCeEens0g
QXMlI2+KhD+J1F9Ok7EKyzf44FgkHtO0a9S9gSnyrX5RrT/bGx+p0Kd9obLylIEjs6PIFysef9Ca
hxOZkEaRzLm/yidC+cTyzYr7UQ6OR1IvE8Er0/xLxJYzoGS71RxaeJerja7lBCkhtl9dGmut//J+
TExp63Wm6WKlLl54h+oB4AgWFApnRWDcjfCyL3qKCBb2pFVsUiG9t56txVxsJ/5BvArvdmNlsm+d
U+iMSZFikifRdYTT4iw2/USDPpEukxBkxiAje0PVti68hyOHNN9aDsgVrjH4mpoRjaksvkp5Mpvm
a2ckV13T1m3KZiA9Co1EEyp+NIV6ql/CWstsfPdVuncq5Q2pkwZPJGNV7wOhMc8QIGYA5lYOa4rN
HGG8xlGiRB7iXWPLjvcCs/xkJCaBHCKj/AnDOPuHdDKBSR11vSN0euBsO7hs5gRFsBiVFC1ISsvZ
JXKmzAjki+ROKaJ0BUF7e/ebZf6Hv97ZW/Ql+SL5WFL1ML6UeRnloqn25IBA8tIE8JlGTjwamqQd
Ecsr+RftcjluzEEnotDDrNTTA75S97AJ/o1Mkt8QPWLYY4vxL48aNG2bk3ta+U+7AMpYWJWS2UJV
Cxe1epl9CzgF3nM2MRY+gqmd9zvbAczHIkTs2J0y3pA7NU+N8qC/YzJ1TY08ykD2PdWwebT8zGY3
lyQRxl89gKOIKq9vdt11KvnIeXqTnr/uKIBO/J3x3PnZc7AMlm+lIk9EH6mJ8bXClxGwPb5YLTm+
vqM0ClTGh1kvb2YzlNJu9XX09mKRSGVYrixoR3UU9TMJJXNBtOkQrMw5Eo4QGL/CtyWVEGm1I539
9Aa8A0Y19N4kbcDuOGUX+Upo2TdtWoAjXxn+duvogyHLEOjsGo/ZCLgtDTBIyg2/KHPv5Fws0Hqj
HdVY3z9t9O8ItqKeUbKgzuXv7bJn5qlT3E/hAIUYI9qpdxsSgjO8/TfMHfJwjr2XnJpF9NsShYXl
QXoMToVDHeZBshtKQaAYgiZY/chkg9xR+ZNyAxj9dHND5kWP2xGfM4KLs5PyNhNlcNCOItjOC50p
1aJm1e4b7qoQcbA3ISimVEvjRUQRvZIYpAZ7M3wI6Kh16nGzi9mFiHcVsGsmYZGGy65SU+l9lVEj
XiB5Fhbos8CU+N1ymTiCRpo6Z8s6FQb/K9h+a1ZNWNRPIpYvfyJQOANAG82NBGYrCkm0QzqOaXAP
eoPh7ad8cqMpbBcc4vA2CNb6ZdObKAbPzqCW23JA26kf4wwwRuCcb62RgpC24G+wNqyHG3z3zte9
QBeqCfkM6QSrte6bKgCGFdI8jjX6BrZoLEW2W4ToYH4l9R7IsdnhbgE6m/I3FehA5u1ScKOb+Qoc
gblLZGxu27149QwPSiWbHbSVCKN6OB3lYbG0d/g+fRzxNjPs7KqlaHkLMSWB1CvMNwYU0Cngb0zB
iggQhx5WmCjAHD9NDQpVsMTFdR6aqCD0xjY4b4ILO9VB+JcTgrZwzEM8TKISf9ecERYi/TrHY94f
NYyF9rfyMJUWXfR9miuxk5uURZQwEf7dgU6k33Gix4bL5WWIi0qcTniN/KM01BHBnPvtU32/8ne2
DWVoVwC9IXENiSDPWyvxCqVk5D5MJdGf1VIiIeC7h424p/n97Ww30kBJvfEM1dL6WZsQJzKg1+qr
uCLFzoKr44rogwXDIrrWidlCWHX66tu2uhg+r2qvBKCxAVJVW+PiESNhu8m0xIfAAEW683N9QUy4
iTPSaWI47vNPKSBr1fgnJieABKTG17h4+rivJ9Oazet2POcs8i2ny+Sp+iCE5n+5MqDT9kV6weEr
Ce2MC3O3U1/JOls+lAwGVnuDcS53doUF8q6+6TDoWSckr++yszwikIVvsMkJp13+TqAuhwNM4oO1
NAIZG4j6NFzrRW8gCuWvBiMAgG43ZIfe/G/QF+S5joRxPyfSJ8VTTT6ahfi7jfco+YCDqsaFxegN
f1+N0ZnDY2mK0wj+hpigBWLI7PXVnAJpFVJ70LVKQ7H8GXqrfiH/oAZqaogGvetBrUwSfxyhLjik
eNnK0gZ7itZyZdid0PmbZ1n3auSa5QLK8KEbQ7NXSTfTQ403p/ZWqMKO0byy3PEjkEQNswIZvQot
WsfnRKl3EmkUN3JoGwVglIsKW722diplgwssv8YNu90Cy4DjJuaOOqPvPiC0srPkk8FDLUoleQ9P
O5Q7JMDJr5wl733ceWBNXgvN0r++SbdBO7+S8aiImtx6iW2Ea3B/ZvpkERGj2MSRwqOqkilE0l2i
ZdI4mbzZowqCwwUieAE7qkbhaGRYmJfvPubm4Mp1rD3E8+4pCX46jtIeLSYWvtmLhkthq4an3gPL
xzAtrFG9f9jdbZZHC4lA7Mr1TZL3oB5bz6k9Wxx54Ht+1pYwhKBYt0AlSPeRm/z2FXuAsbeMZFh2
7dRaCTbhL3QHYV/VakOlXqXItnlE4ECKsKIxUfNNKU8r4+9VojiE6XZQTnw+eSeQd4OFSFCno91J
NktfWqO3h8wlgnjhYvxlYFwpAc5zb2KuyZ/IegljtO7ynKNVIcov5eBMBQxoRh/NUyUNoZtc4arB
YHb/FygeoyCG4WyBv2WRxtQSUmGfoeRyDIWc1YhhNDuAiJYxBxfNyUwT5JeMNzBVN9J1eCKJRgRG
rYm9D6v+v6PCM72rJ6rpMa37H9w6XtmPWS/68BN9Qi+dVzBBmHGAEm553zC0GZ6D82QdjWJkoJIb
bE32G5y0cTa4aba1Zx5kx1sLcMfuItk8KYR3j/6TE6enjPfJB3fKVhU4tTgc12BFNYZldzqdNQeG
01P+mnvjlX9o/lh7gNHUlQ9/tHxHRhGhiuKGg8stNFuWxcpOXVHVgVz4brLoSY3DO1OpdjR69Vam
ehu/J7w11sEi1Dnf4NOPHQvXuK5qFhI1QGOvuSzMmMw8D8Vi3pQm2r7GcOrFEsGcUSbl6kwaytTE
W7kPzlHivVKDjLCy3jq68wFRfARQq7h43x3grl37e3F9YjsKRXkpbtK/wJAPnwz81IQIpFvX+riG
kDJs8ZnbuNbOXZw5b0jYxiog3TfkV2E58y2v8IKZu6mxnA7EnlNgGN2VrPjBBRdqry0F5q8RR3h5
kWtXzgiQjN2aTIEDeZ5bKhHtH56SOllnSlczyVFXV935WXoHGymcIH3Xt8edWswhCfZ9/GwA45Ns
7Z8kv8mIf3OEU8MYOcbxfkg+mGpEjU2Yd5ByOU6ohFKjKcauqPe+vn+vMPG7/4Tt4NuJzKkx7wHe
VPDQrGFfWLgplsLc61XePYqMtzo0L4LaNW1TIlWEwGfhEMZznIqc9hqL07c23Qs2IM0UcWB11+20
R3eQGpFp90f/lOVK2Pzz2zVKmKapkAlYvqo1/a+4dwuj/a8YlIMt8IOjnFM+mzJ/J+oqI7Y9GR4B
Rmbd2IUDo2Mli3CT5UuPMNZrG+mnA1gu+nStH8TuDvy3piB0ltShDhNf7sR6qw1a/pjJQg6u0TCe
pLQWZikkeHEopY6W2/fiHlk7qEkmP8G2utmnqLbgmw+6LOhkbRlgYuwpOU0CL8/gSgjbFjjjgyWF
c+Y1yBBtvAWXB8SlFQC6+MPcLfrUbZ+hDsIuDS6eNGb3/SOalBDM3FFKPLXLU9ByNa7Wh6F1JnjX
EWXWxywo8esAFJXD+bIkyRH4yxSyXjJjrC/gKlZ5RKxuMNrG3CVMv1xj1ptaTnuRPMw7A0Yg6/fV
wo8vRDG3olcdUmCszRBaldOMbKc9bz/0ShYsJ5Xd1QtxxNwFy4hv8+CpW8ZE7Dq6nC6vZs0FR10f
OkGnYFUpHxxMJlzSY2TTp6TA6xQl+UlMt8XbiQIF8zSp82iexaQl9A9Y1kvYIwB2reD/QhE4xz+6
ZYQW2bSA/4SuM2x3zca+XtgHtIsM6O5STczfaaB3GcR5SsfeEc0ap3TB90jJJGSxcPhIGyPRxxn8
b4murYm3ax0dWxwH4oTnlRJslIRXmgW2V2W1kNGRkEJpQO6QOY5uihatZeT66hx+NJChXMBwAQ/l
cySIPE1t2HQjFPvEQei0URI8C7wj9DqV1aZvMUGMIFD1Y8ZWRoVbSDtS6vYSCOrSPj/97nQzkNC9
IKupZ2KdHngnxk+fAiap+HajSNbB0K6IxrUfR92R/ePT6uszAXxLI0MmqC5oShRJSmJC5KhslCg3
YK/Y33BtdQPEVlH5+kC8jmb9xM2WSVh1Z3fzn0wjlvncKCd1GosXGhwzrDvGg8B/n8x3Y2JvFKdR
uXnF0fmXZHXahdwX0BJgPdRvWqnvGu/z3Y7eLqhiKXl/P9HFdKfylBDxSnJbSaTXgcs4oIDaUHNU
4FvwcU3EriboXoDBZfvbTV4nzJX/Fi8NLrVVo/DieghTDgPSSjLfvvRrZxF71s1BUpEFEzBUrAdc
AOm5T0ryv+JQVMulpGvXkdUSl6/s0O8WEfw53oLpfBLKu5E6MaKFBj035uGqzKraSWphptr63lar
KwyFp5WqKRHA9+B5zArZ7c717cqWCfDoB+qCZEN9MhvMJEFMcUx096a7GnCCzbkTETDi4HxJ7GDf
CJtdKgpwPNw9B6SmLvuqeqb73bb+OVXlwVOx+TfQYUU5qhjNpjTbQ+b3Yb9vZb/AHkXNXLgwtchE
NEDMh6ZGwa4eeuUmGPrlJCrtnZh/z11+TP1uUxAVuz/lmNJNWoVYWptLFzueVETLhNUKToq8HwNj
cADAZa2fOfU+KWrYa0MFKkbq2ALdzqXMiuqqcEWwCwU9siKeY7zxLOIwf0TbxvXD11hV1Ba9FY4I
NtUno87STOlBiI2xTpk1p6gZNp3qdic0JVTDc53LbcoqxFKR2xAd/CDzkCJwttxLs/N2djKJgnbr
uHa8Qze4ZfOFijVNMh6nw4RMZz8FeLXmQV2vlVbutL4n7RBXnbNxIsvBr57C1bSesepMLMBfzTsw
KaSymfhY/7VG+aa3TON9o6b9iHVr2X+qhQ9iV4MyNS/YjEGSujiXrA058D76yq6dUgPFhalTZu2b
7o6mrDxspEnXd92vRVnb2BMTyk9E8hmY/Vao1dhWW3ckMvYsVttXcxn8ZX30mQB2309XOXISOOJW
vytc6ILjPrirjGnJcRmgl/Shzrp9kcjUFvZ3xbzcMj0RaQYLnqYmfA0iqo8yuVWAjEcsu2pos0Iu
EhaHGYVDjIF4enfYKNrgnRTVbrkkLraHpkJiIMVXNAyT8+podRDRFmtQAihxUTWxScDoDzs2/AAa
FSBfmYhahZxHzZqfgDMUuK9q37MoQfEioG9vNGbOupoxysf8BAg+pXBStP1nM3HbTXU1j7yupbgD
MuukkAZ8rYwnjSbT8LGdgGx/tYJzqSeNSV/0JxfW3+3HmOvJ0qOlbd1xDiNQ9R0u8yDR5wk48P5g
wrm5UScbYEzHXbF2G8BB/xQRMr6YmLJfBWXx+A52JNrRdwyzM1EUzIkZt0C//6td/y0qJpZST481
607+H/TuZngFlTYdsXBIHLS4u3VQ/F5UV3FmaML7oWg9gW+aAgxPZw6af/KYwXc/oR1yStTarDhC
SoeyfGzl1V/0xuMheKJNjv8quh3Grkf7ijOqHxZUSt4k3CxzmzSQAJqvFfxZwalKPg5/0xkkrJau
9lGWXegfV0DpE8hujvZMsL5krZ7OQ7INVaEQIzVojrVkBg4QJm5D18TYaSsLV63FgM18oQOE05uN
HJLcYR0aOfBoP40xSueqWKIGH4z6gaAxHmvElHbKeo/ZmC1G8ZumBayF/QDykblgnzOldnzdDOSv
sMu6b1L2IIc9KCEWigRE8tFV8PdWHfUJi/IvwvQf5U/mIykjn0Fdy2s9bLz/wSAUDH7vLP3Pc9zn
I3K+gyUbuIP+vSiwtWMxIaGX2UBt/8DGvfmT5eOIFBhIRcxXc8HdG0Go62hSzCk6qb05ZPiphLr1
3V68HhgiprFsvUopEKjrWIybNVQo9ZMQe7dwIhwns+naK87o7U7fr789jSttR+th0S9ePWYwKnSL
YyOIob/7oywkw7hQTjGrMgQUy4IUgPVweOofb2OlpZpbe5A5dYJJE0Lu+gNhp25nkt0LuHvIVNmO
YlV39FOqCPEI8Elf6HoMX+wneE27WjM5Q0CRdbZNkiivI2Mrhm560mgi+GkypENIq6Bcmzu9Mh/S
CY15H8UvNU7dbEAV8Om2zN8MDbr/lZQefZyrK8qycxTHuF7SsKuNep5Nyw27sw/nAW/suTEzXrWY
5Bl+6KhotW2VMqmvjdSmQWCchzbjfG0kLZu+lA3Z5WJbcUUTUSOhbBzGdy29gq5s1gaes+ZExUTf
dIiV6pnUkBUpZXlne9Cv6mMaShdVeBJv/SmYEK8rUPPwVcHh1ELYFtEjo2i0gn2RSL6soXNiskI0
uN7sNKhiOK0buxLePjtjzN+8sHVXy2YRasAoV73mx1Ro9OlDhfPlPSSNyF4yevfqdPg+nn6Uqm8I
pVAkng6dWIc1iP1OC9gUXvMiUewTa4AMNvRgp+qWxcx8QVdFcTvnETAhNxiASJljUtRRXNCs2zgQ
k1pF8yklKCvHQjPsLkZGrlRNSF5kD+JEgwOqK3o9WQRnN24BQVjhPt7yDpPUE/YzZx6Jk6iP3z5G
PkeQaub/XXCS2NbS3ow5MWboQ6QWOLxgO0zzGfaQNCOYyJ5UWN/Z5XXh+KFG+aHHafE1EYGJ+fEF
OcFQclu2eChEonfQyk7TCBt/B1Kxh2CeLE0paYdmVzcQGPX+dWBFuE8wEULoYld+QcRwl3qVV+0A
t7kS9dV1+dCCWrmPbm/Ft4rPJLC6p5NInkaBJ1UuNZoNPsn+Jm7q4xG/ASMAF50b32Vx1Qfz0B0X
1gY4/yFS18qizGwmH2sOZD0W6nzCf6YtLG3JDU05wKtMVJhGjgLx9TuJvkIJ2MKcfQ8GmSVmInTV
DQ9YvnKs9MTZyYWeNKWpJQNlEZ1pWqoz45xGhPhhr/sbFm64Lyj0kBCB+Bm2MQBg+FCaNBvXYB0S
/6BmdYyeK5ag/16jtRdmXdy8pApdTN+sjf7fipCixkm/Kbe3rGRBgoXtkn7yQ/1V0CZwxZ0EcZQ4
n9nABE583YGeqmfAsGhx8MjnyLDKDbQDo1WHb0Q9l6tUXWGzWZt2pYwWWLRpfI0fBhD/+7FcdOTC
BcUjIeVjlinX9XnOEkDk+dynvJpn0K03OSYKcmLWT73gYRwcb7DFjGtPyOydoHJyl1EjtsGRovJD
hMVOWRfC0cgsbg6ooaDZoI465qgLdF/7JRj1h6VsZHpX1B1idsymvdUmP3yFQDF9M9BxBj5Z4PIG
3fy+XMhKdO9GNHOazmpoiUNBdOndekxs/cJlehX/njTsLArCYcdbSqBq6hUUwli9vb823DA+mv6q
2YDH6uiEf1t+9rOdKMV8iEm/pOdN0yAKa2Fj74iRGHJ2ManLSRnFG8GZLBrQ830DSN40wW3NYvp3
2nXdWUhJjvI7ovV+o2LXDPT9URkkJ3HUVfK9Ch7xbPlK8wIvCh/cawj+8Hn50pair5MfuUAwFt9j
dqx0SMYOQBVUr3tGhsuevdtOZCs2rikEn40oimORjD/QAQ9txkn+liEgnMx35Ji21a6pdsi8+BqN
4FHO848RolukBjk5/Fn+j5SsThfVPle367pfxEKrn/KI8UGHYJU21a+be394Y2blxBX7c1Swqttx
RVDGCNNVypyboEqetTUxbELoA6uFs/IJGPGQxcMZU10c0Ub3zmvdqn3N8jCkaUIUsmK+NOqRNa9x
qvPn+Sg1fKamid8MBbVJvBgx/rC5EMm5rIcFXxPSSHECyWr46YxLu20j8FArKH8CPO7Y0aUyGEZt
oxJmJwu6GbY5AItLbcEoa6mvnhZYsq8ymzX+Mh79bNvqaJ08jA1Q83AsPWwEeLKuGwAIlHiWmG2h
DeBNHPJ/jI/yC/pvcjsUJFQsXcmmzY39AFag6i7hhqnETbMccWt8khMFPo38vqmXvncD0PXoqb2D
ubsTS+7nm7KuhHQXp6cHpbf5v8qe4eVm7LbAAhzxmDDkdFjMXPWqd5NFOFTm9as8EsapKlnXVyvF
Sd+fB0T9XinE6tnyokjf8SZOUQXXxrRGkeP9cHtA83P7QQG5ap93NfmiMxGnPWwJKKXtTX2LpuYv
+QAQuMZdCFzi8+riHNGthgfpcMcoORsenyYE0tM4KjlifN7tMdFUQ15K6/EZ2OLphXLN19ZehLJq
dA0vF/J89lCT+CY6eXQDlAb0MEyRidZK0MvbufRrKQG0M4mGNsgnuTB3trlAoN4nXNFQiNWkegRt
mqvS3HmN26yO3oZCf8EAyH4RZ5XjFwaoP79syiSxhAfll6boD9+Um0z8P1uEcrJBFmpuMMpzNud1
Ba+3T+OST8ZEO2QSl+L0hwz+YVQ57S9Zx4rZ45kL1GB//+zUcuzd8cJik/e09Db6X6K6mdQA0eJn
3BLaoimt08E3Xyhez+/e2tWENwieBc4iQswxa2BhNJ5IwYWS3eAUulorYGCmzwAPD4H3AUnBX1Iq
ZG0MZS2bVFrm9TKynWmSgdPI7/bWlpw92Sy8OP3OnpbOz45hM7GOYkfP+3SdwgaRVbORo+t8cVEp
VSFoQrpBAKr1STRC1/a4MJbPm40vtodqdoHG0vA6Dz/S40h5YT53Mdrs8pU9RJakESWOmSXFqPmB
AznBaegWaoUwq5jSeZq+yXd2tU8BdViA95gyUztC04ZHsXLvg3N25G0H3Hc+fIPxA5IxGDsdScMr
D+XdoJoJ4A8O17mafDGB8xQqGymiIvs1o1vSQ3ydKudWON/QKI3vpz39xXBn8SP9xZPKs7iMrQR3
DDkR2QhDA51swyVq7QJEKq84StsQULqf96tvVI/pBcKaSPHbCIuxleCB95ElXd4oRTHvYlAPOV9E
hSMK6if4feuwbADi501YLKkRfBbXwkHdThm/78DmWmW19+h1bFu11MuLJ1T6u1HGyicCDns5BFlv
ogjbAxCuWZJX9x7drspdkEAMRzMCHQTUzabj7lwcmuAnm0EcWEbQ7uNj3xEdcsKmF8FjliYW2tl3
eZyamtR63fuGfzyeiW4cclhw92AOfbmpWd9XjxoPmhkBj/XsJ5om+sM4yscVNlriQxzjiJOaYXwr
DG3dEtEyoAzDEFlZr4WrO7cLEChTiTWMhYCkc5w8xch9uFR3FxmedgcQB2n81isCcmV24k58huW7
pSgmm1fN91ANQLbh6jdYcL8codGEkBIJo2s9v9a9fSGr88FztbfnZeX0La2SPI9f0BtL1wXCgBRs
gRlXMx106sy/fu5+z1RIw9g3WjhcfyQBpRwF9NG5XaGds9BQ6XJz6qdcI86fAZLeD0spkVaEBcdR
mmptsvfkcoG1U5TEA0AVVMNHc9kmDy8xuAH2FDkUsOe16Kj8WzVDbytEKFJRA8hca/TPcHuYUZKX
IC6+OPHHxgNPyBJRYkIlmPiY+Z5Nh+RC2T7UeThqPQwhXA8T1szJxj01/Wa5pVv4nL8h0IVO5Dpj
gPvQ8eyyYPcIQJurKbaF0WlnsQJ9Modpk/zWF2Ai8czOtz7CwT6mWuQVxzLA6AbuPOmwUUI0HVfm
FAcpkFo/rc0B+EFBIdQXiMW+E7htoVOL2TI1WbSApNfnFeLZaAKQ+rlHA9U2+jiGo8xZfk8H/G3/
3KUto7DWjIoJ9ml+mpGe6UKgoxrMrMzhIN6lHftC1RfnG0LkEZvjM6TQIjb5u0oGBVGlicCSlo7i
80u4xP5nqZOTM447zfYHbTf2H98VA4wTy+4s5a2C/iLLGKuo3qzbRVk6hacPU8RnsFuonUj4TCaD
5NN+Q0hE26cSVQSiTqEGDqAcKlb4JZ/1BX+YMsvpHGHgkKhhXh8RPpJwtbr8WhCSSBmsDpO1e8DM
BQfNtgFwnck2aKfUPCOSxRjXKQAp9e5E2vnc24pC/eLYm1uoG0xBTdEa8lVJm/WoFYr3J5wifo8l
7/Yl8GxfcmKx0iSjfJjAf7FLGsZeLXcTIGRwxsM7L0gT1Nb81LEek/s6RPbdmchBSDyGMnJUbRJ9
OhoDnKsMgdvhkdHkdCHCIGlrEKWAsJ7o43fvyJWiXcbbdL92/5ns4K1BxH5b7TFnGvwyxlkOESul
Yi+IKZlkyR8pmUXPiRkjWjrBA5cZ/xtjcqUveuGZGIXuYtA8xXkDQZLBUM+LBLRICopJ6zT3xY3h
dEUUjuCEpjaLUKN2hCTrJHDBKJXpJpKRualpQmRzvyh3pKPufUi0tntTIrDfAo2th9HK4JsOGMV1
SmznBzo3GyeaYx65YZcCwFypdyNbR0x/L/tyDfG/NtPXWE+PvoieVPgkyaD9DUKQXZgSHF3fleFE
EY1MtwdsROwDFObBWGBATWDgLT8SqyaGJANel+6olNQcjxkBHpFDbdgeIMF9o9MtzlZ7vEduLw9r
JPV6+13yS+fnc1KcE12UeWPU7rFjMRRTxTHu6pcUvukiC0eMLU/XSDeRg0YY1FG8eP/zBvc7OcP5
Ssol5ivG1ujW9XEY6Iyr5rvweMBHNaCbc1S+lxcUJVB3bY34aMdspduvQKsJYDu5AArHr2muGwep
gOP0eTHiD1ufdl2/lpgq0Q5BWtEXsSAQ2V5dnQBOJPDrCtdu8HHS95D7zgADZCH36ngrOGSeBp9G
4TQ8aRlcSSHQn05PuvqGs9fu0TYUnLcCjNEsfoUXm+C4zJSiFmcf/7+oXgd1kcXZF7RNITnySaLc
FlTklU3FK1sO8f/PeojIMyUS50tsnGuSxyQAr/ZY3Q1H//J1mi3J+iuhSChJf+H1JIy9dZSbPOD/
L6dQmc+37X33zhJXpoZ7JTotAsR2/ULeVrPfR/Pj78mArauDfx5vZg5250F4BvX4vQfONAaOvnM5
isN2SIK9FJ4KqdOWTSKW45CKtoPEPORECwOEPnEMLvveNJSX2vzhdhJJ1cAndDKut4gmzLB9E/gx
rnNyrjGo3SqIP/HVTlK1X4hneAVvTL4lb0wMsTyLODYPrM3b1n2JLjE14+Q83gVcMcxso3SMCpa9
pOlBNsJU3b2APw614trHK7g4gIMYE44mm8f7u9VKg9Eiv+/tVHDmI+XeTuo2LR2tPuNGmwiiC4l9
jwh1J5XmiqxwLM3iF8SvKVScimJReY0TC0R7H4UXL+Wl4fGjP0VuOXrwXywWKHPgu9ScI3aweRKi
rLz3Bg81NNJekvNub89n9Ex3KohWEXCJsxVNhurjcdatfE/Wz9eTtwty3v1RVa0QZuV9eIFPCAKC
Dq6pDYI9ggmSVLA3EHkfxAK5fvauuhlttigY9IvsKZjeIrSnlzfKa9J1vRKKp/6S4dQJEjVOHtiE
j4aT4kOA59jvFBcOojO5Ro10fJl8rXd7olm8XQy4SxsipkxjnDHBbBZkbfOZwVUGLEEhkKpTvV9F
t4JrtdBytACJlpU2NOeUgruYnxQ/SK543QEG1FSrWYdV+sLVVtk7t+SDyPfM12Ym2UAbSAHDPthG
3Rk/j0dUv9+miZif8PjhlSKq7W2D3WoFV0HBEuctfdfL58OcCPrxc03cpw2Fz/loaUVw9u6f6pvu
Rlwor7exd7DcWGQ8ujgjJC80Fk+JbbfB0lVpYMPXRsUBSaLdSmZRZn75sIt10ppywDI/O4lLT8iv
ZuLGj8fL4nLLoTXiU3KZSXu46qz4r/jbrlAbeUjXpvzhc5tMh1e7591GkjvNv9RtIYIXuPbCnHvM
tShEFM6zO58YqMACEpZnoD2f1TW0amadnYNVBtkEn9jCiZ+qbKi9I7mi1DSuW05XknvfBVgzlgwx
yX0sW/oYUEiL7vGnGgRh2sTky9pdcG6kutk8/DMHdOJ2rZbeczgxTcEsLIKSCkw1PsVp7Anskx/N
GLjhvWkaxP7w5DaCi0UOxOsi4l5AZsRPVHf0wO2uLvzrXID9j1noExPpgjhtMinwoDlBWFkL7d5p
acT++dL9ahxzAdlp9Bljm/bYJAr1K7ylDaRU0zXF/elbooUACNqy6DkLLj3DN5QFBljt5sMHtlQn
Bg7K5m7MFUNVjtF92oe0OhHP/5Zd5S0FXEqn4Y7AKNpmmR+a/rxuJWtpGg13vcvgcprFJXu+Y/sQ
ofhaTcP0Yau9Iu24krQkVLS6m8FYVTfxmqNhuTwAtryP8WPbpBLAhF79upb3mI5QQTcOzNWfs9Bf
qzoR/2wDf3nYdYiEm/S2qFSXMIuZbodpiLhCVpKAgv8tAMweTWZN3PFEjh+rpWNghJOtAR59mTH8
drFNkCUI6ziO8QeW4a4puq/O+0DJUEOjiyEWnY2DbvOFZrKyL1Mn2nvJg9iuZF8RqObq154xeogC
MdYxkuijoEPn+V/8zte/iYQJLU29CJPc07E/1QUR8GrX7j5QJ4fmOApCU8ThQ4/h/pdEbMr224bN
9hmw9tUvXus5Q38O73DXsEaxhx2GOJ2IBXk31pDAL0IW5O/FCwHZIKrRztByB2mmGOZLH5ne/Ese
pLeajcKw6D6hID25nnlpglLqClrYcsbFHKhLN+XHbtH9ya9eWSrmFDydLA6ZsvgzR6yRgyioc2oT
q/5H9VCsB1EQUf0HAxt3FkdwhAgu9KjKKIoj3+SLmmZbqOO4gO+ngzOGIGdLURoDaGsowvGvmzLi
F9e+TDVrA1qxNnaIlwnJywRlnbw4YkrcqmrjX1681srADTQr60aGOiDyT+1moUdytVx1rM/Z7uPh
d5gCW0JoEhE0iArq5tshozoU9Z+lswxKIeMv4r++6Hee7xakMqqiM+6RH8wRxVHheCPjpRad7Aqq
dHYLt70DbxLiaz893yU+5nvklJ0WYfaVOeUQ4i50lwxlehckT7vPOfSRiRxbt4A4xQiVAYe/8ZyV
0L4KYpRnxG/9IilwXJnRtambwpWhi1Yb+6Ogvgly1vuy+UybuycwgkmxAs6/oEZweYfOzb+Zuh5t
eLBus2RBPhvtXzRjOQvA2+IsJRWVqlKJAStwzsHip7iqvMWq44dCAzPuX/MM2DZz+F1Uau+koGMQ
7elgyL6+8LGjdmcgXH1h6j9m3B2vZ2O9nAZzPm1FDFyiGYMfa9nwgPzUldx2NFsRHPmAW52zJjq+
tdApTwBwGsq/OQcyWEe70oxLuPKPUKNlO8Uc7yNPlHS5J7jQgL3IfsnxlJ98eX/9HTAeNyD4faRu
v818le+nQBnui7v9lxyZytNfXsah8IoStJcJ0qXes9xQ5yIGMa0Tx0JjLlqbmhswocMOHHSEoAny
g9yCjP3ACDeq+dtG3225B3hEv1HlC0U9WwsRrj64Q0JpUC4RSWO1bpMgbeoTliyNMkNEwc3bgCm3
HbcjhaM/LP/PT2sfvd8z8m04KiQeXHUJnqZ2wQ9RqQPXMM/nfa33iDgyumOxZGamlE7OGSVgdcEe
JsNio3Te9IlOzm00xG7OaBMJ8tR+cyyjyU4dwPFEk7r4l9o3bXbJk6JPIz2D/aQEAFhAENSF3JTp
rh/c/89U2BWMa67TKMs27TIYfzvm+yAvLeoG/AIhsiYoj7RtWcOblz5zXXCFb1VxI01eUfnM2HEA
986TzgmTKFYGJ/RIb/pQoU5pFFqcDnauYNLFJAdzOObYQpKLo0MJAZnYrEQ7Rf4jJNuInA705iJ6
SB8VPgVchObzHX3tNdnMC97qp+ednhRuUAHlZyJekbVVj3FLKSdCAn65ZKuF/ZexrncHvt/Sx01Z
i/ytt+0BnQlxLZDFV1bpXOezQXYKT32mRiB0BgFS7mzY9EdebW0ioGsLL2a81qynH1F4mf4sNSBB
Z0wlYk/jo+t1gMnKjN8vNpIJzXjYjtj67q5Xh27zYagEByyyaN+f4dKaZrsej20KtCAo3rmDKrak
yNzdq5VNeA8mmjctz6MjoyURlhVqYhx+E+SzIDsIcD7d4kHX0fYvtiF55EjXNRlNC1ZEwN6h4btp
KgaSv+75E8bgVvNfmyTM3DzHYCPj+COGHLcv4IhOA4iRbrgAeJVlOQcaU+ZMlKOAu2Kv6GynKDx7
rxwWhVsic4GB1w+aXY5qWtBT5atfKuE2VxMAuYFoNyqBrQ2KRfmFQljWBjtr62BbC3oCR6tSO4/n
IHmbL6/iNHxbA4/xDPrmt6xWNgCdyGbNb2K7OxkKpiiVhXWB3gUch8xtiWxGsY5gpE4WAYg64SLM
AZdUyxKyIMNFiozufAY0HBzbqwq/wfz2FP2+5yJMTFNdGbwqoM2LB2oAGUbXp0xtMlazmMu/RM2M
rTHRhO9e4RFkrjlmVyGnmx2faqeQJk/A2S6LPMM8lFqWR53EkbLmmjjCHoaGFyzOitMpKyenROog
IBb0jUZp7PHnLxzX3OArDwyonVhBhldaVObs7lw5jBJk/2RfRhus5YA/fJrYN9JWMzm6Ge/ixi8y
EPQU8jgJib77JXxZwJUIxllYf1t42D2RDOR96F0WwtUFCyMRSKKwU9Sj6HY0gJOf/LCKpd/8qV8z
5kB/z8ZGjTovhjmB8kQmpRt5sRwB1NH5Z9hGLMd71thOzAeQ+3rKE96q1ra9y+8nYICt53JQkdP8
34EwGqUDk13Ms99EeyZDG7NsWRCpIlNUY6+U32ZJ+7QzPccmZQGtit4kyfsV/324rCVmOeXouz3J
rohmhq9YOqToJnv99ejV+2V82+XthJ60cu0laJjKU9mUWjUOlD0zEzS+RCgtT3IcvowqEOKppSju
VvrAOXJVJwtp2u4S791MGCsHHY5Of827me1WSnq5yF+OC/WHKeqJFiWXg5Ru+bQHnTeXfJ/XWpl+
GxTj6bX6UcG2um0STaVD4D/kaTk3PbCqnZwuV9GdGVSFjhOw5GSwONeDcegz87Ws1uOjH3yKLCq9
xR127a/tLjkJMtjVq/gs8gB1a94lEQplx5DbN2QW/J9vGHGtcN7nFD8yvQ/Y/X42rP20Y4nSX1rn
iQg9ehPT1XCI3UixMrKtORPjIUBBPtiCQyawxqEmzyj2vfkyv7cOiPRzWf7ff0n4XMS9B+NS81QP
8UfEZDco73TMc5tPL3iKduOaVguiTFtJjaVpwCp69tEeqyTxAgcKhXn3MVZ1Ed7+9XTC+Z7nlT+l
tqmdkVjmm+nZndgM9hWtB2ASTILQ7qKwBsk+9beGlZQJi5XQ/CSLTf6oVlrYMDKS2KBkyp8dTJfA
Wnaru7Id94by8W5B/tgsPrp8yrB4NKpbBTGOwXp/vLpKaU9SBgpN26aSjAzrQEi+IyMh9zxpHyTc
Q53JFzXhnWTjvT7+3CqMBsCF5/rcdofzZXnzKWLShr/2wAWxffPSq2xXOjc180Ytn0idWMqsZXRo
zDOAur/WAG0VXGYfnMDZAukk5zZsy0yXXuXKL77hH3eL6pVtvlw9dUwDeV3sWuIxHvbPe9vBz33R
Csc6gwUSe4/TXV1tNPaz06bxL1j1BuLYvJWWP2adiophiwcy6KIWWw+a/mrYfq5y2IQ8mwprXHqU
d+sU8/xejxh1qJaCTVXEqAyxJE/tWhK19RY5RzANjr5pGOOfih43xdU50LvyiUMtW3u08i/qvb9w
dMPEa794K2tITAcHzjZreQQya5I/Dh+BSnvGQld5ATiTclFDUARY5adUSa1YnMaPBePc/DbGRelx
96EnrCI/0PgvUM2v0ONlPwF5mmGHrDYVvOzCDVP95+hobOeDsCBvQiTxaRiotDIzjoKglP+co4/b
OD4E1WbzEIfKNau8KtgufkB+nD9KddRpT3/ZEvJSP4kf59YUE55GkA3NDYjjcvdas2RrMqs+/u53
VRALr9EnpYqifM9J7JeKhnXLvnnH353Uoy8fhwm2LEwyX0nQETj0S2frkKf7f+bYQeLfEDHwKjew
s83Wp1Jz2w5kggOcxi49aPY93ewq/NfkZnDBhjA20lOqkBr3U4GhlTVnZhkCjal6LJDGLfVh+kBo
7GXUgAcSRYYgv2IqJ29TYkrjpwjWiF+NsPqY3wj+J2qGR6y0+/JM76nOQU2c49qWaCfQXKufUlUp
7HWp0/tbM3YBvF2jpA6NrrZ8D3+JEsgWDdSx1vie7Tn+aqkSaL5XRRQjXn1vXo1YfO9ScSlC0pTG
8hIyvXfk6vewCEBMj5Tse2YhhF1AjVN23P08MlRJMpGYAI1oI8B72TUW9PdE0SP/xrmzdmZZyybl
52SEh90KGR1n45L+ezZutJZe2jXh9DXxSuL1OTeXqNEFsqNxAuS6E8v9sLWEs/r1E5iniQjjbglD
eUeX81p6Q2SWbjhw/bx4cKvJRPxEYzWuBoTloMQI4Szry+hMW5jMVdhRzD7bg0ifu/SP1Z29T8sl
7fTqrfLYqxGwXIETeDX5H3MwYimZM0FWt/lAUtp1ug9OWBwkQeTH0znMy/orVs2mnUGpD1sbERr6
u237MDoQzBHlYvRPaLW+CulhgYV2PAeiNHh/v7r1o1kxFlXPaGpCO/OFRO8rfivgp1WzqcDhuizc
7ks5GombYkDeLh2fYvm4H2kOl8CN67aiK+8bYxM7a0nhsyGBjAdXSRMPkIlMRfcPaFk53Mog+W8t
6bXeXe372VQZbM6jA4WjJKSc6S2iWK3dumPzmuMQPLMEvMIPJpJBR/t+c4+W+Pk154Y043+copXd
3NeZLeKKG6bpAACaYljyI+vPSSeLmBwjHx0CbwHPrquIuw5KO1Ia8m5hG/JYFfFf+m8mVdCa8Xo0
IuuK8LNgD6XP/QOxQNMSXBbrkNNNfxGwwAcfEHDQUxE13AIyYnfAJ15Cotkc0qAXhzshoqoZDa1m
fT9vmM7JS8tijbIpRCMj9ft7fwoGIrtdkQWmXo9W4ihS1tYjGlgDD1U4OeNXVzmd/jnUfUwcmI+y
8BrWzgcohRq3UZjYxXuJ4Q6iJhugsQs7x2G5iWn9oT/Ivk+sbjIKEhjVGopHJbHsqF9KNFtsYMU9
As3VZjBPDjk6b7aD5aUD/aD8OYb2DFxHLpMlgNXCb9BiC1H7CWCCZPG4e+g1mOOLAlIn3/ZR/EPj
Q+FS0A45n6yXYKw5TftYftxgVVzXqWz/WkT/zTi6wZ+qEKewQ3sHICLSl/U+HMx/aDplbyVxysAW
78331UQFKpjTTmIafqULByLi5CNbNvBGCfmPsgHEmF810Jtt8C9ljKO5rvCjv3pWNBOOVV+7PoV8
yp+P553Hszd/MYsVdsFjGwXbQv1z6DKiKFGx5MDllQpVlzmAr9QkECHgsOqrO6IRx4EZSjV1WcwD
b6gEJ/b2phed1QCHmJgjay/t63haa0pdvbXnq+g54ggaa2DHVr35+xAiKdAWGYMN+EDXKZICsztO
ZgrXG6wmGV08Ba8BI3IE/fl4H63CvOF0oBqyNZjxc8DE2emkaZKjGozD98IneDmyvGY52lBz2uqF
7w/TcL+li1IneP0VvU+k9afjbHi9DbHw5fitcvdqBK8YT6svNYzHkWpHwB+MWLSsfg1LmvBme3Pv
NQ5U3MFrhGHR2HQcLqhwv3iDzyakws66MHd/XjAKOHhadwubXwy+p04tKJtL9yb0Pz7g6PS6b2hO
jU/sOHz8hAsN69LdXq3he8pI2eq3wyGxqGWeUdDPqigqtMQrCJObbQViglvs18JN/+W99ykCoTpJ
RBc40kKx+/xSFJCIG0Q4WI0nE0r6yvzwKcAqKQN16JGLsOuUzw2NteCn24Wpy3PsE8Giy7KycFwx
I1rMZVSH3kuYcaSdYy8iBZZUrcQ++m9xUsVqQ5cOi8jnGikQP1PIwwoVZNqQsagtQWU/fqdgr/oK
qH4nF1IqWJHtbgvWo237w2O5N/84jC/OLuPwlkXXsv+RLjy4Fk9a+78Xjch+m3t4rOPvTxzv+qHW
pCJ48yE6z/tk23dCX2EN/Q9fz1LAbcxh8SBsRY2FQnR4f4S3yps9y29mE4wx6dL0eovuOQONuZDc
82Qroh1vAUMCVy6lNYkCanJ8+VnyGjm5+qm4PJqELI4tPoIWqagxLhK0UJz0hbZ4VN/iwkwPNzlt
d01aqLxv2vrCyCJPSFM1wnsGIJHs97zOEJEztG9oNDSw/y6TQcms/ZIocD1bPJNgszvue6ISRI4G
bgODEnLhkvN/Pi92u6Es1+s2dORZOqCzNDehVmOe5vM/jjd9759yqiKQgQh1lzEX3+PGjyD8pQnU
2E5VP6m56+MwlQm6DLcjK7vTdg9MUDJTGoE4/HljOvm7lP0S20tp2TaCDB7zOZGJmgm2l3CeQ7Rw
taf/hXDG2msSwRnVoJy9hGgjr6SU5w3C7StzYplfYpPHYwDWli1BTclebtdzoUhpb3bDKibdBlC6
XlTMcAxHQe7l/Zl+u5xCaNeZsaZhKiEm+OQICronVfTRJWlUzEWLUb8od1l286bzP2CsXiyPfJ67
QUr7FwOxVPK+JPp0DN7eaGbiwF1HocYwLmEiwV/e1KxmGrl9GbwlH3vMi3w/1XrOC8x6fD7bEnLB
vfGSfQYCNnLdwJNmrWHgq6oOzEEuwpzfELuORLYVSRiEzOHUCKHdq6jJQzBbhx4dMA7Etz7/2jiY
y1qu6eEPzx5vw9xD3h6Lgf6PaKO+lTxzhssB0zZzH0MeFf1fZrgLQqYQ5u9Qo2wdLkpDiMknzjb2
wseK2C8x3qhiI6IsdubvGO7ttVtk+v9P6jaEJYfxmiv3bTiTZrUZk9uDwJ54pHR0Cll1fUXaoSv/
9fZfSg+aNodi3fHInuSVZVn/viysERr7i0ymXWiBBYk4RsNKWdLDccGpB40pNHzXWmj0ue5J+rXN
9cK36omaa3+aLe5hz7wW0Ua6/BFii9n1c/5cM2kqsiUOOOE/BmwECktYvPiKpSmcviXeEdZCwynW
VQIvZRElFC/SvZkrbfGG4Ezjd5p5QCBOa1T7YQ+UZz19NRa3HqP4cTgbPAjiV0yAepvxX4s3fnG/
Nc+hyTFk7jAG+JODmLQsW63QZJdtfPdr1L4WarZVSqnGGAlfZG9Z9MDWIaBgC3povLMOfyoEqF0m
S7QBIKkuZ+rMdh83cG+cfHn9O/b1rCoTsn/Gra2Qd11z4iqTY4mSYISPv+qbDm3ClWM+NxMh6E2E
Sfz+/J6QHPUYvetJQ7awun3hvneXXGYVBkfD4c4aqccPIWTBnz6hZR7oS5+4U26GZ1gR18Y6nVLW
DHxmKm/ID9V1Huwi6NiE3sElIaoxxwuYSgHQZexM0v5E1jVxotYm2dFPCAMXwdG0BXiUkFMDzSGD
xuZ2bVp6+wdfmPN5wsK9em47divaJJSlF/Y+HsZUVefPFA6jMcgUEvBiiGYlVWnuqyifdpvVbb1a
25PyN0mrpp/+8XNim976gQJcW2FgdHTNfKUCVklhJ/ChjCnnIPUk8W2MklgyQVQfVu8M/aD9OtfA
+BgxTIa47FrEnM7cTy8ULs7MRJz1efqOAgWMRjW7ArfgVC9+zKfP/TRH6JwFSwDlcUBaqeiRY78l
8mZr8X/kRJAfxdBu7/mJAy/VLa+NMyUOBBEIfU69yrPL+B37i8POgmpFGD+YN14ljx3+1o6mlsvj
IkVuqTDROFOOEYNRiJNy6RBLc8Eb+d33RFip20RvRDk5dcxTdgz1Oesf0bWu73X+vs9vhku8+MXO
ukUrMVOZ3zwh3yCzgemq9u3Sq8Y1A7GgKrdDWc3VLsp9Z9tT443baHgxd+E32cWtd3YR/Z0e8+ye
a6B4YPsvm1JgGRZqyN23gHRzc62oyRfvZfgJbG7i6ZR6lDnsTX8xo6JR4t4cSGKQZl5hvGjdOqFN
YG9mELOaZswF5+IjtSWh1lIsPoyuv3G/z5xMLsbenU4HouyuaGqBORzz/0QtLuPGvUCsrzW/XtBO
D3BiDucCIvfu1Z3wU5VrDyqL56Kq2TUGisBCMgcl+g21wGlmAEpy0Yk+2+VGwv5hipOPNbIfg9uo
JlamFEJ6Bh+tGQwSDKZ9UtwfXZ6HvqX37aANuXcrSpOeJZMcJGe/d6o+Q2qvmVE/GxqjHKIB324x
z90+eSBe6qbHLLvbcvnxxSkXpoahKCwKdvZLIXVOcxSYpssr8ZppDU8BytiCtWVEE1LT8f7R2yGI
FqxuXBBv86BfBBaEgOR3lIM1PpBQ0fDvNh/oJ8ZFWnzz1pC4oajgTEJLUhObEzQnvmnzPCoyllLD
WnGqeeTVZvdikBLGiPcUGBTGadLncMgF2bIFeU0EtY/ffhd99OKlZnnlgEztvwDy2Be0CJ5kx/5J
0kMbnjQeSW1lRKG1FP1KNnAIsV+aR14uU/aARTxDtigt4BJzbjnIfcp0Uf6aFL+SHt0NZD6G1kct
qk1YUkF1k1gzP6VB9Y9ZVaJOITvmnrz69K1eXri+sdCC0ROBpqO46ofx/iW34eUF+YWfTk/JPE2H
zQ+gH1juxGVX+OFyZKdym5ztpogGl2LsTp6jfPje7UVUhwgHYH1hTFrFxcXjydu2B2Llg/aBwE4F
uJtB6usAn1qEuVu8nEmOnh61cHL1k12HgXFabCf6KhcOk1li1hbi7BJOCv/cObvSkcVyaNdu7ST6
VQHraZPfa2JV4I8C8nemZGtnIlE06VZY2svUKw7JNEY7lCtMoJu5ldDz3K++EYC83m8kJ/RVFyju
lejynbjPJ3kCCIZIlgthidN4nF3WgZTXRTR8aMoml70vpMMXGxcNb26kKNlO61DUyKEskF9OSpb0
bCZBqEGQpoYTe8rvmRoCyHHHV694u5BHPgqqW00eIz0YTXXw/+TDJ1V0uVbBsqteZjwKfmzlBEjM
ei6NsnSI7Vw/71Ly4boxdOQ3hn8LLTM1IiynUcGSSPZ6EUgSz1+1mMXqJHuvmKLTTFfXNLLx2kNN
GuRNMmf47R53LQSR/bFS+268cq9muHSh296U9OScRy+1zXDW9JzQ5STy4T0thOJDChRZPFYKNxyW
Vfvg22kS/mKlqm7Ot7vJu0lJU2cZkDVlWfNKcIQDExgJyB3w+rqY/XeVSmqY4+OAElmC1nXOWSwh
J9frsg1iTc5PSs1ntWjiJELvZ5X4NRcGMSYKSFLrWjMkO7uOJO61dqOpYdt0cnrbiIcpaUHaYPdB
WjSrQkRDzpYm02IX36xd9BhU8+Gb2YS4xPuS3tzexxy6oQ7MysprBTi1ZHvrsaYyciadFzMqSFkn
5OrxSoB8pGHQGemF9bj63FANpJn84S0T3nMSfI6j/9tWUNU0L9/MgLFvVXAA2jSFCCFL71ic4j3f
+kWszJcN4FvTx14Q9dEjKEh45Kyw10bip7RCqHIKF81GuWAh894mplzvR6XjFGaCMpAUoE+FhU/L
z6Vfdh9DCSInrIbcJzmikTBngF+6sisZgy3F6Z2rKkIo+y2HXklvkvRhJjvHmFUBsX/XycdtFB2h
5cXs1//+leXut0+KmCuTidnz7FKiP5WLKnnVDQtxbsGIqp9VrnEip4jsExG/0Bq9OnfZTDgBVkij
H49TmzwBgw7w7d4LOvXCZGYUEAjcgOsYWgex3upolaCr00W96Dc6lmKPZafN5Mwlv36cxtrvEGWn
FWac9o36MyHLbX1wb528yY08wnLCQJA6VOy2I7WtvShrL+mOJODdGcfWSbAN2l+1Lpxb3kjRLuFj
+VPYCZ/6svAjpbylGQFPICHg8HFvg1gEDN68TcJDVk8mYsXXgxnRMI3ltBoq3OFfePQGCQf09gGY
OfC7jmF6TtkpZUxuarYeHyWkAb3Ag5loVtpEZ8GPgiYcguoebVvYHGbYnIVmcnq3i3lDnYAYN1/y
raaLfFRgqGmhKJJymjhqRUUth6oepksIwgWRV1EZGvpzMWa71AqkITGI/fVzqibYT4/7mltmJm3s
SBk5Vy8Nz9AP4ZywFDbpJsmSRgqYZNW9I+7us/slxYQecy6cdUFyA7Ed+QMDWIHsj7Zeia16GeMT
3ryVHERcmzZCkehwYAElIzikt+9y/HIVJCkfvtxlgftoBtYvv/uwuE7mmDFh63Xd+tTuKQRyyE4x
nmwBvV9kinrYDgmmkyRYmmYTZ8BGHmpfscxPKZqUT3wK7cyv4NhpZo5SU6UCYPYaMbK8npO6q+1N
m+13sKzWEwgSY0CJntgFEqgW6ygM9R2/Nskjwn1O2Dd+su6GLntdvXAu0Bn2HzLKMuwiI07VTjAz
06NsTtrQoOn+7VX06SUhZOmxRwUBuBRyDobwBEmPyWLrckMwENtKjuL8z9ZhwcqQkjo8dlGPLCoV
sVSa1pmL5jJEKqnCzJieAgBzeWxCSqwTnHnfMTcDo7aTpWCIEo4okUxdABliXfKyOnuNOCwQHyBR
p9tr0fZUr9FXuV1jwMQ9F0fZVMX6UkaaJfsCRXp/DSqfjTvSjq07qyiWT2Slxjk2Mw5s3YKyQAE0
Uis7/jXU2hBSdiljrohLGpIRZwovjFr4MCOl1kz7yd4ZhiAzXskLc+2KXYW0GsVZs49fP3ymHT3G
FuoLaVLQGsa2tlto2wvPP/ocYr56O/b2FcMGJOq4zGcg9oae4c1dEB52EF2YZ3DAxnqLzFhJKK4e
z6OdYUtZ0qdpcRLAg3uLQaQpjhdOnJHdyo3ZJb+1AvEjWwqLf0f9bX0DXoF9or4rAl+0ymDd74KY
0wKn7GpkX3+OE8XZZLy9ep5r2JAJI1JrRQjm4Wh0WAm9RFCgQuK0Rb8DHjeR4nrmAvbN+stjYOvt
VZCpkG4KufD0lI8XUTW0rjs+hN5PZ14dbORzrdZq6bZdcL8N2We7ga5v252AQUJMfgYjw7M0K1Gm
G3fJGoPuuGJW2gDH2ZwtavqMPvjIvXPnZPlTWGtdUbRNdBtIHU9fBFNZzvbN6vgYeOYfF46Svszf
DTS7N0jFAFTT64Jz7qyecyCGQCN8rREhP9o6l5fTRlAZ3BpJSLJ5w9mFCwGwFthotQ2UWga/cvN8
jIGWAsICA/8jbJmr8m2czizLw8Xw40a9Z72gaKQt4Hkxpck4LZShilxTmplereBwOQZdP13EH8Kz
F6LQj7OMnAni0pxkhe/fS6chTVg67UGtqhpu1gRPEEdZACBiKUEhTHtjaEl+/1Pvtci/ZAdK9pJ3
J8uIoR1ECWlCXJBwNzv0+tbYPj1WEOpG3559XDDlHDq46aj8zzEY4p92aP00DtR68BJ/BKbzIhuR
NOvGoYu6qLyYeVr6jio9kzjEUD7WFtTQtlP1+CCEZZqCiWBp4bdJZ1Qoxrz/yx1OKLNhXuSELCZZ
tL+Aa7QkFRfut4sE/2M6de4s38EQ4J+CoOi3xpcJi2JfVUMAbV5C9AqvADUI5AcIHdALY5Kl9OxM
hmNJMIewabvXdHdx11DHpGa+UOkdUg9UUjHGEgaGUK+IUBhP1us8Edf18zdou0eWpFFbGJiaSfp7
3D4RPcBk2Jv5OvZrgfcvPW5aq8ijRA9zORGkFggUkxAqak/sskagVuC8Tuf3hpsGFJY98la6X8nY
ka/joNVUi9wWFH0g66gBdcKen1OXg1lcyej+WJQtURaekJDPvHZ4IjLfetsiacxryyRNaH17I3HF
tJzkzXNiYNZEMx8nRvaS0E4UZxqPh3/MC4v8ZcaD5Ig6KWquOrNwNDRUKJR1v5FqvbCgAs3U2BMV
ehnQt/4lc4OFueGCDTuoBNjrirFSZsRvUAbkCnQBKaSdCwyvVoR+jQqiT9IcjfPqLs7IaWlH94bS
GgP5T8LdB2IS/IdXg/mf2hCuW+00SYivPNcbhREEfszRWXb77UfOkwjHj01uyg6gg7eGYRDkCkhA
8/7IifGqjHNMETZwsepdZ+19wAbaSlFL00VOd2/d1MkpWjsSQAbVh/wXzr9RsLEXQmi4BJ+fWCct
8JhhPFhLvxmYfYZyyBTtmMQTPHgt8Z8QT0S3mdB5YXz/kcdyevrkkCcOLZjWkdgF7IECR5sH1T4Y
5iQaxwIhiALm0+SQGx0ZqY5lQf8+XPv4dZr7mFE+qLMHGXh6Tl3LMmwHtmNARgdICrTZpHt57euq
3XMyEnDhgyZGl7YAginZmkZDHHYdLVN5Dil7c7LmmMgQG3LWPOwOqxTAShYFutIjJqKIOEY1HE2Z
PoFYG09W8J74FXlzyX1n4ttiJYKVYjB/c/PEnznce+dAH2+QliXLZUQlBLlqquk5B5zkYg4vrWCX
p7vEW2VAP4pN3B5zJNONN61k7SKc9rnt+odvJZYPKwiejvOrHaGtqlj5/Wr8tQHtW2q3HTzFag94
aVdP/3qU4wNYvS4WkqyPvT6T1xfSOwYvEnTNLO+iRCVAVsYBDAxHEjByfSIcwJLoOBkwz8eao1qj
KiELfLF91TubppmBD0CbY6icVlH8NxscabsD6R3qeG7i7D3eQQxUwC1vgr9QRL1rOayJNDZygIRZ
GCzM0Ltpcx0G3citSlC0SpsR68znBFzmytwebtC8cNsX1wj7MapXyKtI428sS10hSsBEi6pkzDP0
RNs35zLqa0BlsWtooBTn7AFqD284AcvObdSZrZmXsCp13KwKjHJ9mxjnFXDH1CzR0HDG6/0hTPDw
3jSjUGM5iiQIMvngW44fZrb9tjSoBCKgKsKpXN2Zq52FQ3aBNh5yG74BO2qBKPNraqpYZrtfmryZ
ZiXwGYdn+T/psW68AUuxGzb4uO0eskrBZ/7b+F0KUYJgWW4oEs53JECx4iNIIpHwj3OYIwUS9eXp
N49Y6u86kIronBNzeBgpv0TjmkJJR7XnkZ68llxTX93U5SePIKhVLONGEMaIs0jCDaRsItlbkKTt
3GQBcZEYgeCEzezKVhVaV38Zqci7DTwBHExtp2VrLtZjotrXqWYHbPV3eOZnGSabdKdAFbE38iMw
c0Gm9wxq99qvDfBh9IEsSlrB9+1jMTciJtsgQQf1uHK77WtMF/P3RVm8ApKOuXl3WugeOqMOi5ew
rh+G1KnfCKIPF/33WAFY1YA4vn1NcD6/haz1f4ll/Eu6+w306CoHbyI1QOaaPlG6qaCtZswGpFDG
KuYMCWbjwaGXXeGxP+CjWMQCSdVXYnxil5RW7CpfriZ7/E5Yh6vQOzW+KxPGIVbtUZKXBEt9yhO+
YYYSopJp3/3Q4uE5xJy3JMaRitRt1MOAWhaFEdh/1pkg7YWoCQWwCVNQ5z7rsBvcegT8/4k7NMhC
/IzNsyWJrM4s0oKJ1/nHfKCd6wLSp0hA0HHqqPnI3eXCkx3ueT4QdfFIfAi8HWIic1Bb6AY0C3xn
Aj6vqCG/JkY8KbiTHXrfpCRfvWvW7FO51mdwbYBoEdJeyMwZ02sBZZz5f4R1TJvuOnB6Lg3eaKMy
/6D+bC258qJPInqjLHfrys7oYJN+4whicELzpbSy5pJEJ0BW69Dr0G+EwROn2mHJrcvduajGMu/S
OTfdv4nBeIx4+XBgXMzsLi0HZYNuxfl+U71wGZD0HiEQUgDjfEYe65av58/F88BgMp/wLrErU8hT
CAfyoeKt+zjoFNWDYkhYgma8Xf3EEzegyoJdOCh0LDqRqfV6lXS4GF+yrRLlQ7Q0iu14uY/oUvpv
ufSi7dhAy9jojvkVzRPWl5OYdMlWGUEYuI8GObE1qpVkn5zJzztOMSo5YzPuTADP+a+grmiv7UDK
G/oRgrs7BraVRY0nXR1AtPzX87nJXP+oniq8UyWeQTw8kJ3+lhkk08/2PJzTk4YXtHWfdqRLQOh2
N81hnGZU97Pj3tvgleVXXnsORn5jKo5VvQq3+oA1fctnpQQCDpp7yKZa0+NkrpsGgP2I+dSguQl3
c2C2Rot91Dw1vrjqukLWnfDxkyTPLZNZ0hUTrIGEAfEMCz75xObwOKdCecy21IACyDJ5GxpNoFLV
TjSDwSOE47fLzaNgX/XJ30+cBXg6EebwVVOQ/Tsn7okTVnV4G7lNa6xXkVvpUe4SkfRn/6OY01Jw
jPtrZdkdVYRKvu5lsiAgnnz61amSGzXQFrIa4rPxMHGhLwKy0+Llz2Lth3pybjtJOVaSDamFbo0I
FDLdew2e/Jl0LC6CcPmSBEJWuJP4qMrJs7UwfHDeoZ48Li3oQ1Z+yA8UsGe42N9sXou4g2r6WpLd
lbQVufwyDtOiG9YNlbcB+V16nEybtVb9QzUbfC6qtwtpxmv/hmtOKQPyzpv7d7qvTKjyoJcl7Ix3
Vfb5Gr09q/b1Is+RCzHISfqDxQZ+wrkqyK1LWiV8n74YRwIfxvpHC0p2IDwESXJ7aal1uI01LuZf
8a7+dtgcOxevIrxhMOkReEZ+Kl6wQfCF30z4ynCshhP/bVTSaNYenpfUdh/nGUtPi+AFw6y/wA8w
/wG1D3E5zbgr51gV8A0rCE9rDmtMUiS2F80aBo3CQ/CJGgIy/NAMlQLbZECcy7K5OLcC5o5bjsXz
PgBi/+EdduWXPDwNuYI623I6OGnLEqBrPhJEmjkW/T+YX9SEHSKqiBpP3JwDFQ9g4gAutLu82rOK
5SjX2hXsdsbvbuKPw3FIr2gyuwD0QB+PIRzJxL5P9oc9Zve6u2VVeWP70VCfMhxObLJ8yGNWbfmd
ouXCugXaGrShwNsJRRNdydpfgBZPxERDrmzLFbyAMZEk8nKG6wPt6izodFf+RvvCK7Xk+iu1ZyMj
W2fNSQocY56qv0gSeJi1XFShHwED+UumvmojncdT6YXuVH3YPe9a/9OytQD1hGSfIR6/cqjJpfpB
1VXRd6sNG2/DiRW9m5Z45GavTf2kUP8DvlEzQADnvUjnh+WRpphtYDhTiBq1GnMItQ2J9gdj8eh2
QPyu9L8UxShRfZyL8/GS/R+XEOM93eAkowjeCTMQjoDJphrvjHM1a6iI/2QLSOeDIJeFDUMRvqw1
vyPwA4x8AWivSteKWADu0z7nrl1w1BkHjeq6RsnPoUuaCBbFZTNWfydidX5ZA7Ks8bQrkAvDIZz9
3RiQ6MVEq0/kDRDcNK4lXqpYPsUqvE8v6zaD7NGTO9n1YdxEdGG1RJuO0RWu1fNrti8owcoWv7N6
3zskPq+eu/hGpu6bDUkvmepdGu4VhnGmayJN0sgXujatPDU1G+W6BNNgpml26rO4aisCxBJ6amhR
7Jc0+X8hLKvtyAMJmS4BDuJ4R2QzEBznBQegMPQYguVNhV6R/7BBSl+fne8MSfSTODavtwebCJBx
Bxj9U/7HeTTMV7u0or9SpJFfFFn2r35DiicMzFoPxJ/qcalLt7cthWeV+1shLy15/gKIAnX3qKNu
p5gFplKwdWfSSd8nXbQ89Rhah3JYXHeI//BfTjiZTVTXqnqRTf/QjRrKSjUFQgpN+0voA/yxyiWU
8wWEfYnF4eWC57WExaPw9wRLH58aZKoor4mLCBnV7tmOXznuOHr91aTP+BSHvsrDPpvdWrwpB2l5
4KDZb8J1O/fcdHXMWvVo88wrMaCqlTwkq/0diO0eOepVQx7mDRFmL51pwZv/niI+eEdZ1+A8QkxH
rkNDMRDUJ39tw3qWcYju6K+ZgBZgwIodjkoQpTspngPBB2JlMwWjnbn4Qeh2ugcFLfM96E3EZlTZ
UX5eGX8Dsoho9MuUDw/1mESb6q/Ui1+fsRFh6FzsIQfYczS3b6LhyK8T6+TL3g+Uco8Cnu2QN9Mq
ZaG/Y2FWUn3YctxOySTqFCDqIFRByNHIMRgEgHVW557kl3ByTRByJovFGnoQ795E8qCu7+dLcGAv
2hbzlXeDL9ygErDSA3l/qjbplTML3uVTKXzL1b4gus/yse3bK0WOVYFL5yjjGkZya7+azvk3t0Jo
GlG4N8CdB9lY9vxnBxjrGdUk92aAUB20mxvlN4zKiGWqNg2JCx1+wa64yocaU+wRD2KZzcy6KaFR
Io+eCnNBRjMM5lbHBmeESk4GF3TPZUB2vFMo0wvF0Rdjma/P37k3v8DIHhdwr7ThCLm85GEaaPDl
vcYKXLfA0JRzmp4DfBQ0HbVFcMkx4+YtzXV4z6aSslK/hvlBh1OVwEwHfBXj4n6CLOfg01tRWKBb
iDkAGsfmZmtGdYiO2bWg6SgXEMwO1YJ4ye2OXgacMS4dN5ccOmLBNBDL/qTnJHTsJn7bM1WwD2L9
eNL+PA/+zGKJoVM7u70TB8WqXLaT6r1MQr8+I6HJdf/AmRnQARj2G5KdGKkEQ3vD3804wLbV5cAy
P6Rq+1d2A9E1G+9DglBnpfYF7Xz65l3avAkYUjjX14dPz/2fMOuy3YCYm87D8cbgBWy9lmnfDUYF
RtcKt/nCoiguN+It78/6o+4F00hj8k1qQAN4NLFFbIAWvyi20A6TxafsS3J60Rn9xpKeT5L8EShq
mkKOgSJFtuVaTHTzqrg9h5OffveF8NNGvz7/ml+XchtHetrzCYZPcU4cVOJElywQb0iUkYAopbsy
oYA8WbmaUnGw3yIG54tJWBXuhjdxohDfma7ZvBpGdtM8Y0OBIoKWiewXyq/0Huqfw+iPV7cQfG2c
WJubiWvR3OfeUodPNUvKgB+W+dDsv+rRR644K96b21yRnLf3pO2tr+G8YeaxbyDYr2aXmbt1AwlX
ZXWcIfI55qP5Z8GKoaR37vnSvDnyis3SimTkmKu2JJvrPwwf7y6li8PGXEygt7TQEqPextmhj0ec
cfdnuyRZck8ZDIaQsrBANcD+EJ7lSNunQ2iGjoXNpAtKI1YS6q0tCVApSBW60irrJ85rdBQ08p/1
QK+LJb3GH0mDO/RT+6iD9BKnHkGoSh2MGgX4Jn/b2D2I1PCes+2sW1zA47/68uYS7fip4rfH0MEV
ikD/e3HNcJEpFEU13jT/1QBCkD3OLjAYTUyknuUgQh2HUO4qm2k2aXSLOEmBZ4vxVQhtM7XrpqhT
v2tCvpUs1PBnjWVne3gVoy5/VirWqQs1RplCiZTgoxV5MweK9F5pOGdz11V6VrVhnFUYDSrH0t0D
AC5J9o0vrVRc9Nh2puNXflUE4o8WPrWUucmb+AIfUGBpM90RKVDLRnRXiqVDPg079bCrF2VuC90w
2pecIS/yGrQe8f91a5U1S2XDjAxtAWQvZGo8dUZ0gke8EQd1znBu2yyubZYnubi6XlIvNQAtNA++
vFWBbxF2tO8vljrDig/cefWuuRv31EA8jvHXISP301BCL8MJjLRnvqTtf47v8TIiiDy96AmjcghM
PxTCCftiWTC0GJPAghwqhD1p8FCfhd6uUKckLaWV/kG8QDPprotcesKHX0PCOUv6F+l/40H04nIX
ifeP4LdtA/ijJpPITL/kRiFW/OzorNbDOYdCY+7jbvUjU8JTi8BGjAga65ZmD4ccVrXhoU7Y/fTG
YdDsgImJ+3tvkQuPb9aHrdvPm1TXufUcs6CBAAl0CBflK0hBNxeOCT+YkCNHQ7mMECFfJJ0AGZUy
WjPEh7P+7IzSpACk2xsyGJbBYLBYbrVvvJS9KLYNu8e/D3TsEM5VqhwKqd/hwtMGuwP0djLap512
6IC/QGUDeHYoTzyk0wGAPa489FDB1gJk/NV+k/H5Kil2f9osZBDj26NlrBzGtoYjzBp+q313IABI
U/afQ1KKP59LQzprqnUVMkYypdnZVCe97Azd+16jFjvzDnVPw4J47HHPpJbFrrPERTRCfxkqUzgR
+3hydwTyPAsxSmi67PZubzMJ7dQaGhOn5cR4BnzqM93//oWi5tK5kyEMlcwQJ2Io4kV5fyPPVaSr
KT1V8b5TMH9+AUaw7BXjdEVJp+3GH7EUvvCbuntl2HdmG8vmNb4px3IUE8kQaKhrkubYji1utlyp
OiETa9DYH7YudtCrpFgrOddoPqE4IPVxU2Af4zXJJz8O3d+/jWF7YvPO8DCbZPAOXv6pqqJ3bk2w
piu2pGYyeLL8h+bj9LlarBrgOIEciVx3odEMWwo67E2cjsP6uxMOOrIr2HiN9xceZDg4JKcOgYnV
oVPasdLcQO+1TUUxE3W3PIc2lipvupZ0G3HEwe/LKEuIpZYt+WmCqZBTMCVzt5C+BNj9wtrvGIMN
88rWFERsb8CIc8xfTqdo8yS0lhw6EtPdUGS9C0QUTWS1Hz2OLx/AVQkeRNtqCJlyhx4Kb7A0M3WH
b1Htd+clhelvcy0xSfc16SVDfElfN3AgtSsz3y1O4gHrkYYZ0JCeKgXpdS5nrUrHXzROKJdRqoF9
y8qXRLEptffnYe6NMnJEXw42plAzJhoOXe9MsNZTJc8bzLSI9Jk0L24mPpEXv3gRrcVRdNMBwjef
kSmZTdMuOlcnlrFqBJFS8/GAxM237bJQqF0dYMq/Kg4UGa4L5lAm783rM4nwWRIK/cX+lNh5G5Ee
KAp46btwj6Mun7NHMHD6DuCio3ueXX8+nod8fHkhXfGyQl0ko/5H57V77CR+zuQ5Q9ZcCFGcOkgS
heWRubtdWSdA7GlXBWPJcBgU11+bKHhjkFtBY7LUD2z5m7jQJhOLHYneCJQMtLOgv8LFZv5UEqrA
2EdIh4/aKcUd8DkLIpzoZT3+OOL1k6yb1aOW3xycmuHY9mu7i9UTo7qKzgoFP2uGtlwawQL8gcMs
aDU4WHvgEHRj8/3RxgVeu6tggUFg4ZevgOb0rjIF0uRWBxdawCJusU9er12uxz4vsSPw37qjqpH2
bzsUTiUg+tt/r/yTV8o7y54sIClVnKBQR5V0Wc7G3HlvjF8/GS+Su82K9mtPYeKNJNgXT+aCfpJ8
flyBszkmq937HEwi/YJ11PLaWZcB1D+J52hTkTHmN801cXF5jm6LU/RDHmRULClukGpLum9eBRr0
uIyuqPRQGI433Kai+n33LP8BsNILZ1fqMBzJkhpXtL5IrsjLUiy24n5KgQsiB0YTfX/Gr+BKI304
VA3DQYHeEkCIpTr0CnbF+OaQ59//oxf+iCqDWKoOisU0pafp9V1fjqkj0q4zxaKUkl8wlzHGGLmO
SrRWcq2pvkdKevTkq0XP29LK6HF9mWEjDrAc4yl3bvNtbriCrbV15PqSTeId6ayCzGjLNEXqq26i
4x288fC6A0dpdcJg0t9XcHHP8MjrnP6gOWQHLiBISWbaZlL2jGRfcpSAiA/61CEOIRN+40rPYEk/
5FeUzdykBvho1G9J1oUk1qJDGdCMzykEhebzXSJ6Q12dbleXcpGyXKNqf09uQk2iaJpKfJQYoY85
DGkh8b8mAYQ6SVZvRX58zhZuM4g+usYyJa1vpSslmmuESeH9G9ZMhhakFiHJK4zo1e5ijeytSaKi
QuLjkzDj6GTZmb2UkZbOuCQbVXw737ABGYGndgSgl6qU2i70yQ6oAJI6v6XW6uV+LSo70i0UMDb+
kaIOe3Ix2Ze59xsazD2vQF0IKYGwK86F4nbVNfKtrz01tw2TgdvDXyac98lBm3ym1Bqe82mRoSU7
4idZCG+AY2CK9SKSKMtY1LsHfodH61LP8JgGjH8eankFJp2m/QCwvOWvt/7E9QajZzyWS3VOGk2S
ROAAWlrM52EH/F+ZdRryP1x7NYaa9k7tcvPXvLtAmXyNAALe6TEPnfoun8ZiOQ03tavfnvn7pgZP
ZrbEpRoNpAsPJlgEd0t6RIiiISUUa4zV831yLN2hdT03qiQxVuxdCbOsuykubqFN9qU53mDQj01p
ER2u/ViZpinza325JqiYZAjVfWnVPoec59hSeoKr/NPSK0ybfF3k50pAlHmJoMyhVdw+6MpGqI28
OEN16sQBXVevHyv7insgHovMamL88hB12GbcnavnyIkWDdWP4hz19f1IwTftzwhpapf60a/t8hGd
/ro9jxTVpXg8mm8HA9GjH0VhWFQonQDhTkA3kYzTUbS4x7XKe+gm+Jr84cB0FrFfLbhpxjUUCu0E
wkMece3f9jeD1Uc5EYkHEnO9ENWAsJ4FxkmQNNNg3GvtL10WgKwraVvSyrgT8vYk+K7p6o4YC3jQ
wpkDiWRe5s/DXaQfke2RbDApDjtlb+2GT2bCug6Dd1Zy21hCcEpVWKgxGAuIIvmfVN5o1dOdgx3e
9PGV8pcWPabh41i+D1rrQ0gvf3UrgMxsnoGOpQdJiHIkSP1YV2PtKj9YfiqoEcIxc2YAzyRlHdBP
LL/BciTWeZfgegbTJKbm80gO+BRLqI8vP+xNXSEIh0tWlGwGSHYsKXC+U1Y5JofsmUFWM2EzZTMX
LnB9N4XWFmfasJ4wQI/ZLZI4WTsUY0esyYI9slrgBckBBp4KZz2W+HHJHgqoLiuozBGAS619VYov
udvHJBESZHKK2VUVFTI3yKZWpqrMVjL9N82AbOA5ZSRZ35M3TQUWyNFG6bOcshzw5k0K8bvwoXOP
6XoZnVBx1E8XvP8h/JR8ZfrP2UPJF0gkEuNindcsUMQOFUUr3VnkKFhQ7ViQbyxOQw/3sS3ICMJa
CcwhQlbPRBYMetjRRLvCHjFMugMSTDe8Jvjif4kvLrGy7zuc14eQE+mueEQaizuKU1fU04pWK5vQ
kQxFD9BKYQw62mppaEypDoUqO8Oju6zhSq81/PHIezGYXZU3QIz2rqdSoZpdcMOP3T0RnYWQaf7A
DwogY2eHaFB7ZiIQhY4bv4H1pS23lUujmcZ8hoMGnm1Nwl/vYeph0qD8YfQIHInH3UZ5kiGPuryb
zojgAsCFrSlodBG6jWtRRFXaE5dk+l7pqWtr9+RPnrEwC11UeNrE39RuWmvsqaqKmPRXtcK5jdFl
bfx/Om8l3T8EUB2NpsZsIEfVPuVYK09hq2Ud7TXH4fXbH5P8CkiSZ2YgD4luuizPnQ7jVfSIvgur
tuXF33vgtog4AcFWPF3dyBQXqTPGO3wxX0pxU4jNLe4f56G+RINDJumNA7+kd8I4z9W3VVpzGU92
Q/+M+2AsXAp+8GEd2IVK2X/8IoNtsJdDzXX4oZ1i59bTlxW0ozlRtJTzVm6VDkvBzQwQ+hHFMhPO
UXtnEuhk2f2RZuxoRq2ciRA9CdIrTPbPt+PTOzTkL9AoQgd+ss8VVbDYraSBDpAkY+k1T9GG4vl2
6tGjLjUdbi+aF3391SlblpHBxfDeZqX5QUJCmqefno2B6TgixfzJE8JP6vdrFiVUwiBw+ku5zh9u
EXvLEx5oddGbIvNN3lf6bqFhiR6eMlEWCwPaiiW7p7Gf16QwaboDO81s1tOondZk7txJTkZss1FS
anqLbL9/fS3/oVssfztc8frndWmG0G7jMrN6nEVKZ5aV0T8gLQP+tvUZ24S77fjlu4euiRDeQ6uE
UzBEXoeZO2O5RbGvvoBpP0LG3sOf9Efaf4XOhntefwBSLmtWPyQIBJwvMDnQPekCbg68R2m+Gfis
SjZGhNHRqZ/2novTuwxqoFkYBzhQ6RJJF7WftkTq4hs5zwiLcrf+L2cyhFXtbDByPrMMWx6pMwsY
9lahr4mA5GYjVU0Jsb9AAf6HONGYl3gx2pJNVebO0Gdq1GK4ZW1bBgI8cbEjRzIYwBKUf0GKsS8X
sMFszf0FJKSDyBYD5YL4iseSz9eFGMgjWuj/vcdEEdv8FpyN7mIQncbkbRRK7WxBcO6xM5AQM49L
CgYAG9sK+ue4UNmINa29oUlkhjbaNm+8X45s4KnyacUHHOfNWRcEcMwMTKBh8X6YApsZPR9R5W5A
TOcE0hJYg3eZeFbj3caE0Gejod1QiIfvU//Yanlh96s2YllTr1r4LgkQv7j5n0sJVlStiSiaNQIO
XEp7kThA5bfjpW2anAXSYQsgSgoWvdEybjLzDuVh2LNr348VApQl+eRVNwJ8w2eP4PMNVnlBS07X
nvLbJIFnEyD2VjlC2Fw8uEkmSABy1t3XDQ1C52gE+cZrYanQy5t46GsL4HogbpLYD930KU9+O7X6
cTZQFzHOn8Tn2hndKtRgfqcM/QhHRw3WDE6ZiORFjM5PJJOXP3HsWqgQWS3YVOTDlqFQOyhtJu4/
E4EG20hRvmIS42EVvDpn8dNB7uUOSxhBiXyOKrOhlpmS2RLJzknew76QSrcVL/UJIPmz4oHkgNr5
sNcrGhKAE9xvMOUQTqlmrkHY8LEQwI1l6tiYzSCES15y3wy7GXwpBPh63AvwVC7Go2Wo7z33999k
9YnRowXdzFpysC3ioDhZWRahwKOD8TuYafGKnOG4GC1MM88rzUCdocBHmoN+4rEw1ZAciZYSI0gn
Q2R0JpBGX4qZMurkITqbnn2EjD0TJxZZKteJm25LbYeThzSZbogvJPsQErK6NoaS9Ba8Gh4e3yzs
xgLHCxwMYFw/6Ya923fKrPhc8RNR/NWfEPNlw+M0Yttoq4fnUS73qU0aAr1XjoqbtHA9dX8ZtiJx
QWpnt2kFVY0Qj0YerbErjBv5hYqjTtkAxSlnOwOnxk/SGvzV0mLkEYDj5gxu3m/qDxuQ8+pq4tp1
o7VDDXWqMbLMhyRjC9H2E08PTQ40gJaJd+d8lGjZeZzEjzG2VezjRk4p4oC+e27UAE2tbx5r5cPf
2Hea2M9gaYP+/MYVykn+nZ3HEFfb0k4ClBF/4Mdd1XNL5QPnw1WN0ni3C+SNo6YN8kAbru9q0B75
utTaOkQq72QvJmsnkySXGvkvGYr2Fip8cf5o7Ur9+rwOU1wHggdJpqUpAL7mXUelMub082dXQMCa
wB4TbAsnsXg0ZFi72RHH9hvLDhvSQRBz51CGjq7LUh5BRoFIGEIwmW9w56WksxK6fc6AeJ0VbllO
GPWubWzH8mKE5qwbPe7nqw+aFPQBDjBe6dWX6XUyh7lXTwkpvtKk15IAN7iEyOMYoSqUrad5OUii
G/QvD9Pmavus1A2vxemWIjjxgH6XMrnk3ACBWXCcJLzMGmOesb1/2stp31eM6rUaTFMh+5zXqCp7
shb/PDEl/OkMC5eSQtnFsDhgTOxoRXaroaCd9RlySIQzpv2WLOF2AI8FcSu2Cck24VNMlpgo3R7S
bGYhdkU+ebgby7FVaXWN2IjqnwMTC7CTXiBTmhTYFP1mamABtbDl2Ysj8SwL28dbriz17vh2Nfa6
jPJRtOP+5vp+Ezc/LlUCRhAi8IH67oWol0oaG6zTfRMTllCrTHOrYmaX+sE7WF/bnBm0JpXhEwlM
k9BpoMXCkr4spjc8sg2p5FKcpGEYR0vAp/MjkkkFVqnIxReA0WmqTZWXvIEn4mMy/dOUHfYbhkv7
rfRfKX2lO3WdhatYzwAoOLmxFj1BHv84wG0gDq8ybPDR9sVrn1LgBk/T2RoWqDa+WuFRD2shG+z5
2dXIaCdRV+rwE3aSe3QUignpnpBIQKCWS8wqKvNDnWrvD9iROF5+kNDIut6iNaxceHje4pcsIpCX
xnZoC3AHbYL1I6Zeuz/Nu4P2OEpVcmdrc5OPR9D7yOXMCHTasxpVhg5UU9wFlkT5ecfbrLdpjeNy
tFDzusoTshqEsve3jBi4rzRFTunKOrQuLKicfCF2WDQZpPNahRc/UTyhwPGA8Z/K3ntIJZAH0rpL
9XPOQUjKPZ54LO3y0mxT3pwWxggMScuf9HxyORas1ibAc70i6OGqPltGAPWYBHOqS2phgYQjAFLb
23Rae0KUt+1OHzrVdL0fhUgE6xjAzNsxQO5l9tXI5C5oKjbUkNWexbzpD9tLw5UgALzdHAER+MPn
f7PHTmoRmGQ3JE04taS0zzEPz9bn3RP7Yu+221ldsc/b0NYIK4/H+R67AU4w8yDfPc12HYSLWOLS
rok4Qk8zG+NjA9dCJJOAgIJYBMrnWpqRoP1q35bGUZc0Gm3itCKimtof9EcTaisb6oU9VyNQjdUb
wGbDhY15A6nE5Yx2hwJLtxA2eOEWOmwfL6vnXWsGKyEMIxacFFKKQhoSf8NmC4/0n1zXUL8zUp65
qbPn6xybSEubj/6vAeWEXFtpQlOY4Bj2+YO3HtOy1ERHYSsrQuiid8TxyQEWu4Bj/3xl8xAQp1kI
DQ7Qmosq3FVpOChXlB1x20mLxhMjWTUOC7Le88OXY74NEc9xQOOBPb4gdsS5ce/AXnS79xnMF6No
oNrknPhk64M7asAGrBLc71btsCqX0Jo28pGwtRbHomueT25w67vYI9FjwdpcvzEN4QvIBxLePV19
mxoxfgyoSFlPDhsLUlDq40d61BJKt+A/ZcUWT+MGS5Mqruc8exueE1ZEZxsMG2NXKCyKluVXILfb
O024UO79yTi/fs+b0Y9PE6+6Z74W1DKVOLRMprkmAldkS4bruizKU9FJj14Yvgs7ToYCZTSS5eUC
bV/ULiaeCzxxlsaJ4gWW+olbEP1UXQIQlR+CBZUaoR1SKWUvW+yhSqBXjSlhliQsWzWR7ZDEYpTt
W4L9W9bA4uQ4q1dqs4PQANmbY2Sm0Te3oNVCm6gwSblWN1kDU+fuA4eFFc4kH6dzlHKhg/OWHxjn
K1rWEEVkGRpsYjOwwu2yz/mx2vb3R5PkoL6f8FZlewbj33hrNddpXlQ3aAEYi/sJaaGb9BmB02XM
Nk8cl8xyr33KOdqtiGZd76XNpdTy+bXcdyl0p/SK6gRI+x78P3BBSaXgIYbVwYPGC9axTAMp231E
63UriOT/suDHkmjtajrPxKKwjcm8Zr24jrnic9VZc59Sy1OTMrIiRGfFceW7PQ76pH8CG7pKmDBY
7FG9vORjzwzmIHVK4DLSPMo49LTJT80FXhil+a3Nghc9A1ocAJ2EA/Q/jOLGTi8J6R6tQ68nkVzN
69k0GDXWp/33OnlXvTz1xNahaKlMec7/huwdvKoRWZvFRTBvhltCl8loAPtWCeMlqAc2sRiWL1xP
0dlhtbF/oHDGxWq1RQCywiYc3l6ndNhmhlwuwk4utBnGBRHRxqdxWhK2G3EWVW2JnrJAGCJ1JeYb
c1YwJB1fe2kLFnHJmWFroQen4S/KP5RPePYC6CHMjRvLmuFd8puCB/D7W+N8eqW8/r6vdTtFLR5P
bU9y0FbgbuYmwVyCqA42MI/kdJfxZi8wenUgdwfR5SPRKyJ65Hpe6gQFBvtybbvNLreTxLqppgh6
+afrEeBKpBQpeYRUp1Tfg1JCZtQBTAaYW4od9vgdS3Yh2dLDBpxV+01BywD87T35uwZ0qKyiY4PN
hFArdRi5w7r38ssqyHawKITcLXU9/nBZq7uakkWC0Ll4WJQkavvE2+rn6mAkZd0y7u2AikDFLuQ5
B2D9xaH8d1/+9svq6JuPNZB/Mx0PHCcJnUm0klBlCcTQ7t4B32C8EzkSKzT4IbxB8/KzYJJnyEZu
Efp0LEGleBLXVwlN9pEu9Hi5Jhbjh5cUQyxrIlnDZKvQ5aVAsN/x5wmXSMOX88fjPhwk6KhbqK4K
0apyKW1TLILo5KlApzwsxKrpDQE9bW5yCyyhoM06xft2Xm1M/lXKdyD57JKiPzuWlAQBgtTvEH8Y
6yIsa7ntdrVNuGLmWVulIcuWUHIK3xPZsz6J6LJ13LVLNV7CCLGJ5gdDhXZufJ5nQpKIKZ/luwdD
NgGqrEefkGxCLwFMTBxjcSIzJIvkI4ckEo+g0FNxwqj6g2X+jm1z8nuKvBWwOcfBsDyG1JcSiKhj
KgOtOlopNP6pP0EFTCWkIVKwJcO/qEwAfQuVSN/XXq+4bz16yXKj9yX8TmN8B/gc4ORjbonzabT4
y4WlPWgQnJqtRFh1Giys9yoNVIctYiaKJg4CpHSeowGy0UUMDv7ItTDj/cJQtOUwL4g6HhYgmIY4
qWVXY8qQeNSm8nOLLwzIit1xMpodkG9OtlbesfLKsrpgDnzoP9AChBr1JAFrelIsIcAop8bo71t/
mxDyBlaJ+d3WtRlUR+jo0A9VLSnMYzenAKSJuCJ6SlpAFEtA1d6w224kc1xpTuFxnBT6zTJO0nmy
kl81dFqjQiYj09ZOJoIA58akcDQTKT2dR2FOgGVvYwWI4qcoXaDNBebysnfopzlD+RKyShgNP2TZ
QUiN5hdHKQV5z2NfLYk/fJzEmD787GPsNhyFgggD+eyxJbP/BXsqF3KQ5/wkTmKgWN97Y1GlRTts
Y6qPpWs7xH8+vM9i+uGm+DjtswgD8YY8McZjXOcN+fBtiIXAYBm8DHaghuC9Jrg1P7zQZGm09C9v
tIk4ufWWjtFnZEVt7YXiquWnGiHDlZg6SEUkImYxe89xeDL920V2eSOcPMvUydzb4D3VqGBb2paY
J8HhjBOphvKs9lR/sBd20pN0IZqPxq8EHAvm47zZFL4P9noewReMBDwwI/tlnTSNc3ewaxn4b7w3
/WcR+0yFfXD9dSHoLOXOwlONuthfNSirZaR0iEIABUzWfPSlctMNdVUijCEYjBdpt4ZDc44csl3s
8aIR7NhaGhSQ+qkHDfdIdYRnm0RffFPGOPwfBal0/eNm1gaoxBZ922L4xICnI4FJT4x7q6LMDqFw
Ui+wtNwr8WpjJ4k4ookZxG0XQemMXnB/h8Ba9oidpl3zcyrlDYbwFIKPmIO5mTkBY60LmppfSs9y
Qin90cJ4fFj9owVPjo5CL+xC4YWRqfwuXfqkfR0Mx/9xBq/JVxIIDzgi56jHBbT2cVdsqxtVWY/q
PNPLbclSnpJJnuXUgZNa4LXOjHT4ohfn09cekkKfG1o/jCETbYePsyTJExU5CJ/izM+iX+jWjcfj
aWUNX7t1El5U2mv3puLi/eq0+MGpFQIVUffrMd8gHnV4EtNW54AuBJ2va/k9O+TlVF3XDC6+O7gq
ki3bS4wn8Ei0IG4ZtKiL8SK4iKUe1cHHPzmuy664KdPKnbftl9AlnQec0F+S9BGARhAOmwfErcM+
MObRtTY5+rCdyeMDAEjoMA2JRl0yzzKcv/rJNQrTm1c7ebhMLVEMtnMQoyjrylDsachN0uX2mPq1
P2MhdeHDTuvrrkhaM6HTuf4vnrvXQzH5YclVy07bS05eO8kP04/+WWAlTLT1+IUCzEaxByiKNtcm
mUsQQW9mUsCCTEv5Z5K7GuJH4+LKI6EJ/Hxp4M26der12eQ9KFBXVFX66g9tjNZU69BXe2jVTKgd
YWddq5+HGV3YifVIKRTQqhrt7AScjww8ga4EQVJcOqYJ62gfjHiBLlUQbEp1D9z5hgbkb01gAUoX
/ADTT0CVyDfHpHu5U0Sh2SGWuGMrJ6zE8/UN0RBXXe5LB4uZ/3sQSEQp1slVIAY7CuLFV72GnrLN
unGRXkJ6BzGctN3HGiYJW4Tw/7Y0q+PEXNqLELkfuy3vMyeiT1d4n1k+TGuhJvvDLWhLySNABRE7
2m8l++mEqMbgSadxu3+RN0G0i4yPZBdKGZKc9QKX1+t/ttxvdJel4OQggyxmUCAjpQ5caSd+3vXn
9JT1QVbPZLLHw8N5hM9NwPk6s6MbJUjpky5QxyvH2m7EDMLJHSW0qSKiDrP5ZDKs8GARUoAH2aSs
9yz0xHpFZqGWnzD1VKBGrltQ3GlGjn+SSreDZQ5qIREaMBtP1X/Eh9TDtilStG0ALpDQORA0X8Ja
52Gq0cgZWysjDxJaGVtFLMEXHI6YeJhzFmOVxHI7IXpyYpwmawRGeoxhCXwFYDilnfXMZRlhzwxS
qhDWoW/hZMKaxm1ucY/9NN0I4y1dz3irfqN6TpUba3aiRHzxm89gnPYbD462zeU6WBa2+UIIlHux
Em1QSM7gyWvr67unSjkV1EJeLXow0WY/9pZtkVnagQx596uFMPiS16Zp6TariLNr3UNmgUOwzIqy
gFxUOvlRCH/p9lUwDDSBJpP7JjGFpjgXyYSbsQAT8KEQaI80VRv65cGICvy6SKwXbcGbbiOiB9mU
cAaYLJjGVgFm4Pk6ehqjd7hvTxtYEjMGwt5cKRrdd3AWTV9YMuLbHORQn24ksZOPVtNlHWy6Dr4d
GbcmAUmPX0XQvmVjU3Q4Iblj7C29KlwBE1FgdmNCS1NEcBApA255WjPsmMbgs2n9JzhmumcJGhQS
Srjsy4qJESki9GIElAR+5MEj73r4SI/AEwPxaLGbMcE6YS11wXQoByQNL7paSFpiuS2nIxDhRX2v
0QTFlJwyWILBJCklPY1hIIind9n5YuQNJ6j86Lftx1Y4f8g1NBogSgN/9P+kaurxX/nhjC4ZPXE/
yPEiiLaoBi5iIQ++PxQMp56XSs/3KXVggjlZ2fYUVhIYVO33NGsNgP9WXfKOPqyyzhi5/rJEaRJo
U2MEU6nndFwFU1sdLYfAfA1urp0wGVN5BB54U4ybRiNl3H348+T7qCNb7IbUl5BMjJP67U8iDKcA
pv24rQIwEk7jWDe6HIbfmEsQ+kerWUeZJ0sR5jBJHmJYrcPTJzdqq4+rtmATvjtx+5W8dd6W+t82
2vcc1W/ljJRBBF1p/HG/exKuQVsi4yhD7sgq/wVtCxnehlt1HrTES2eQgNa6HI9RFfMsaXl/2mr5
lT2Gg9NObydrKMipczFtDyLF4AmJ+ij3/r4KDyGhdQSwGoUf4scBWdweTi/QHioGvT9FtYCGEB73
0Bx7W7aomsUsotCgH2diVpDlwqHaZ5Ffg77pr52tT/F0XYnEpSCaJOv0yW2Rq0LvToiDTcvO/R6h
gfzC40QUWgmDWyG2dqvm91NlSPzBnQ5pb9vK0NhMT0ybAVJW2yGPXp1vO1a0umAe4Msg+9JjQSRw
ylb1EpPGYokrYJYEUDo/OqZ8T8RakOI6xH5ryW/R79RIHGwURQ3myqgvfYWQVwnLnlACve/rDvT9
bpFc7E9g2a7Uefi6zf5W6rErFo/zufVhuodOPcJ9XOmN6qkHpP726MYWHLRohkyl7Ddc6W0MiKP+
YPSGm9AEN1iIO1WcKGtg9t7TEJRf5eNIlnGkjPy+4i0AzEKyPhebJXkucEKStWdTPcHv0g5pRnv5
NEejxcdv1RekaDUFH9hiODcYMT7HNerar6MxEwaWHWCbqVzZwI7qtmuk2OlhBjJP9UhSjRBPtMIU
VDvuVFB1VyCH0TDtvE7miixTesZeLQoC8NCGdwhedGeNnwGNELdpOCBO18OXKnyrS/g6hiDQ3RZ2
R5sokp9WBv5sa+EMt/pH6xPSm54+72iIaoD76c2a4V4HTB4kwE94M4Yshj2SqImToB2tJbkey+Y3
sNIbbPbHRiZ3/ob7Z/EqboV3wbEUJyeS4scJLYruOU6rwUuNbyHKFn/WIxFnA0tiMhFN5CZw3zFD
VFRdKaRPWw+lPRFVYkucwO50Q4azfdBRRCSDlit0b9w1s4HrJHhXRyxTSsWhAA3mdUqrjdG0CKhJ
zola+riMwbFrS86DwSWRLnEs88q1JfCgW2vg8K11M044YVLvVM8n+iUi63nrIPoq+bjzgcs45KN3
CmhU/4HMjoPMUuRzwElE1VMB9I9iNKAJoONjRfS8/SIZNU8C7+NLOVe2uQ5Z3ved8CejXBwEZagW
80pNHcxdwn+Iyi7k+X3o6VUcEiLGs12ANeoUkThb2i+hfQGTVp4p90Ov9zovJfD8iar9GK7ZYXhx
VbnSB8ewrkIbrDZn18/tHFC/L+2iNXLEBk8Y1CYcJctFEmkeHUZPY2BF54JFc0OIywtW3xB450yX
DhyKkGAtwdrCuI/2c9anwpRzFSzMJoJdvB2V0UdtXzRWWcZc+xKKdKSfcc4JFrZqgB6tHgwdaJuO
jGCC98O1sZjfAABextqKiDxDL1qQ2CXB9LrDZnAKoqDW2Y8boCa7po7Kbmp3IgKFUAKamPgf+tII
7iY4SEYSaoFrCbu/cx700jP30jMYRy8nYsANIW/N4nDv72CbcduBjRirAjVd5pxwdrlZknJYVbT4
nTXQ8PSshG7MgHXgdp+Ge3ERHlSQWh004dSf9CcnQNIsBOsGP6swLgA3vzomdEHuyQVJrQRNe2Ap
w4eH4o3eMO7ZOFK1Irrb3gHy+vUin3S72tAByR4pzyTPjuFez9ufI6V+Xvy676yEZWBWPTrzrzkG
K6Ijdj20SqRRchuB4Acra97z3nW8b+lmsbOilwLwwB8/rHl693g54FiAhR3BYGdIRXBSZ2gKaYWE
IKE6kZJcGFVrYiuuLs+4GQhzBrU9p1lcVsYSNoJUNffKcS+w0b7mlmHaCNZ46PdQDT4wtr7EObcu
Qo1xY2q4q0VJCVM1XuUKh5fq4tVCE4Fhaim/WLkZ48EqIx+Q+fWU9SFGhQolfzt1iM+z6UxUj5S4
B75O+oRi8NNvUVnZw22I2BKSbuExsKp+g5dc3oHjUj1gAo8tbk3X8mijd/H21mnHall7/M3li0rc
ZNVZhErGDv66Knfrsq5r9NFvtrmCXpw3HJbf1QHJ5Q4ktg+SKX54fXXjARlwLZvImiNGMbE/2Tf9
SXV5pR7m5S16fu0SoiXjtC0dTGWCMyOLIlqTpJhruuyzh+cuU5436kWYrz5jD1Y6uQzaK1k0HIE6
Ow3xKbEPjtxIJESLg6UwReftcGkLQwGKPQUrrtMmdh3nQstV759QfpupTvYZwfp3lp+a/Gif0Iqq
oB4V5VvOtLvsOuFMjUbXse80XZ3bA1kvWNYTeM7z4PKJlXnOXnGjsBOuEhBIyMQgZs26nKJcnYAD
fCVmWVddU5YobOixbRL/HrDI6eVXhT3HbmsbaB0JQas0PQfZYuVLg+KOJmd+RQkazZs0LRn3SxbA
Sj9NSvfMWTaKrp1PoHBc5CcZhfISqosJQvLT5m2ZnJ34BhKoLviSU7gkJmQC/+/ZtwBnwTCK3zh3
FnpRUpBjo19MvTDfviGKqCK22fY73pjbc/jPhp10dTXxhqU2Hrp39rhwZb4wPxag9htjsRNOqLIL
s/WLzCMh1UBIRSekh22i7VkgEcSGUdUMHAsPabX1CTFmmH1zbUoz+6Ku58UuhFerWhV/YVYg8rmy
MG7298SjqgvLqmV3WtrRYqhsr8nNdWB9sESGC4EjznJoSIwwKQfREQG/pbFnwcmPgSdDVTcjuFsm
iUR1QjuSbdJxNuTJilKG0JydcqVWvtBsGdnoGAUfSjPU8b+MuvX4ze18LZNkM5aya/OKugDjQOXk
bgroLRZ/8dPDjKT3ZSg4kwm3ZUyIvBcdUsykbT1pw8Lzdz5a9tuiNd/qo2viHbr3+nOFrXQC2BwW
kYDRcSw+jnTcrnuXezcrxdkOKJUE861VkED//lGsGIhu0vxSPk17mQOyDZBHqgjQmZ/Gu6N1LIo7
KKyRPeYMq0LMphez9z/dQk7cazZoBUdRV797/GHJ7JCP8BrA+Ibza6/SzJTYUAR10G0PsSFgCHUs
jWiPuYTB2hQERmJX2YwGn92f7/DfPpPxlImhLndMJoRM+JoDp6DTx5G8HF5K/h5y6orpEwUhMM9F
AD2UlKw+9VNM94nUmW6IsXkRVrV/tE15BKihVBYeIFRTDpkmbqjEOkezrAnsGjplzgyS6G3vbLhF
V4+t4Awtvc85DyArGiV2Im4kRd1gSbL8kWkSDSzBd94qaWNZr++JWx7U0wbrOoFCANMY62PinFAa
fFSgb19Txng4Z8BlWpu9RIxvyWaUxh5UgkXTI743j62RMmPJJgZivWjI9+Ah9MadPDkYJPqdHZQ8
bLmnPmpcoz7T6CV7Ov6Kbg8Kr4FFYAzx1xZ2/2N8y32vP1vqqQBr2YC8+obCvo8FfQTwQg82cSWt
jZAIoBODFFisJcPv4QFiLgBKLO2aLQAO+PLFKbLPVs3gfylc85S8SlJSul75BnXvI+BtJ/MpCDoQ
lZ/0+U5XErl4fIesK/dGvlDxxgdRKX3xHU5IowuntMneRapPys+qLQKnL/LKF0mF8rRcw5Xf/iVe
jcSDEgxBh1PvQpNKF2/rBLw4H7YMl//NE1KxVCRZUyhTX7EbI86Ua4UV1cHqzP+e+c/mdkShRnhy
CF6tbQyYq7r2uolguULCHfirQq56Nwq/IGqXDRWdPYu3k/nDU+Pe6mQOTaNTw9a8PCFDIQ+wL381
zIxOKviVKJLuc8YSe6vl5grw9qaw573wl2bKTJ+2/uQlYLIy1N2BMzgI/3cg6GjZLXIIWE3u0HAI
5z6dDKwp3LO+6tqJWbgC+fh4FEnqI8cePR7Wqz+P/NiUb4y5d/Z/yn5uNTS2/g9WpKKn6aSVmOM0
V7tkrbJXRWYsubz96o4dON8rEgS3UoiFUpqt0o5ItaBTzJYLytzdLl37iZsLroy7C4BfaEvDWwN7
9ya/4Dlhhu1DmvpfFkTbiHiAVpyar7m7NWIbIupsVaqEzppSEmYEt9pBjF3Mwq+csv55DeQGXYqE
GUHTsJ5vKH8YyM6Ol3Jn9kNFuaS3cc2BVQbyZwZrXRLYjvqjkiEhHUOc1D08KGwLLSnCFPLqtQZe
6Po3bJ8mdgYd0FXltWP7v3/p6L0IJKu2Xz4Oevr5cPPhxf6st2ypRyWxL1CPcVl5lhUBJAOTOzEf
Q4VnESn7ssm++PzaD22GhHQgtVkWPGDtq4YCRdSUlqQambJX3VWa/foa76UhvBYWPIxGPIzcKq1C
HiJYDnAF2kAwfOpZ2sM5KI3NyZHuSSl+6Vd9SjTS9uIaqoEth1hGkCFLKw8OcCNeOu3nIg/Tp7WY
wLpUoSUV84eVtgE8a3ccuQgKLOBlXsx7JDhzik6uZoZn0LcTrcln1ZPNqosO2yJFmekWUthWWASc
jEJtiUBhipu3coVFoGKidOYFMHsM/ddahf6IHWlutphNJTK402ZOVa2XseDvQPBTezJzCd6G2/fl
avV6fdEWKpN4KONjWHWDfvsA4R64V/J4ij8bCO4cBgmmvbVP9A9A4cSkDb1y7k21+AvRCaqO/lLM
tFQqHx9EA4iVB5kvd7pFOG8M17KAu0VjWUp+FBtLmpZcwTxiAp7Pnrc3XSKMhENneyIrXCg7/MsA
0AANmrqH17owYZLj6StKwUbk0hDzBAiSD3htxs/Elt0aBVQhOLr7DMSZBI5pHcBY7SI/mxOMmUP2
rAKRhvWXNsWZu/RzENy2/fHfoTzD+ZS1k6uH7ubeOU3zoT6NEAjMtZ955BAlUbcGfOwDCUmbpka/
CRtJS+bqtW2+RAykb4bnemAJq7MsPus8Nu75MJEa7pBkDuyi1TMokcqu2UGOK2jaUwafYRI3S+oR
t1JRzjr8GpPGtGBikeQ0cRD0Sw0Vvt1Y0XpD04tMeCygrF+3fxx5poAzXaVepZqHOx+o/lrtESC7
TAEUkN6kyodnJFT2sf30D0Ry3HexdJ4ZUpy1Hq5mNtNTtUBpVkMYfMNYZVDkp3eP1hDw9S3KQFQi
upBiUJwgNVV/LpytyslDtDwRuj8AnOEDLZYlSxdzJ1t0Pw1keXqgjgWQ9gwhRsSBAcBzfhmWQN1P
YeqSXflAmxSKC1DQxi+NH4lI/zSkeZJsXJovtGka8gQ9Nn5cXi2ChXjsZbpkjfDfm0hzaIEpuWRA
EryL1hqiMmCOOjvGkkhnUkN8CLHKhff354l5bKksMExKKvwQEHe6YYZVrhZmR0CdQKi4eoTSiHB8
C5syIAykT7Gr0KdVT0436JksP3L4RkRRS14NoMXbWV9rLb1ViFH5IT+jU+feNy6JuwRUkYtR35Sx
Zrvhh3GwJ+IJTXZN6A1kZrwM8tU3T2NetxJAJGaj/1dltRvDXqZc4esn3tWZwIlR07KnWzNFPhic
usKMIYHOm7ybiWIOF3F3QdL9BnlVBeZxEkNZxFxZ689AGJl+2aW4DGj5iVK0MeHRhl2bGj2guBPx
DrEPiIgAwhNBD+jm43My4BzP/OybKVEyrBS5X2NtZsWOJ6FX9LslHpYXECADT/7uGQDlhCVgft4F
X/f+0KOJB+dYU84VMMdEHsx8XqrhLiuslk6roBTvVkTg/H7fBuDyH17jSwEMI570nU5uhEF/B45D
iJY9cNuN24y3KrEvg2rBZXG2y1dXd6JLKFhZQHLSSfx9E9SzmzhucC0T2zMk49BC3mQpBSavhyzr
YyU7PExhRcoZLcxt4PNY6xXTlSKq0JBtqU5JBcVJ22Y2kfED4dHx+iGK3qdjJLlxXrqv7gZZPhKc
Bsdk4YG8WcqkFhoXtptcyvSgqmMt+88G3GawVhCmehJy2j5JFkOw5BvJ53ueWCa/JIkTo0FGQ1Vk
G4gysBYDW0Yxazu8AsL25fFsZVkGMA3w1yLTRhgaHlxL3uW9nw6sqVB5F1g5ceCqW12f1JJ1kNdO
+k+9XeWuCnssWAaB9GUVE6Zo5SuDewqQ6kibea0wA/ONGg2AkPDNrDworQ2BZ4+oFWp1To80/gXf
Tiq8+R6HZTDSXAxg2p4NbaWhjc6VzEsYnF0qHrgfPSfNWw6YZxa9bweK59qF2593qUTMAcwdNF1+
SQZenEjGizUEYD+YxXneoCbXfZzDBlGTvA+7KLUZ3TEgCn/h75NPDQ1J5J4GyTmt1C1+geMPn2Yk
1/IqgxlcztrLsoQCmseILQw7/rSgzOyNPEPUq1ClCbLsQOqn461ckIPu0umMgOa9O1xWPmJ/hAdh
MaPAynF+uh6s0r157WlNZcivyGsYpemw7AI75wFsFPheoeN0cO2DSTbP2JZmgayc/NvMRXzgEbmF
yHguR1bMrlRLuxLX39HM9cV2UVh8NJHyo9PGHwbIEEiP1USLWEKSSWIA08JfV1zrFGxRbXfC3dLz
gNuJJ/lV+7yuV/tXb9W6Y/Xu151ailvaqEMBmB3yCQE08nI0XcbTU8lNszoljkBqd5GJR5q2Yp+S
1kTdOiAjDEotblgegOYUsI+fzui9azuQd905Xc5S2KghiLq5vkt19abDwfeMKtCKGcWUxbtXANs+
lW4s25ByT5BewB1BhZEP8DnImP7SG323KSscmX5bYctNqDIhVpU6FrPvfDP4+3DaTp/e3FhqscFC
4AGqAfoDkge0BMYLZLb0KBMVLVlywRdspMvssMMQ6AnnyjzoyPZE7rLVX/6E7q2GljCGCE6Go8wZ
u97efosfJLCziPL7AYFqa1SPRwVi58lnpq6a44L2AsShyE2MXlg5CBfGGx6sfQUmbyhbZ1NrV6QR
/P4OcgDCMFBooePncguImb8yyRc1PkrSEiccHVxK7fkPXmvcYjvVfxBo5fByg53W7/GbKdpxUH/e
BSCi85KC82WSK7AX0kvnOtHmk8uULi+Ox7PVELC2sy4mkrNIi7G5yjVGQvySQumkFH4qm8fVVPlI
Yzip/bytflH5d6h6fcvDIoUhsU/trFjN4VzyjmxREnNcO4tqg3bUE6KriMI6Hi0RjEND/W4czEIM
dll4VrzzF43NE+uuWEqAxytQEQlMgisupeVMGK5PBWpnPGWbJcs16TvAdZs/VaKsbZCbJLCzS3s6
6t70FwAI1v2okrR0Nb67Sb/VukS9DvScQxGjjgHh8seTaqsUaqkxIB3aZaadLN/V5fWkPRFhOPOL
nsztyURVdHXRrbvJGNtjWLuFGrykoTxnpXj9SAWNM1hfsAGUDMH2AsqO9TaVd4207VKh3VlPB1om
VCrjfd9rdUh+AIgylwXuJPh1XLPXKg5g3X0eppKng2Aw3iUAN1BI2pC7MipqQ/MU7NGAw0hJcZ4A
gqnzV98SsN/GzNoXSXJfhhcx/+8hUCaTAPKdq7I7KBq4l36/2//pcCg8uOBhltwTzkLzTj3tma5e
r4UGtLLNx6Fp1PffABn8zLWYiGHKbFOODbnNR4ujZnZat32Ud/nXFJzG0OhbaRRqUa4Z30yJt2aP
2tKMvt9t7OH68eRjh9MfJxLPUNqoHhep5LSLz/OQb+oVAEK8By+5qU7ojjQufcI1PQU6fp8DpFph
ywJr7iZhOttJhdY3kNrSKk45tFo54hM/aLbQyXplToYOPiblN1PnvpQbE0sApXNiThTEw0g9zaIb
G2RoWUfMrvs8uBRcl+HOqhtoF/R8r7/VE416Ior++lselalyCIiOHdmIvl9krzFU+uz/1ZHfQhC9
4mY97kiQs8NbB5vvdDcNJdJ2qC7sGfB1munlmaFKK22dN8j8Fwt9vW30EoQuTw1XxKD0aj6Uen/P
HJ5XIwQm0+zXfGObrc3iGLR3WDnI37MMuT+ogz+4v0OhR3AHMemMVMjIyVSSsUgWO1k0XF5QFwhO
hZNsnm6y4U5dQOWwDYLVQmGKgJQPXhycq0htUgOu0nwQJJZ7h2YvvZlFvphleJ1Wnf6OMghyGpTp
11b9hPq8Uqi88eZYg74oiYTakI/IW+kSUGgcyN1CBzxh+0F2UceBjMBmJaHlm3MngWwkjU8tfZpx
DRdQHsBvFN7Q1KVe4XFdaV4lcisYqXQ+Eg2IsLjol6/5/bSWcg7quOEskOYzB2G6qkTCVlGd89hb
4c2FWZ1M11hHumuqmK8ENkStMepD6x0CQbsfTXjQ/JbYa4wj29M5IbWVh1S9VZuYRJaBp24PFbar
Erho85JYV0TGcn4irFLYW5sJCbwRXFeKp3cdzULLD6SuCARhx173guLMUGVIgLk8rk9MCMOfFgTy
0HIoYztO23Q0xOSIAtkZsua3xtNyo1rj+/Kzlz8/u9QYmKydFp9JUY6jUtOdntsfZ5NAAP/r+xOg
6nYqKyUoi4BfSQwRoji9X6SyfGmYR8mL7fAg/zZ+PRMOpeA+JnPPgzbSrw/aVND8CH+btUfyKQ9s
s41o+h0nB8uD9BODle/pSSpQPJ0/98uHD8++lrqxHxmnuYmRKOeFSko/zDiFW6XJiv8ADDs6VI24
uAlnyA924ErhGNAcm6V0bGrGoDPrtwf9Ly2mPbJKwwLsrmTb5JTKgaBFsJ9/LVbZHLXGN2JNHmgx
dhbwrEi5VpkSPOnwhdAuRqtyT5zpkH3cwFev1yR5cd0xnqvsYNeaxV3znyuhPggZIxl8BUgJuYuW
vthbJ8iaND7zV4RstNx/2jHIbxKI7yURGpeE7Gd0eAcwu0Nf+nroqHqumB0aVweG3r4mUdf5DQ0P
f5ERP8gR7pCDc9nIAVtoQx1pIrBwxJe7+Y2eOQs/anueI0NxICf9KjXjad6CWw6XvpIcxaZfM3kd
HZ8e7vF018jH/lJEe2ZZsks8Xf3NyrCWXA4pUJ04giHaG06lbu47FWqvh17VfFGREJtTTMB85N/Y
2lKqz3zN5PHFiEijNINyWzVVjQph6NzM10JjQCI7c/5zxG3hQHc2HI06sxv/05fPjLF26f3Jvr30
BZ69DieMef8NPr7pbzPXkTzwasWJ86PxsmlmFDmsM6eVGLspefVbXAkhll0kkylZkXvk1c1l0Osr
JOpbPzMN6loFO7pR8fo7wmzzFExRcoMxz0Y6+wGKnnIU+9nB2YZqEFmqxMIuetnSChdIi3hxL1uN
o0nypUeBekFEdl6dRGQUs8XbtsuNE3J6X4gLKOYj8MRuTButegN6i2k9hd+LpU9BctUxnVyXWFAD
JcudrfyofeC9sJi7tv+Yc06X3q1lcr65w3mfiQ7px31R7yvOj/6uaEilkV5JKfOV42qjB0Uze2OS
BOm1JJD+cEMnufKog8ipWnaN9d8vxqlFOhOJQM0Wfq0NUec3vU7coSgfJkyxhGNtmhL1Mm0EQKhs
eT0wiqqQWVUkHopDdOaA5HmVa/pBMRofE45ERKELLgbNTU70xvr+i/ImFrjY48VN2EFlKggTQEHo
0TgRC61mFtQHJegNOCqzbRE1/ObnowmT2aj3UgROrWqBTgURrfDJ4VQGw/IQkTk/j445R6Syvsc3
UjaeFHqWao0yAJYa21RPrw3j10kWHh0MTTKLp8NqqE/TDfH/+RYsJ65KkmKW2uyX6Ypnz9gR/R3A
Pqb2fq3mq1+tI9YcvUJ1u5BzBvGgVUCie4WGJmKv5DLmKJt23QMVprm2bJOe5Up5vc2FvEKGv/uU
T5IiwLh9Yh0nFcXFQLQZ4NNWy2Fb8jvc91FQZPvtkErC8bPhhcgkjylDXPclYfuGHHoxBtOCGp3q
uHPt9AF5stBOYSK82LZmbe5QqddNoI/lKk90NFnDaixz0aPsBkp1fV15I+0ppvt5hyb9KNXhHeBe
1+C/909EP+a3wyEayLjKYGK/colPVQAHNf23D+zfZDd5dg1UWO5fhd7GotZWuYv2bKc0axuiu7E2
tWat2IwISxXFKg/qrIgAv8Dkmoh1cJ1JcKOUX6silgbCoz3pY4BLBznrGbMpSJjtGC1LpRGGAnSZ
oEbGu3X34rZQO1VHRudZGkIciUFFCIAor3p48wOKoM5tZph+FTplno9TF3CeGQufWM04Gc9a+ocP
/yNf9J60xc533QlfgTIh799KH8SEL/PraFSiDlOP8aSCVxEcV+FluBHA4yZmFb7z9Hj9s8p84nLF
JfcD8MVg/ZhR9T8BtJ5a3SQvLMsLNy4MA/TfNJ4a3Qrn0Di8rzGgyjop2uOdLlOKNhXOYTph3ZWH
+nJ4QDQhyZd7Wx0SngCyaRTxIwcstypvCJQeWPjzHh8GNT+xHShDJFTGwYAsGrFTrEM9hPrRtwpy
loE6k7iHOaxE6Y3hLuaqh/jA6ycyrJYZjbzWxYRXIR9CeYqhA+Ipx5SJhr7KU7TLAFSBjmYYJ8Vl
YTvuHJp8udtTOvP3yiw0KAqV8YiOOp5/rQOknWmP0TnaY3YES586sZqMWd8DHM3+Xx7eqCu9Smcs
wXnIdzLg58j3MFzoi8B8fme6pjFSWZIt3an7FoMM4VJJxFudQadmhp6pOu82zxYE5xoqOxWBXkC3
2mrSqwCIZOnpFxyjJzLYgDvNuw+ZZ/4F8DrhgWdbmcdLgM/UxvOVnlrdtZ4YKwEcoYFR/luciRej
F1Q+56OWkVI9qo1AEsdDl8CCtGKhbxQFX2b3NfSnuGjphzpdTdt+VXQupbth+eXMWeXILg8gXU7Y
H45sB9GOzcw4C2KxeFDUU/IYaf4nNK9FP4cQuxBZkgva/m3C3HpTWVgxvc98tvmubNgIvOXehR+W
JCDZxrpq7eoGbp8xi/hZ4BYWOyIFrYACxALQAAg2AEPtqs4MDq0EXVT6oCVNykDKA8/i2eyD2RKI
8f5LpiLCwGCRd04sEmF6qcbZrXLWyfc3EPYmcpnIg4nys5LZXFYzxVzSnVMQyGxAcOM93lUnLvZN
Zo9tecwEokAafnUZ3opqKEPoHuCtCVes8aS0zxqon+pd/6/otw2UK+idvlYHQ5aRu3XcaiFD4PPS
RLFc/FSXLuG5dDpktt1LUCgIEASy/LIUDestasxp/El+tIW0t+DiOnlMi9af/Yy9ixS7jcfUuC3Z
Xqry7ETlO6s7r1JC9WTYozCCpLkEkweTzDWllOVRWzQBlCRs0XxFOS0oFEnRqlSLcc3+8Jlv2r/5
mxA9oPbw0k28P4J4NwLMUvs8UM9JNXo/qmQdeP0sYx5iMLrLqukR217tEVqpPDc4qix4KNppSIO9
giI9KBix+t6E+LFMdYo28YZkd9phlmkutrKl7z7Dsp0KlYVqyueg3Uvcdjgzr8Ms+obQTJyDu4Qc
hhghXqQoJriypGDgvxkQ3+GwFgrtaxIj4a1H0QV8h94Wq9jojRjYMPt1ucPUMqG7YYh7UiIqiFww
g4sawurpSgUOn6iiSjaC2aKNe6KdsxG5GOwRld8pruCPlNRGsWEFmouhhOoJguc1J0HfGkndyiy4
zfaJPbFPev1MH4vuuF3kGJzOWWC3AXJlTKcT8K+j0zN3x0JKu86hH1DdeHSMH0XgK1WJV26IGtEs
+0+zCEaoUAvxfRjxCiQ/B25RTejc/lCQA7D9C1ELMkPkMHVUlF49QonYi3bN0TrmQQt29XPqpwlF
vjk+HJkeRQfvpN2SIuQO6uEroaqnts2JdzwlKv9S4XgigYJwju2d3iWTVsqKdFlK51ZMdElhl4Hu
mICV3glYrKkpDVDrvUGItvgHjTazNdReELm0PMLNU4rx7/sMojqZL/gM8aquiToIQ7ss3BpvWTEs
zPIZ1gjfT3GZpOkHJfJdhORg8eR6F4BWq8pkKvDeru7ZAObkNalJKdTgS2JC75V7sIFfrdY0toA1
wpe8p1g6QHtKtb6WhLnsOnDOaTLg6WfRBX/nV8UTX+e7hhVDGQzAl6d6nhkCM62ieswp1U2rlL92
yLb4X0Jaqhd20XE/PRY01PCJEmlYbXgdBHGKlS+59IKjeRBtHtAjTERxdqPKh8MHxPsm9NqLj0bo
6uFIoJaGVEgPaSN+8NUIeMYvejrgiqqToiFuUqplOLPxq/Sv7xjkbl2fLRX7K2Gw5ChPWudUbwZi
ssV0bgVAWZ83XrdBRwKw+4x62zzUTa8FNrRog7iB7k6++W/zlXXFCjSAcCEoWp0MNRUkPlQxgWjj
1vBk1HGa84sHHiblfSRAUAddwDJLwC1c+4HkWlEoIoLs7fvbEet9lLNcoe7lsNVJNZHw2X3MLrIl
wCmDjNVFaE0oBwAZt86ZhsqrXLf6KLgdjOuwYck0WcDTy6ZU5wYvRacIkGHjQLqi9KmnN9PeKVHq
uiv4MWXwbYuXsqdFkbdL5S/fuDcAY6bkiuRz9GRJzcKKpkFzhgmuzg7Qw3GkpLsowVyEVuTAYCSX
qw8PqxKXq/uM504x+36Hji8SCv6+CkoO/LngU7zrqrlMV7RW5hL12+PY75LDAFEmheRL19gCAya1
4az4JMpyuf1k23Q9BwZaE8itPT4HZjExciIvIPfYjTd+oRWTY5nGmvjIp7UzRE92Qh3LJOsc2lDt
Ct8ZPQovfReRs7hJkD+GEbx9h6oNPzJKI5g9fUUlh20c7HRPqcp4ZXAzzOT6rbdoylmBqznxT+5+
0WMDXZvYTdCC1aTSrqOTMPt/N/0HaQSKtC2+saCDwvdRWousqbdG+GjECgJPDD0UEV5qOlsQiGK5
s/3io26IpTGWn9PWFLBx6sx8KHTTRlt5urTelsOiDGGNlcj+8ty+2yyWhz+HJD8+d0zJQxs9M+FE
unCY8P19LIbs7shE1eGxnpeN8rMZ/rHnynSEaWBp+eTciQmQHfCC2NsyYRiBZBmq4Di9URHQkaOb
fwe1cjcEa4ShcF4Qu3J90i8xKi2AFSl/9QldoXeepIggcTorknQW36KCB7qflZIhxftxrJllMgYK
tIyh6uFjGxAFZjo4gXWff/6jXKwS6Zltgm806q3UcZjGe3tIAX2Ybk+Lw3IgPubcG6bkSI9f/h7H
SJYnB5Dreo4U5s8Bbp1Zif9TJir8WHVMMVNqicereLRv0IZ/QodermA8sjJEwBlZJSpqLcP60M6M
DWGZECfaFE+08+nFLyq1d1zMFfbGh1RVNL52SOJd3tYWr1rbChBcTCrJ6B9YNBwpinYESCIj1UhM
0QubzO4v8n7s5lKJqMO8HaSGxq7PF+YjDgZrD/rJ2tNZIv6XelIdjTB73wSSbGjkbIrsHLX1Wamc
prX2NOUlFGJ23tHUWOPVKLslQxslldq7+xq1m/tX2cVO2bPMFmpSKsNfZfiysof4xyXWDKVU6PJo
SDRhR+HxKLP0aI1Kwr7FnUKqgWkaesoZoufq5OPndzSXVeJ8FPXG49lV5UndAegOfz7UQUYtEYJe
23JuCG56Y3dyZ4vXu48219TT3Kv1VfctWsVHz5x90J9SUe4+nGwH8rp7DtYNXR1ESJFQrhuwG76w
CimOpKOWr0vTOCJtVhzTTGllLazzWfYpKoJa5FPwGn3QpOKcvZWCBzTQpkvlavztJuI217+S/dlc
IY1nW1+nEbYKBYl0YkRZB/MzcyiXcnC7ORc5SNHYqctPCei4aslLK2YK43MhkoBqJ7PCCGMAEwJy
pcDMoHdDb0zUubqYaadNEkTe57tC1oiCLjMw5qCicNt6fYoYkF/6td9ndx84jD01FBCAgSa8k30y
aFr/jrTyuQ6MzAin4Ez2cdltfabrrYolaMt1gyzC32vEfBQVbz0j69xEK8aey7JNgM/oW9q1/LGY
R2z1ZhH/PpoCqLPF3eTRydi8PvLzm7uW6OrwnHRVjKnvtOmCMON9R8Y/WmMstc2+tCfpKPNGvnL/
PMz05lkHwVz7Ke8FqNzKaZPiUfQ1X5nC3YSZBwuoBaoL1FRH1sDpgfMwgkq4HNlPSPXnasyqNpLQ
ntdWDmA0oay6D4Qe1WUjCUu0Wz5IPrORkWlLnXI9pLEwzYYFYfxz1zqjQr2cMW2t8bGcQHg9gVpQ
w19YBEZlhRDPwY1nXKq790MfWSKj1YsLHFA1AH8kIPATfDbx/+d1h8l/0mpjCCTUrjfRKUPZbPqS
m2Ctue1ckyzILpIMr7Lrb5Y/xyT+LrP7QmyE+xW7v0/ud7sqYK7lkUs5iN9l2GfLHXMZzRg9rgz4
a/MQdg8+T4jYeyIiDU+8dryygQnMNUE16qqmJqCN0Xsh2bKcr5NFCA7nBWrX5scX6FUVpOIE07aL
en3/myPbfAwGy8wZxs/x3uGwmW4W6tQAtKJ9xVQj1UYSsTWcCbZY0Jiltfwg1HxYTiR3JOiJicfi
VoLHb/jjEAtLVymKWEv7v63/875m7f1QeyztL43buN9ft/DG7bL2RouxB8FJbNuUNKu/aUmXEN3B
MuBUgQeykZ0wy1IQavwKdBNJumHkGZHNH5vav6Br8X7veLZXueAF9XLrDqn45pALfLx1yK5GeuxG
DZevR0vOZBQxszkZhufzvF3TnRFD4TD+G8Slv5mfWQdtx/ukfeS/+xxGae8U9np3WmnMiz37vlWY
pZZuRzH6ezvUzqDFbOeiL7PTaKhOhuHMQH21EpGf6AJgYFo3Go+9qJNZEeGkfl1yS9uF0ec6tN4o
qzt+pzzJN0xzA/Wx77XbYePKLkdW8Dja7OY4jRQCPI8aP+FXAh+zplqVG7lDo5wtD3sxgx+QHeLP
HiNTdmD+TIrfa5V9wI+TEPNiqQ2VixTzK2jfTSkLVLDNcupVsLtmSlYR89KzhKIM8wu821P8BsAd
DYxCX6zTAqu8Dp6CNXaJ/v7sRKDzyeJCrLrjR7PNb9BOrtgVu+Sy7xOwTYgbnHOBc4yr98qG1iyk
PxKxqAvrDpPVwdDfW9mRrY+O0A7WHds34LQcW8yqXVPKXQHhmiVkv1StqxtV9kx097ZBPRksaEJb
DOmjlXZ83S8Glj+xQ8TGBHgEnw6Db+1iRBPMuNMSxIzTYjY7C9mJ5T818Y0oDZoYJhV9p584L1mx
+zGk5Gv77LESahOVOf4K5DVDLOKrPAhFfsOQLCuauDUcfHlJgQKL+kXtxjtAPlimsIo3kaZQn6BL
NPXQrKLxA2fAn13Z/Mhv9RE9IHsTDMIXCpy30Y9Oe6TU7I72F/AW5XbCMeVBQ5jX4+sUuGRcrKYq
JWTsO/S9rFkHPyJR2tp9TYIxWekCKxxhke2M8+3+oE8V8/lFivdyCMxbIvMQNkHVmGHTB/SrLuGF
Ha2+JqhNbQL+BfTjwtlp1CBMIZtoKcxTqO2o6laDUY1OvAqAyWYQd0o44i+U+QGk9840w3pnTxxe
QgJDOidhqs0IJ+NetbpcBXuYuc4Ie4kKADvOcvSXamYFEtrk9e2CwvtIJZkIsjECXWfZsRHBvl3+
ZhXzE6+5GhoIxhC01oicBkyYT9x1Es35vG8A89JNbMRNAcudzpWOLDObJvRc7PzJKQ5m4ZhW+2lI
nrm7lHLTEQVM11+2zEJAFFIQJfWmBVKbESLlAbgLxsqF/w3nwC7Ysy4Ell7GMjiXRsw5Xsc4MRI3
ymEDRSHHt8hQ6Zc0pw2Ee3Ucze/LoPtMFx03rsnwykP05Ce6o7savg4uZwGupuBURke2dDs33IBU
eSgliEsoAeJjYWQTr9C1uCoQ4NPK7Y+ke29sqUSWiGURV5x5tKgmWfCOJV5zdyyMWxMtSZ6vjluR
PC5rOjsQIbr7Z8NR0QvV5otT0U1KCZYD9NsclM/8hyr7k8H/VYFsU+zxlMOZCYOYS5aZ6QPGA5SS
uM+gfqZk3VKp37f2iz9dLVq8Cn4XVCoieJrp4L62g8AZejHYhBaeQzaGT1M8IaqdB9xJk2P03jCw
a7KzfZQB37u52xXZFbVF+y3tbgs31BNUlxXHteNxSzng/DLyGUMonH95UG6ck87izZMeGiiX8xu3
dj8y3YdgkZJ/9TePDUgeek4homvoaXoC7NiWvuflmiyUGRj7U2bLjB/GuBGm9lAh74GKMh6XeGqE
yMKEdUg94tMxzLLtN1TfilAdEPLuasIZzOzfGwk+tdyZeuJeBmdpmb2nMVyZJv4pVVXjthcBeRZI
cSuj91WOk7VV2lnpiJ8/NVEecymorA5KDvQETOYz05lYd0H3BPVRgPeTxtqOYOITgamavMs1bcE2
XcD8c/Dzwvx+VF6eaSVmLsnTt3NKigPr7a7k7TqFdCmQ1lacnYXwW/VQUi2pLtm+pj99Wl1JTprD
Ebk0eYGM3IDIJv+BDPWqmetOn7cl/70RcDqivxvhWj2Ble5a1MyOrN3PzVNzvKTP/k9qwqv1wLng
bWc3c7Ou3mycCdpcW5eMwV16z7Xa7QQxriG7hR5LHcyKIju1tBKu16+3zgqquE23Ezx+a2gM3bFS
yUcMnxb542JK9XNu5Z+dpoqRjzlQNqMO6oWVPZHruF0gmRNE9lUyeKlI34ybn2LBAburjHkiV3Kg
t8blTI9+AGvyc8+KHgNpm7e2fa4n0PQ3KQ3/XwworX9PpHN1Xv/rUdDryAw8R4ShdOuGYZMZk12q
loHtSoBA7hN5Op/zwH4295OmGaYHRYwdQ1ey3F/F6r49wQ+ZokIzsNcvZOBytCYjM8pKejdgkc5q
K9kAnxkt5JRysEnj5wUap9+Mn7rkQ1s1xItxfUYcSLk0WcMjCw16CHQrtuZD0g2GqF+uWDs4j2Al
tqmP7rIzaOMPl+1rfvEZeI5OisQRi90JF7oXUfLW1so/JxKXUT+18PFC1j8w3LdYG7VYgf9m58kq
y2zuMqm3+y2wdkmpqv42zJr7dkPgUkg4aYYqQqpZpvF8mqf/n7A0Q18RBQw3TkcfQ8Essg9o2e1g
Ph3u1uD01yIfPCjoNk9s4ocGUTlF90vSdHf1SYPaGy9nfm4LDSbrBWKMSAJhPtd5dkdu/x2f9eWD
+BCPPRNcjqab2TgfNTiPu2PassnXNnrbo3J9CjdzdAxootMdKg1XUGv/X+8shFC8Ti6FEwk/LB/i
YUjRA0kbuB6+nz+aOhKey48TZ3C3Ke4DS90KoRx7dtXlCfaMhFD8ijflUzU6BxB9mJGdN13jQJj8
F2RTdMeTPq9XOX7kBp71oXPq7cTVtuMOigbPvspNNX4pUC2N5sIbm74UpWbfLuMVypaFaqqv/qLt
teQtvhgK7bdphzHUMJkj2GVr5GwvyVE74oZ3YwgNtn2ctKjiuGqXbZs67yRlLUD8bEbb7AU8Z8lP
9r9l7vlIeuY8q+ACx9OD6RIoO6aF4Z4+N6+LdOTmgdQnPBXKGA+wuVBogEb8+JoaX9wDocKAmtIT
205g+Sv36aiGSr0HMOix0o9zX97bD/r1r58NwwxQ75+WU/PRhnN0y+mSfrHRRt8KnpYhto6tOpbQ
j8KmPqn8xQHVeUoasK1dV2CRgxfqSzjyewFLw7C4rsNQTalnc3bOqB88f23qrSmcEfupwAhbMLnz
fO/Z8j4jE/Mmug0CTgOaZS5gU7M9Zr2eNg9lLZc5p6R82Mg99E+0GCQvY5Rd7kyHKC5cO7laeDRj
HpPI+mNkOU9suwwuYuH9hsFy63iD/YE1gnqvHd7axbRZJk8n8l9qHYLBnZ3fNE8UmAm8qpJxJYQm
IuFpdvT0UznhAausPyMcY2FC5+lZkYNLCcVybH8sCkjv+IzjlHHS+TG4ERAZOFX2NsTJoN7FEj4S
85IiGq7e8GhPnRQGbb9Pdq3dmKKOyYqDrOLTB5deaw33zVxStlLCsKhi1ORsQh/cJp5aU4yE08ir
mExwK/mKu0Kwnjth/hpdiG+h+pRrl3e+LD7yglmyvize6TQnp6f/HTiOBjCdQwzG5we49wjiVN9Y
6VMhZyVYFbbo0vgJfCeEjJtjQTJYByEZQXIga1Pusq3SM9MD8FHztzqJQYmwOw5uZKb5vO/1/9UH
1RLkygTAPW7OKqdcNSx3sZs9HSJSeh+aqyer25U3S3alYsAoNyWreZtCQZ7+1C7HCDzpu9BlwUFD
4qISTfscXMdmDk4nmVosQfQRthd6fr03puiwutdcBHnhRNWG7pJ0C3fe6dtrorAhNa1RcXUMliSc
exFpe9TIcdOZvrLlrMXxvDo5aJfdWj4AZpd/HtfbuNhdyGam9tVZlFWyrcyQ2NVlB9jtOMQIalXa
MCa25cr2PE5fxRH6aXpXfgIF9QaSvydUKpnM70VeB+tCPPYvFiGdWrt3TWGlbanxaoUW6R/evRpG
4O+DOYGVTzpCePamq+JkzCwd4DKsk8QaQbX9OvEAsP97AnC8HOCN8TFlTU/8ylXA/EZCQlJ5PHDk
Z2LjxAtT/CowA5DREBZdSbafoU3sjsAD0j/Zg8o3xNJAf9qT+3vAaJKCdle9UUIcVyCuQUASnyAo
Xrw+61uF9UzisgwBmsND20GhZ2pTE0gJ49MmWZm0KzX9adgybOQWfErPsUjHZEa20pdsYx0vuoYB
EYclivtyO4T6wRqT0g5QvdG1qFwyqi+gjAnZGZhuj7q06bsyQrBgYKHnDc57UnPUGJPrSCJaldQG
3K4KExKOmMDZ34wh2u2od0ZKcAQE1kVplzEdBb8Wz1qoCH/93lHswAspTXj64IYJw7pqVewTkteK
mxqBfUTOAyCs+/Kj2q88WTuGsJM7vV9aEoc7V6lpj5L7icNRtfD6/BVs9SZtVvADCHqkjY6Yc3Qe
6Aw4JY4X7ZaR+LY7fUixykzYiNUV7tWZ9eOH6XpOhHoKmrvBTwAlxJIJvaIKC6xZX7GdwRu9QzE3
efb7dPiq3cvAcKBvcfo5+zKnILPUqRhVhDUDVB3MRGjIoG278qFWH5UgCNR8zjrBWkl2RU30TM5V
FmXW6j5csucXfCMUPfheEREQtOZ/f8iSaArRSg8c0KbwuaokKvW0nF9lzZTO24UgAUBKHAZrFkOm
ZhHupOumIzGNBo/aUz7kfcQQmMvNMpQ+ShgUiGE3E14BPDV/SVppdU7xwTVtFI9ykHpEzJZc33eG
jTDuj/pSEirBsgxx3rj8Q9zuMjOU2sz3rNZ09U2CKIBtjUox6d+5bqNkwb/1rhaEpYg3+LgVUIFR
KpKXHtSEPy1Q2T8SipwQ8J9sfVI1sgnIQGb87TJ0hdruf8fonrgMvv7ySut9TvrRTNXEQEnGWg4m
R05GgASQPk645egIEUaAJNWv3v0Qw1BVn73Gt68QkTgMirk+uKNOiI0pdBKlQPM4xpDeVONwpO/W
CRdiBYYVBqe/RXx0G/7AbuzGl7cW3S0A40GotsBf1NslyDzRFixRELJNtPJpxL+wDnLmfR+h7aVP
SHX0Q/cRfRphV/zJuEXp1OzshbegyNJlfdCabYbQFsi6drL7tO0ixiuKfFR5hXKu6bUfaMvEveVr
o1lpevjV8XlI4LByvKKUhLymlWkvKMkjvXQY5whzxP0oLOXjnO2waJKfQtjjk0pZLKubf/8lvhK3
OvGzM4nrDR8moYEQ+umFtC1pf6u+yKvQOrNe0S/+RJ8ruyO27hp+YhXeRpS4EhgQF2Kgm/64uiK/
tyDB5d5jI75f5YzxTFn6z6Bb2LpxFTF5gIYmUJG8nHY0G2I+WYd/emwC5uwluJPeTNLI0x3E9nby
MATDE4pmfxpbEGYMA7PrGy8Q5gbo/ylNdZEj6ITsA51Fg+9ABF8nVJYJDAVz9TqK2xXbqaFkRyeT
oivUqhLp+6wBJ86G131SkeAPbuAy8FOS3nlzpr6+k4r8zwOt8sVLKxWMTYOf4GJPRiQbxdUFyDv2
2unw9OiEmF/97LInfBywCMQ/COrtJlVxWMf/Ncbywh4hF7M1fex3xHhr7pdyQPYqGzs5fPhfegbm
QOCtR5gpbdyn8m7KxV0EOjFsIE3IKC/FIbQ8HkuQfJ6t5DbBzs0mMcVG2lGbHqn37p4n9wTY7LY9
odHRUEIqGUyUdwSDxrkcnE9JFGWn4LiWKVwX6W70+OLq1wkAljzd3bzWB6WDNdxOuIWhczUX1meS
3UT6ccWPdJVBTFx1ZRRwdfBRuqMmVe+Hxr2Z4dgC8BwBN10j0JhQeDxvnbEJUaRam46oMUw88Dsc
LllDtZ0n7i8Hjz5oYAJVAKX3I1bjmq/erwQms46XPQWaH4eYg6lkEfGIBkL99139NoRde00SQ/gE
w0eyIKPLwVisKTD4ARozbhc7Z3iWNEiTEoNbPJsAcnROafIUWoLZXReG+47RA42E3aRVFto5bXlx
1cjx5/HzKFB4+Z6HGoxgJ/u3a+YBfWCAwQE1+IH1TIMVlIZtbFbhltPZ2AvCIKWe/f8mNrul2B0W
wqCzEa0pcmlOvrqKOtoU1cA1RZXmYUR58xy6wVgyj4Q/Jc84FQE7radhTzEImi73TrYDVSy7w1i1
+t8ZWbGDgFQfMrfr2vu0Fbz+4A2DP6TFsTyrBPd69sSinxAIbyzgKbxNMx+oC3c2ME/uI4+6fy62
XyCkvGzG5UL1ZF2Hjmsc3vKYcNFcgMMqvRWAlJH7heXjGT1+nkkNDq6C1MA4TZFmzoREda1LzYpl
RC6s32pYz8ewyNxA1v4HzPIyGpmZCb2TZTXJznZsohgOQe9x+/hywmM+3chxtd1pAP1roIieKpGZ
fNFLagr5qL1KrhSN5YGDDDajruEEzh7B8TTk9fmTF45uv4Flh5XaeN+hMuo0qsHwM7O6qfwl0KcA
jYcJg7NpgJmrRDs1z5ziB1toSQhDRhGE/Ml4PsChha7BYhptQGECGAz4c8AykYdi76fcSXoCsRAO
HDCO6HpKoskSJDCP8p7WPnz+JMURJRpbvR+svE7DCN90YyDrfOeW27ZxXj90C+59BQtsRWweDG/n
OAj4LjefgJbMqhwqzUGHaEjHYgmXpDrmcV8dkHrvBxcMUoZY6w3CDUOEVk9hZSPPqHxJ2G7uNyAj
1snNpQYg5C/PMOtUQMZYgd7q66w+U8wzQ3H2B25fufsUDaVg8qPY6hSI9Trp+KXyScuoOdXFVcBd
6V2nOOIi5i7PK1bafzUZ9HTg70f0g2u7bGfjpzsUXMFXjQps1AaUMV/NfkoNYLmeyX+n3F//SdMs
achf/L82VqeC+DBYygPN3CbT5PZLOjlfCY+yqOqvtUtLIoXjAHZJYyZExlX9MM2zBXIn1Oj5TgAL
BTd3ehhiSXfAB10b3A1HoubhWYVS+2QwFYOt3yFv/N/5+17y1m2K1dLYiIUh3NY0nQ0rv12XoctP
SDKcjQmW8Zj+iyLOK9NpBRn9SbQu1ts2Mep3fAc4I4rtiRDu8ubm64okiPqrecPA0VUUlGoWrakr
cZAU5XMtD7b1gHg2B61Btdjgq5FEb9izrxZDcZP8mlUhuWtuHTNDpJvw0axNwV6chYRboh/BNPAZ
Z0l7KzyW5HDJ85mHMfn4cJDTYSk/eOL71+9ILVxnB+oWjcCf35MAkkT2chN9RRClp+l6qzZukqgw
HhM3FFJREEirMrUb7BlZyScsSCmD997IzCkspf5mGAMIHYbS6AA8+MeEwUm4tTfci/8aslOIYwVl
Nat8uyKKDYV4NyrRTGXKDk9nghSoattzvBj9Ks9SVtxrJL+VgKeK6/XgrE0WF7VUrtM7L6nmIZg3
7S6WF6koRH0lG6ug0VDc1+MCS+m5yMU8pg2ZjNWD+VCeNxTkub28kth0fiDoVwsc4mUtVulEGoJs
EbaGPGOFmvyBqE9yYSDd9bMZyD+Rns8At18nZnBC0DTvr19yrpwhKxFsow68oR1NBFxneEQ73rzA
hel/Nnk3eMCepZRd1g1hpiyUH4BjIjamoJg7cN57pRuDmE9/yxqFNj6AZad9HfvOxlRvIubLmodN
CBTGc3CnWEwU9g/OPGMWJ+PFHxo3RFCzdvQftGL4Jl6W9wnPUOpoOUwGK6E1hhNggitgrJtj4/UD
L/9ZOSLzfVkVFexFERdM5Hu50yif2o2HUr/CBvO0jM80jwqFiFWb4qu2zCE0vq5ElgvN1FB2xpHX
SJBm9dsNlMMZKNfarMZOe+HBDRLdJiDRU3s6G1cIL03tAM43ClH5+XxNoYhyL5zb8s6+nK70VoSy
IWdADbyZ3sODYFSoJfHhTUb5RH0U9MWs1iYGi+vd853SpNcdULvOHdZLAzeunmAarVLZRpD9S29p
Uim2Y8WM6A/rV0num+7XV6XitJYlUBN/4e9/G/gloU4GS0QWSWD5AJk8Ybiu0r7tNiLq6lW7b6Jt
AFy+AjNvwJwQaQmLs3jIyr/ddn3wo8LULItSh6kefOO4p+q7OFcBn4bw3lsICPAgmYnvWZVoNdu8
jBoeFfg8kMS2IeeNpiHFT8/Nk2TIssJIekdZldGocPmAtUqgci3a5XJ0ba8kHJAwoAUeyb1yTaA9
vm6Glk5wNbMbH1Ss7eZDj8zyj534XJXOkF/V+n4PrwNN6GkbaF3cLhU5vf6J7Jg3eCGo7U1AXxlq
KBBVr91e/2fWVqrZvJKfJs8JQ7/yJa29dmpovk2LUfSy/+F/rmxjzihKdGGx+8Z++Dz8lUUFyUL4
BkpHDmCW0ap8Vf2TzlfE8Q0EGsLHlzlT3GHXe2USt3UnOECWmfsA7egSBPjTnk4LU1I6i+Ig5dXe
RuD9hXTDcZuGmXHmFegGbgCH6iuDNE+YLHf6WTSRiTTtXqn9AJGYA14VLSUSJzheqNFyNzo1YL+l
zDd5Rom6KAUTbc8mCP8D2fc868Gct++92XFThg2981oRSQn6E9V0U1ei0DXv345At5GOleYodBzj
13UcSS2LkRYgmYwCJ00yhvHN/JYWgiXWCv+SaKQfNxK7hQXUx4BtQ5VEddSEB4BVw++a9MStHtIi
dC75f6yR8+ia0nTnXL4XwWJpWmB/GmJcr3akqUYUICgt8URSkNP98Ea34hp+UIKC4MQia57sbZJt
TwSAXYFh2g1t/4e18HSdeeBEgNDfp15TtBHr4BP3txz7qZ2lZ7OODJfOdWBOZtX3V2tLsq2hxWAx
YL2PEBiGI5DUAjIJiGDpy0XjPAgojjSdepCK242LLiozUSaoh50GJlfrJpuMy76vUeQs9e9ez1Nl
adB6FXE5xfeoX1rDlG5qWIpllyMXRNtfwkSPAOA6lakOgQqoUsAoAM1PQfHkXE1eA/G1Mq3jEELi
+GiN/47qAFPi2D2RirH/WiV3hW/YOZAaUZmiulA2VyNOSGVROObXKKjPScCdq5sLJ4UGn3eMS2Br
B77nfj178mTYo+1TAw0OQmVU95meoJJ9PtsBYr+Gg+mzyyiNdjD5MgLLSNnJ94SjXkRk0dUsqvFA
3nHIm1xyg11GeR9rqUqb1HJi3/dPI1WIxNRXPUWgzwj/E0YionI4cUsF8Dvw2x0F3zX8dh17znyb
AOq3oN7bDTRq6nQ4qHKrjmW4zrM14TgrPpft5IvR7JZzbDSfPtinhhdp2YzMF04wbOQ8GuZTnFNA
kxKG5QaciIKy2wglu+Pv5PkYtUkqezUCD2L2wRF0JyIB+tDpVYE9kL1aJqDDBR2IzfaT9umQ8PT9
UtQvw4uM0yMK3RpiG3NXwFo5GGkFUv7Pv4VXokGnZ8FO1jXr2QMRuj9S/deHQd/B3nBbka03Ozd/
1qdEtGWeRVIGXZQfeHdcxQjR1yzsj3z5wy8lLImYuF71EbaEuXaFAEeriqD+Nycm9HdK1+DDpRpR
+Fchi6JzFt4Eecm/9GOjZjsdluwlizxSyVZYIWv6E3WP2r3SSc+e1a1lMMwiCHDaEQFCtPnhpZ+a
u6GazRLiUZaypQGRzBILxW5P6v3jSlXTAAE5M849dTLXG169y5hp2q++cU4mFRE4KrPVrHKONlBV
bBqdjcKKdaSDeziIOXM90wAbmnmwAThj7auyS+ZFx74384dZXsxKr6QffhXGzlxffuR7C3UflQLm
7qXMbyuvBA9+YcFxWfkULU4XGlWroE/PCs3lp81tujtyOnGxC9DkOdtkslb5MwbjAsUqqL2QcFuR
R22/0laeVMwBWpvY/nBek6MEJvFzzOwmsMbezJgfabfYu06dQ/6/MKiQYI4jyiz2Bc1sfN4GpG5J
/ANrlxFJeFPMhqQ3ggArlbU4fa3UEAvr3zSb0WKyNq5kHMwro5qpM7M5xWw8bQa/YrFdBwbJSEB3
X8gM41kh8XQ89P98O9P7MbIa2aH/7TwXRsU2JM3E53VmEJ4jPzoZH6eXObuaxy/TJa8qSlmhzpvq
urp04hbYY+He7RWTSnjs+kIOJWrRa+Y5ikJThj3w8SYSSeaxE4Eu+fkD+SaQPxxSbs0mD+gm0Mv6
hiqvDrVo5mm40Ms4BfXmidD15A/5SKbzF4D16MZBME2sIEFYRRE0Z284pcw51URIcJ/5rTWXKvqy
i0OL2smHcaCtUIRCyO9LEOvcMTpfnZnHkA162vQf9pUaTNLbgF6ag3T/Ia67SRdY9g86avHiqbxu
pZ1QOJ9nH1LtyMu+Y6/1GkdALGAbCpHNF2seWju6pt8NM7rq9XIguWSjNIbfKT0xXGueH/Zfhc0L
0L+hwJe2tZ1txb6+Mdn3XsXKAy1+SnHF1TAWqqb3OujlXKQ7MjTA8SXbv5SrbFzC2zOlnvuGyCex
D9jmD65wt0n6Khb/Ei03/pckuEihkQqgbYhrSsIH4Q+Eu3fF7fJ79o6rJ1HnOta8YvgckNxGuVkq
oYxrsx2i//y10Q53B9rrglrqt43jQz61cl2gJ/wQStPcUvxH94Tg5vouADD5Y67stL5al500zbsC
I6lBPlIMzanFmOLOGCfeX3tPSEpOlU5NS3Nd/xvXh/ZLkQuY7kdEFvPDhbS9AF+MKwwYTAkKvfB3
SmU+TPocYLb7GLmohJzIEeaIYqsz7X2lSrwfOS2R76YxJlc6DyygNY41oFbEUJgq0p/ylWQnkDcA
8QdBZTRLHg3Knng8ssRiPGW0YgHWKXYoqwd5Qas8u7xsrSRb2HBgrWyz2y18Cu3ZaPTkAm3RHXo1
2pmJ2pp2AcyRN1pe1rb23Agnl4l4ydNeBsLdCQ5t2C7px/YweeKH+b/j+nP9V4YR51Ggvd7GhcbD
jseqGa3q7VU2d0KVsqTXpffok+sbQ2KpDPC2BCRCns6TiuaQv71TG47g8JO81fGmC//DAavkaZ/1
e6noLsiD6Z51c+KhwuQsR3u4n7olxRUHfFTB7sN3jsOB/uSTL0qBW/jOZT2NYCMTlyv5OV1ITyOx
4Jei8b64cB4D7FHbLf+sK7ToPPtLgzmJR1MoeGN7hT1pG1vA2go7PInmrPIf/A1KMMjKv6cUsH6W
QEU6/XAPA01qMWZHTo/VgunUUNDvVBMSGQpk5slmZLg/GvzfD1apnybA9yStOEzF7KiaiIsWDXrx
vBvFwUC3o5N1iUmqGpJ35mRFJqcoPcw3+ShJfCu0HRd/d9RF53MxemOS8wS+PCcoKa0qP3tKJ8rw
07qiMkg3L8lYkEeQ1IU8rXuUsMu6uwCpTeVEGAe2ptAJSbh4x5tuYm5CWPTUKA9jtEA5RaVNkdIo
pg/VmZAyHRWaFwl/Nvp75Bkez0iFKAH3lJhJQIePG6kvL9pwOND1QdwFUYgr7Nefs10XDMqkTmRX
SoRjzF/lrukLex7m1CTS9mpfrdSVJ3nsk2R0POn0VSF8hu+i86XPfIWpcBuECOMcKBMGyDaQr2k4
lvVzBUX8fA1Rq63KJhPEslldL7F2xHtChpYTxy3FkIiTnFRTgbMSVQiBO7EE9SXJE50jY5JKNYVH
oBcP+N8izif+klRnp3TZu5WLGyK7yanZOvRVW+cV6J69pXdPrGIY4xJPSC7B3Fd3rxg6rwuRDZA5
DG/zQhiZHxeap7Qsfc4PBostdr4h0l7MzuaR4x8MZqJk6N04KzMpVgRql96AqWmkaf9BB0xEU7XT
Y14XwHktkZCcK7HfQnBkbij/lOqh+V8Mr2lUL6/YbC9c5o32Jkn4+udKS4Wqjq+hfYIzsgUui2pi
Yg7I/FcutNFc2l+H4jx1HlRBepk8xzmSDB+LlMvOjGM2H4fgBgu+rZQGlJK6gtPSkCFhc7KqYDnl
WW3UgTGyq44qM7rOA5Az1dnO1dnq6TQG+M07hzSAuEZx8WRSnKxXQvEP/5iy1RzUHEXqDzC/2gsV
TwMjKIQZSIthqqCO8RQueiOk6wS+DMaRR50ZauoBdruUwq95ZcpkjK0zTXeeQAKZs1MNjzaJMDm0
DTjBTMdg1NDwKLV9MWuq33g3udkFlcYrfVVNuD9pS3cKerDdkWz8QhlP2DpI1HcFjTTGNP3dnFSq
xoWiwtEqFk6eF8g0TmDqNffSceeNrcpR05FbJ3m9/oCx87mAfaVaeRXq+fRElhWNqpZClc9XG3XX
F9ZZz8EMcOzphA0WH9PIB+O59uzhkgcB0m/GCX7HFU9Rv9NGUno2PqsXpWni11Y8ECw8Y3T9yIwB
9YkIdnVkpCRzVhC9gjzAZVroLsvimVyFVn4n+3rMgM3RQrdX45O2N3ukYxFfhUiHL8HRpgRqlmZK
pIcXOj4RJbDtL/So3+NCZMmQtE3LbRSRtR6LZv/Zq00S7Q7bcWGsRZG2uROd0LA47YAM7g5dJx/n
rYqfU14YIYm54Av65/8oSvMukGFGN3wPF3u2+7P+IuavQEJ151J3NjnV+XOHmy1WtLJpZWBZ1xDU
as2vZugUNglN6yUf2/KrdKJE+L5yYhsauJgyQvS5vx+ud5hYh+PFkCouhvNEjRJIbUckhigAmKRC
O+gVx2sa5xmyUrGqF4CFt4tzksVZBWXp/GrWNAEk4bSzVxesRVyc9gLy4+eHpKg2YrNc0XThSwE3
fslvvhsU8BOZnyGVn/epOAsQFGxG1/SecGru3fVfTJUfuQfePCS51TmigGStoJp/Z9iPZgB2rAO0
VyDntAG6gajZ738S4TgOhC8kSCx0K8rM+d/uyDntLUyJr3SoxdCjQ1wM2UvpAmT5bUK+JUgB3HPx
R/rHPVCTq7gsM0le4FOd78qynWwDTlSBAUa+wASYunyD9LtOSyIvzJKOIN8sbNtJjezO9Xzu+DMh
Ehu1zkir/NPFhLtffqItZ1zBsCks3EnNwAfdXTgMJtiui3Qqw/ImwSPk0RFOVWgnzizlBdP9HQOO
kzKDsmgu3KhoC8ptHWtDP5JR58haBsfx4eBRI8ML/SlFFnEboMF6QFoIY53FuI6mfKr7i7ETRSGe
Ql02KaCgnYTdZE9EzDQtWZrJP9eL8LZm3xILB/XpBleqA4S3vTxHNTaOoAIObYSyh/UMiw+da9/1
lky8ob9phLpX4Jsd1WC39o3JEsuFH/nYZ3uNMZ+GW5wRBJ5fwzj8VKX1A3SJ+Z4Q/UDO1sDeLKss
1Vmzk/diaOWnIhxXRiCHqwxNFF3b7R9p7pL7XoWiuqJBAnc1VrE6xTcDoQ9K/qyBmM10uEFgWSCD
sJgfIdEEgSUBAfBQdFHymObvi9vdmRUIXccjSDqui6RfdEdkPLTWGhqdTsK65qexoPAbGHbJY1S8
7s8amm7vqWl57ZuOjrf9hQhRE8jJwPBdsRCv17lYJ0AuBf1LAhOghcMOOu4iV8HEGEUgEmtbiRWr
QLLuLwP4UaBoMMAx5dOaAWQM2EbgUvdOJ0ggjbdlanMPGuCd8t/StCOGWDU48moZE9sAT2mouRcF
CV3gKahUTS7/e33nPL0kxO9CrQRH5wrcCjREMUC5KI4IfIMXgaTU+zSATEe+adk+JmjpkAO+EswC
OcSBW7XToaXAI1UTfr1zVE0aZgvHz8bEQ4JWWyrZX9A33Ma4bKeWya81q8tqiKOPAU6pSE0VKp4V
P/p/ZPZenGCvFXga8DKe6uq08wyGZKJA24Mf1SvTxSnypEfX6BdPTYghcZvAbCyLwbWIjQZkWUiq
wadCO0a3IcWmpr6DstGPbCw7NhkLyXVStWAw430kEUs0VPwzmYbyXxtHcm+Hctfsvbc9/PnTp7XM
wwPGta3TxpeVA+dyf59FZmEvxLQVXS7tMA0GEwkoH6JW4nCJe0Itt2U1/PEP16hIJAs8o/X6XSJZ
u5hxHL/aQ7+16qnAl9X7u8ftCSR/I8A8ri3hIdGX61rsZwTqokTZF5nLK/O8qlitR8+V5BqFHSuC
jo8b0vh3sHts/+C7nqo7BV1/ykhQk93f9vswDJ82i6DK6B8Ixmh8LqCLAFCJRdvOixszirDPYXY1
hKDp0kgBaYul8b90O5+XCLbmKDRrg2VB9tDlqKoM6/xQrS6XZAql6JNZunjVBgakGIM+8XTY/pIf
p4AgI14azHVe+L3w4GUigvuOx0Su2jf52xlRlefKuol3jD4Mr3GXFaeNrtaNO6oXJ2Isd2JHZXow
nrJn4Xr9Vz2ChsxOheczuL2Mav38SE0jSpl+Tx9q9dOqHbp8DzFwrtB0c7J0R10F5gI+dW+lWMy2
Iosu2wY+YI2QvG9mgqgNvTy58k1uy6l2+qc5OAqAMgCFhDA18KPMXEUW6JQl/Pm7A0Vupnpy8kjQ
CXqiRC/DzLWdyyxaC3lQ0u97eiSkWqZT7O8nEnbuWDBaAxoKpnCmafGKSYzEhLhUBHma+iwTTesP
f1hzxyPJ5AXb+N4HbBWmZJAZgrrILsrWjintIuIr0nR7pTP8mFl1gDKUGRxK+nFLAdm62xoAvFaW
L9zjG96xvMh9fq+7qAI9Qmr7TYUbUhNaGE8Rpg0Zy2d3NhNFcEA6sRR9o7WkJuBJEZfHQ/zHbrFR
li9l/IgGfxo3dIzKr2f3zvWuC9+D6u2Veuyf7XeuziHi0IYv4YuHX8jxSjWm1ugIPsQlOi13zzdN
8sxjvfW1nkLBtrNrvEoTQbTTMdUThXV/Hm9Fe3URNi3EUHLTTcebdqCcm0aeHmjkV3ETKHm/7tP5
Rmn+VEBq+y94gUzVIt5tR3vy/gCki/OQgI3/589u5qsW/EyyQ/WrBs9rzNNCD7hv6OsjHgl/YAkQ
RlK4eYIQBv1aRwIrK7sqLnKZIYNfZjGw/XhXWRe1nBYMnDsSDjMQbtRwkhd8Zz/RkuoGPU+OMZC1
0aosi4VRQP8eQPBYZIS/IHDo71kmqlbt3B7vHWUi7RAI3Gn1p/FKex2Fwhf4zo6XwuhsndPOsoKF
AXIxVUpNroWWHp04/c8NK5VWLwBd27iVOwwYHcEWmbr9hv2EEvmzfF6yqEIpTv8uxlqVVfO+PzaQ
548hb48sC2n+57CWPC0+hPfAchu6Z75w0LwrrCMQLCEAMu9FtTJYBgXmyNAiMOvy698gRHWWltIf
kmjXtXr3BxhjmAqTPYvSWLB2DC+4Zmm2sVT68v844z/Gbe7vgDtmNouahQiBnUEkbEWx2g4Z48it
1A5JXkXLA3scVlQoeCFUQ2k+htAAUmmd6tjmPy9Hc7xvT1zdpgP8wp8wDjGUWJmpuj33tNLg8S6/
877Y8nVGugT4fcIuxdZtCqU276XTfZtc4GzSN4H7Pk3Jyf7n9R89pY6drdO3vr30xxSVO47cAQlP
EImr6udt4WkQoudMr6bEZdAtdlcZHa0YFbDDq56UyT2TA8BlMm0EyZakqLEZgp38YR6XqNzsxlph
oQRYm0ODEfVo/9tlsbA0nw3WIJuu10ibYiUgKpsxBNBvRXwS6NBLfnskTOIS4KrcShWy8bw3yChu
HS+nkKNQsuDuJdKoZL3ZOZSCjcdjq6pRyOFadHaDgVsIXE2xUkl7SpC5km9tVJDYtFNMrLjNzknJ
ocH9iTSDWnYKYpfNoMC2mrM+YHLFsaiArzPqxavZyHNJ1W9m+tdbCB11lilCpk7eSdoei0cSc4Sg
ImZlYUwAFpxMPPtXrwf6I0Y98VEfaXWfe73OX04L5dZPyciGCgy5aT7vYVAPan7FmLK3kjoAym/A
VmA2YE2gvVA896WPvbIdvR9kEmtEpCdkDY+CEyhz+cSJC2GSm5V3a8bGn7LshzB0cnAvI/BD4ehy
wtdw8tlSYmrDPxG3wuHZJM1UZPUwdp9rMi40AQbo03ydbPm5R/vXY5/o22odbPFINMaZgv+hzFyp
GD2Kr/rNFkCdzXmh4ruPGcUci1zA3QnAi5/Pl28XUQLU/sE3B5joucLCMJ4XzMDk+28gB8rG7L4z
db+KYLPqaMpXskaRKqnwBzC6T4WTmmm4vDJo7EUugA+O7BnIt7op1sE7j59wkgXmqXlMXKqZJs3s
KczmBbtC12LBtEvOcfxPeZ7XthOAjCb7fDWCKyibs6KNOZHV4qnAB4DolE+L+TEClX5ki7Bn7xfr
ZrZdkUXZ8Wwqkuf2LHPIv9tOUjpFWVkU6mgybLhGA/pzhgrDmZx1XRevxiu0FVZRJMAFaykwre9w
agWUC+ys9OKa1iLxaL8JGniw6Fj59RZYjNTzJpnGE4CO0VI7NfFVBKBOwTeLk1WKPxA8wkssuuOB
scji9UDyPAvmqR/rK20QmWeSb8mnFz16n6K4uTV7PIpS0JvNs0ywuq6BmXNwfYSdHWsVufteE5c7
JNqZAWtjRyaLj1K81OGruO4SRwmz35JEg/zHKGxcyXMoTZkDNwGqmb4K7KdLfBZvLlJq1P0zVaJH
2lVt6Mk5sS25jgl3lPVHpi8E8jx/BClRjau4t8q6+RdeSvspBwg1Djx3MTndz9NI6Id/eXQAGJNA
ZjzPyKJ7vq3cWIL3zWq7sjdY+koqCF/xxQ0BJsRgVbSt3SjgiawbAigQmeRoBAuU3l5rWD8+8bdM
4ZJCP9mySHws9Q8MlO2wHGFp5WqfLXBfmUNaeJ0k999pGCXH1w7+xTuS4SB5n9B49Co9d5tB/YHY
E1yMA0DFNBZ/EULey6CxiFV+7cAIH02gE3A0exaLWDnY/jj+4Zfy3qR6GbDJVzNVgJ5Ohn3tc2zU
q/kxuRuY4P5G5UHBX+GHRbHnBH8iYuUY/fThBjMDxR4qBMFJRNK2IAkKEdFVVbqwjZ6m0u7nDNsg
z+2frf4eoILVHYmkidMCqKOLN1IwiRrm+CCnG8Sgv5gna2h79O6XB5yU6uwSg49KV6YjBnrSHqL4
tUcMaMxXM7XZ5CgwJsl2jbftUv3dwMdQMJRzWczOsZMd+BjIua0L6qZSEH5PlcW4WvRunXHibWUo
HpiOEmEPPMR8frO/Qgn5B6Q9CMa3x8FPPDJ7dpug7JeQqkMKwtlZEGCzmCb4a8WO93/TMgWmRqiM
Ai7tfGDdZIIs1/P9Do1habbwBGewWhJDFY5a6Cu/NQoBFTgh3WserftkUVMULqRqSk2B5svAFtiL
o3pA84gBt0p4iN6ZUrae7A5kWrofTAGueGymwt9GGCV51lK+0GtS7WJL09o0rv1Mu3G4IH5HmCOz
dUytkGMnwIXwHdEr0ysvfAilSQVInC1dYoXWEKXu7nYDq9gjS6l0ntULMmerxSxy1FU71Bhx4ybv
1VfYtqs44zueJ2kWDMAgZZUZIyglWs3GE/VuFMAqed8PGdygstoKdGfaLdtEu8R3fYjzeNzxZSv2
I9CQ1R1QVNRk2DKmGHCNoFtsjVb6M7wY8TwwgBsifg18guEkdIKbVqnBH12c2D51i3xsw3AZvUi5
I2i1VysGhDeNRKEJHcmf2iyo1e50ThJiaO4fGE75JldkXnPKyNl4GwOK64rrzZcYODNdFw323VLW
/7oJqeZAufpwss/bglcdewUCYK3ef13upjNsY2pC7siIw6NAaTkDaFwYTKQxk+rVP+ey0xxydIt2
04cswe21gyZ0MLewYk/805PCqiJkaEYmC4MPGhUgfb01MLM2ty1bO45m2NGs3jdQkAC3XyBkZi3U
BhfAS7mfdDUFM6G/lyfbXSRxVcU/cbh0vICR+zWNqi1RHj9SI3mX9lhi74ZhowowlCOzoWWmURYK
i+YYXQuGx+IhnzG2NPoA5A/toxQWh5LEKbK2n6sthjKe3gi/Q9cSepEq7+dhCFRlHG7pTBkLvmU4
NvPS93ppBYze6eSUq50YNoba5tsO3BS+eOgbEeSogT9KmWfMVhGUKgJ7zVW62VSt8B41pL6kTz1z
KpJUQt4au1J7PgLyysgM1b9mFaZTYWlXsvTjKfCn/JO1ks6WU/BO1y7a5tN5NG9rtS3AHqnLkW4b
ikU2e/QddlpEKWw5N7wdT36ue6ZRrxoLQAQLbLgXMDHSmpKnJj2EF4Sj+2gCNnwAje5sUQMazsYO
WOvbsqPn3E0bBYfuvVVw9Eb7/csVDBdiBBx2O0/tQsL9OfWr6rD7w5TmpAlNg30f44W0MUzbhl7v
Zqi1vk0ByB1ersLlyjbJFy5sH8u825PgIUwiQxxYQb7fwZOoYmieVfvkL0mZBncEKFGJFjixNksY
o06Fhx/d7gaIz9pOtx9lo9ITw9B9hecC0Oav1Ak/WuWbEpcRRLWpBNY3uejpGDBmdHUqGDNt0bQM
YCK9OzyLjnPd/Z0lG7iJHao47tqX+TQIu0jLNn2tRMdZTeRwVCWHWHZMjwU/6gTzhL1dDLvNvC9B
U37sJDHu8R/haLfjr5KgjvJqbIMlEpqK70bfMcYkm0oro6R3C3QSc6ah7Ht87eIO0H673wiRhSnJ
Ds5XsDkDafTUQME/W15yIsWxPCfVpeXreTYiDRrcEPb50OkwJtwqUVXd+mJzL57/40YDSDRoItQS
OMJ9rT8MjdDUyBO8eBUC1CvNKknmOMvOoZGyj6CBdehIWOgYSk0JKFMD9HVn7F+6TKLoAsL9VLqB
T083NWaputLGAZQfceMCs3AHqsnJLE4K+iJ+qT6S2WPo+LMXaa0V4GfDvd57smuDEet67hziNT2O
u1lnN8TosJ212Gam7QX4v90fR8ZHpr6Kz463jLlqYSfdU2oLj2QdZ+EqeqfnhWvC/AJul0WY6L58
p33REWey0/OzVjEikSrR8Z++nVgFj2huHlD25YtypZrC/ujMAzAnkbnuXtVuJzophpe7B/wY33Eb
fBXjOcCtP4Nq7Ecl1lszLWb6/+XhwaAeODd0iO1bFK9ds/V3f3TF2oB5mh8p9IMc3H3/EtL4PFA6
fjG2aWT2tQPMdYkNqRoeawTnUs/ok/4iYRXvmhmN0kVNhwg1M8+BP7tEY/qTB4/KkLht2DspSfOD
0xOg/dWet8+0JEyHmYfmYpYTabjSxVPleXDC+HsA+phFk4HjoHl/KbNcauJUWTcMmswq4UA//Gvg
pWe9TZuohelTOIQLejvZcPCcPzWF0rUAhr6oRrOf4wkN0cjU92KpXEBug5g/IeuVsJOkgFx0ul54
XdgCSet5tbBeizHOuktQaIs0QCtErHFLJ2C6RXvAmFe4NIJA/iC/269hymmf3XUOYcST56tcw9+z
3WDDh7PPehoBxKSG2DbClnobU2QK0A1mXpXDzuK5CC0JKcwi4dbV1hGiCZF9jWZ6nYVPGjNPR+2e
Ljsn1C/jq7C7cyM30kstB2ePOOsjCtc80TNKJhIYNP6Vom3hCQQDme7RrhzQ48CAzo1jX6Hg4y2/
LvHMfkiwFQtW/P9wEHK8em0wA5Y7bcAerKjqIJDEkF5ENYbnVs0W+ufRm1rGNk04G4KcGJwFLx+r
AkaOZc5AmcPiZbTh129wxZzER0cIZqapnaO53w1RgGasl/nFRAmz5/CnWxioptK3R2svW8+brYjV
u5edAxA+yy0YhRrA9EMOZWicdc1sm2ByB077XzjrIHMO1UDxEReVeaPq5lJJwPBYZA1jdMZtahw7
KvkgtTkdA2HQJduh++6JLjRYzksmn5D1OTHKHO7z+Ap7/Re2YelIQoEHjaAbR7mMGKg4cxBM/2f1
GeniUduhHMrfQLsfv5v5FpVSrlcGnkzEUjoThRDr0Qfekqq7jnuxGvF8qfS3hqnhxLidtaUGilBh
ElIwGPB81eaks/Wo/P7R+HPyEmqYXqaA1nx08Zd60n+yM4LbXahCrqXbQuwFEBX4M5spPzrHbjYJ
qG5krga9/SglDObNA1Rvj7yZXXDD/HYfo4RqXR4gIreeZiXFemYjEBVzt8kl0zIenhlFNU2H6vDj
2ZlRb2MotbmmdnoR/m/t5CroISVC5cVVdRCMGw7cN4TFZU1IpHHQuSSbMyCzwv2Rv/EZ4idStA6y
ql1x98mFoHggG+5tFtwuBRDRkSBju8CAGg1iXACBmqSIPRsKVWU5LXkH6c6rfOt1zlsFrqKZni6+
z+Kiox4DBxYqOTULaUPYc1YDndej+0uqtTBNLGcKuSnPOaktl8/YhZ2rbz7bDxzRytKAuY6Rdxfz
FJXu+C0u4ml/A33QPfZH4phjREBK42uAllCvKNLHTXQsKATJ9KnrVLp2ZTIzKTe9/nuqO8a8QGCW
L36UWzuQonWcPVBP6Ph7GLRknU2M7siA+RwoetuNoA5t5kS9yNBRnQbdTvcolD8DMbhaE/aXHnVh
0iHXQ5apESaFXrAEC/GZLd+mQNcLsfdKrdrrQnk/rtY4DOV11fzMwUCZMALsGGpN1U1WABpQ7Goe
cDYob9GDBg6mA11f6N/PalXJFmSSIrXtLE4IgpsWgVW4j4UnMr6Cg/gt51ap0gagv3fODxVI0IJm
pTkC+vNTVNxRKW71U+1YWEAAhlrUkNOgQsjiJJowZCh7hjPPqhP0bAPwmX5oJiMU3sqKUqNVrTYX
gd10UB0JcqEMsMciAMI9UxsxnyrsmhltjGf+U43wCyus1pd2KxFbvGujUCk+e0TEiqkMZP/ExkJp
P+BsL/ji5BjO7v+ToTBSZE8FpajF2vqb7Kg+H9Z6biAdC5HwQsuTdYGwT/egw5P3HYKWDdHgnQHc
Lh5gu595HBjYVVlxqxUr3Y46gI+QtwqDYxRVLdj+euYZEn2g/9j5U7USqD38z8oi04QnoEIGwhZl
M73A8Uj0NNbdZly/ogNukTHzbZJbYfHLMIRdL9+v2GnYXVHQuB9bM6LtReMJZuo0QDx37PR2PZMt
h9qaVX38my/sccsIS161I0GCjqGyz7wpLMYEREPY0HH0H7b1EslPDl/KlL7jdZMkqchukJhdz199
04xezmKvSMH+CuZ+PDwaDYvPFigo7rughQRK7N23EKdvcXEp8PLG4Xxwus8mATSTx0G0Nbs80BjT
2S3MVuHNcLrhZsgv6xTKzZr4hF4KVZ8ZNL1RqU04xnK/etv6v7M6D60qRcMIYc9XRwt5XIQWNcCT
kcGB7CSWuX0L/0dY5sLJJ8+heDrgUfhgFghqGRAAGoZFtLrjMT0gLXWeBG3JFQL5Q/Nc+ZOPs8FP
rFEA3xanc4xN0ACkGlZIhrJqaxBOJpV3Csjldf/LZ+d2yAoPAXwCsrIaShoPt1DWvDavhLiv4Vi9
Kb1N3/TiGMr2gzxP54go//t2JRLOP2pLpdcRR9xA4Uc2ZPNTD6Kxgw04bErgGbxSoMasgmLGeOou
PL0eEZn9C6nzncRZNggfsXZW9FYaHRSSbHT9D1mXblP6dMuaOFkIgLhwXEJuE+elRc7RV6bmbcDp
dzR6DGIE0pb6PJZ/ylBnU0k/iA8C5/6+NGpBexZOZawQnMFFRvWgSNPqKM+lPyCvFmDzXW5zrVCe
FU8LkjxMT+Vkml+7zr0cZRZ0oomfbtGHbmlA8oY9AJxC4aYL+b6bZiHIodJQK7dKmb7MMKtfQyfX
sxLx0AQSRs/AkAVpOvB6WbpTfGBkKKWnMtIX/HWlsDkQISSKVQGhG9mUxCFrJ4qiUtFYs4DWdmFW
zqrxkYWNYYutb8I5RHq7OF1jvhlGSBXz6fyyF8tkD6zhTP+5/ybCpmmQBeL1e9eH4i2LVkW4pKan
WHTRA2B1ssQJcfzybltD7CznsPff1AIo7kQfb0GGn+MpZtXZIRiR9NIC/KgXw8egPorkFxI4kLux
TMNd1jFAPj/5EqBVU3xFe5ZESnIX3/HfoTHTfq0pdGjDYWqI/k4qsLCJ5fPD5xvWwDtrAe33hZHk
gA0DRKSKNWwZqW1M8KQFlU42ZK/loZC9Jtv3Q3AQYjCsHkKpU+0qr+EH38r7niN96s01K5hntvQ6
AlRm1sfX0IrgidIOkL08oTxU0agDUZnK+AFwSs8oHzAsTVc7ZVr5xo+ofFrSu6OqKV8hIdVjhRd/
TfCxsdWcZpNbjl5NsvxCkNmYvIan369ZXw1+g5c3GB2vzecrfXeQv7csWx119hF7Pl9N62xFOXfE
fsKPtM+by9nEA9Zgizdg52OPE409BbabMpbSZlhujRYwjGso65167JCZuDDIwuA2dv7hA68ioQ8l
J4stxw6XT1qyJXideZgZc4apyuohg916xWpdyKOb1NusOROADdAltbuhHxh9YO5PZm//CSX/pySd
9EbP4Cd0UuRh+1dbMVOL9mIIR6u24XMxvbnTL8a0UU7L+NB+MveXLbqjGp6Jclk7fEeDOoI94xWL
CZH3Xpj9goJ83i9emvIPyztzZWuCo5ERAh1xaIzUdjWMOavc6gIszHFw7h5YCyldy6RR4vyE7Sy5
ihth4yJCmIkN5cOLeC4MQdaAschBt4HHKgYjpFJcXbjz+sviti2D6+X27UGmhzWwDMIgo3f/L86V
gg0jfjXN4cqr89Xa2kmq+PAK1aZ1XQAivf1+jQkVWa21c9EWC/WBysqYgPJABbo3wEC3U8ngTkwR
WI2F5zQEcm4ukwxLM5GOwaJ9QOWtnqUMYKxE4GkeEuMZ8kFxVkisaVuTMZC0Po+FIv31ilddeC9w
Jl0fUyh2SByF3MeE6GvOa66q5xTTgYzhWOsoAgKv03un5zJewqQ5gSB7BwAU3G5iVyuMk/RNkhFm
YO+dwijipVCB8HeJS6cQ8Ng3WWI1bgT/3HTvMMdpK6jo+Op0vlwom1oWY2/mi04BLS1omkHbuE8K
2cONmo1I2NObAq8RYZidPev9zWf5C6+0aBggsWrafmQb1ly8c/a+6I2nC/zpWDPrJYjYGjS70XIx
3QapByzF95xo6nb15/w+uW4+fL5wQAEeSAt4dEuANZRmwcyxOZQ2Lsyx89eE0vPZT+9lSHtMk5RC
MUrA7T5xCu6/u+Nzf5+xQXliZj5RW4D9bQj59LhM/M7BrDgVeI9hDlAv4L61J3BpyV78NSlLnuu7
ojSOPjUkmHhIHLcai5/bNaw4r1Mh0/KF5JXH/kmMuqlkB78YnGdWHmpR7h+jigFAIRHkUQXQSWZ9
CFn8PYowbDS4Ww9v43sdGVdOxxONj1YPW0FKyVfG9AFZtunQm/FAo0Qvhh75e6tKixVy8I4j75Cj
3ZFGzb0W9WdDD+sQ2cgeRBuT+fNS7tPrTewwaAgvP8bZYQLMQ0bmNHx48yR9r5yQ4PNQlrfnhHeQ
O6g2id7PCXubC8sjayJr2aIj5RNoLzRzR/AY20mX5lrw02/4hPFYN2i1HClltaC7b6lQDRRxjXFY
hxn33G6Zrv564LSUHAzjlPMG+doOAQZSqKDkLUP0UaXSSXkMrQceL2VOpppztKo/fRe/FZQYkPTt
xTQEQT54b31lhIJkbyVP4sIO75Oq/5b6kqgN4DP77mTLDUC9PdHlcPptY+muCUbN2YIypPlmgGWG
jAkLNORpSbbF4B2Bctrl0zyKfw9mtgy4MHp0hGDjLCu3Av+ObCilk3fuyLWpaBkfJMowDTUiA+pX
5gj/wbhcTzgHT948pG/S5SynwFU5QX1pmCOCTZ3ZbKwvzJxVZew6qk/A2aLqETc2qMohIH8+ddY9
JxNXsJXi4oVxX53HSNkf8c+hIWHbDJjCm/fbibr1DXm+j3dgqlt2ujMSbaJ9xBmYcJt/xt7LtReM
Vf0UvXpr97ydKgsEfn+2HbObKJK0j4/ZBsV9zyTap6NwIJSxn3RImpR18+dJeDLK+PZK9eCgQRU0
PUM5qRz7YRFKUO75QMgsdMrxTj9D71y41Gk0dLJfQXzDDtODrq/yu3hZjrpMBhiqT9vNihXTGJIN
mi1xK2+1lwxixxqSf90cx/vebQDt+lmUOoQt266Vy2Nt3uxS6bu8AF0qNXbWQykfCnrE4hknK7gg
tmelA7YXTyVDPHC5T8dcd3hD87dRpuHnXGgqa2or/0wyovqd69khKNPZaFUcLS+UD0MSPxDSbkn4
mK4C9g48riOcLUKEwfU6DJJ8gOpznAsZOtMAeJnqzpkxv5X2iDluLFw5Jn3kfcY/jKoJsfIx4sll
4PC+/3zxMxlYJKgpFWlI6tZjBnSp4j4dJFuRwZ4EZimwl6A8qjK9mr7fSPEI9jXyOLy6dibbMer1
4I7PS00b3rEnypMJAcN5KJ6JGyaGinPA8Ia+IZ1p8G1q5kHJycOHQ+okOjEKSaPUv6fxT1ymUyyw
XfkvEmYhXoah2djvXJZViIQaQxLaUF9iJKZfsv2TuaPUyC2KBd8yObvYAqVA05IKuYgSooiDw7eK
Rj6xrb/HwoyK591f4Cpd2Tsw30E6FYPHAJGNXrdmaffYX18JQx3ifBl0Oa8JnKgTLc+5fI1gxkRQ
Nw3INU/eyzRkZeirPm9O0ZZrGVfSCcM6FgwfryAVOuAR/oRMMM3XkFn/uuxMg/PBB6e+sQA5GGr+
8YONcDXwMZbm/LgoRVoLaxcnzXWeaNmV4RimTFoVnORvm6Facs0fCA9DydKnjQv84nlYM7a6VKcW
B82IABA5SAkUmpTmX6epgnNJoJMzLQ65qfpYEgpOndTHRtmV/dG3VYifn0DmHqdkIzYldYhQD/kR
8NspdPgnt6KBtrdRMrGYb++/7fzylD/1HuuBW1hPyq5HbQsN02hPl0rF5Cd0o6vQwr5RWYI8jBMs
RD/SZt4omIL9zFt8V1uM8TzAbZi7WqcDwXv7TK1035+q0ZY08GB68ZeeH3MCrJb/XFjMn3CkCRqo
qY+c02qanZeAZ/eF6WToBSBzT+msqj8I0cpxInTzNsZoBBWyHrHUhUXIyN6rIjpvrgORevc6PUZb
VxjOWdZ4JD9EvU0Zi4P2C/b/fhMeSajZ2YGj7IEMvf7gXPk0+e/8BRbCzPBHB3eN9/58YqNy7JpG
qI/Ypqn810hOQiIsOOg2EHnLbjugsABnWuWntYf61cHl2kpeItiv3XLmwa/1TLj7bTafHyxQosdS
Ki5VwGMmXiG89lzFw6vsGparvrIEd47k8zd5+CTePhJHqd5gg6zVo1sYqYYjD9BJEJC/tIViUXIN
aiEClFU2B8+kXNOGKcbVHA+1RLnWgJZ/3+/8/23sn4nA3J/MqAIdKRG8fvX9OQoKJviOV0vTzVyu
PNhM0PiqtQg6h5AXnwjrkfO42cTiq1/rnXD6cTF018q7TbExScXGMGiHKkcCaEAYJMMwwNl6+fwA
1zSXP6RofeTyv3olwvQ83riynABb/Piue2brPs3zyhIL8c2aDd/nxS+sil42lCPN+xxQmgdzbqiU
6egxF2NWlEhea2jnMELjPrUKXs43vyAPK3zMQNMnOVDKWiLA/Da4THIr5SD6/3C72XwUxaiBQkRA
3nns9gPOoqKMSvPullE1DIs1LifBs5oOBp8dDmtA2t4QRgquQ4hFQfMnTXk4JP7Qw7O3wDINNJYK
x27Sz9r4ENTEj2dZC+Oo/AjBuZRUO1k6q/Ea7NYWgP219yczrD/u6jVTgeoMz5t8PKUkommmjNHp
yLs4RhVc3SomMiUbcfiFyIESdD+BGht5kTM6HOnFz6cnRwrEjjZc26YK9ypeUKeRsOJYoOXlxcsr
mt7cYIORQNVSCbXgQ1LXiMc+ANbpo4OUBTkLLLXRUCF/QVDwKALUWNFZbeAKSlBhT+2ZmAZJCOEl
pOUwgGEzcl1yvoLHUoZcC14fiTDQykxqM1JGK04dr3w1mMwY7JBK+7YLhK3C3rrSV8EksjpcYjav
cjfpVD7B7PKO7AF/VoxeU1CITjbq9pdN9p2MpasxyLpKzdEpkpqVrjJq/oEakayCaCXkFPSYeKzU
Rpab3S+7oIM/eiCU+oP1TegqdD/N633gfD+yBy+DcC22QmWEtymkG/somsu4aZS7tQ1Go1AF90fz
0ksUUyz8yn8+MB02KDNLHPdq5rBK77135QzbLV/dcwYtgDy65xLwXpZ9xO5GKcvl+nOuAPZs5gvi
pvPxvFz+l7cRTkTPsKToTMpPORtVPWuC3TUZjkQ5BPQA2hh/hVa8F/RSSBhSt8ci1kQETwQKygc9
lfNSYF3NQBeP314CSircK8QvkEI5PhuPi7cGnIC3KEkUbyQ5KbcnK5Nkh7l8OIOdVJfM/8mBrYUD
alamUMUkMTosNmMrPXx7h0wSU8pbbF3W6FpNm+In8RV2gz0vF0QFiCof+QgjINCOvXfuo1zPKFY5
PfqqmnmSkXxJFHV9OUIETIQMUh04UaxPujRjoFm9gq7u4wSTVH0MTuQzrgwGIdO+cvKysfWpVrlQ
r1E1yKSzNA1N3BlroKg2aB8kEzZkEi7x3/v7X+TpXus2aRoj/cga3fX+E/UUCqlEUiziSadsCbCx
OKs0eLsT4R25BdAC0xqLQrjhPe47BvrHxbSVcWsidEaMAKAgBP2j1KsokOOc5k8ZLo/WtdbbpEHM
QUux0nbFVgWUavNbhOhiwdF7npwfZPLshmMXa/kAHMsZHUaNJIMpqzbmMw0qoe1yBpDaML/LjEVL
8x1Sa8ftpLL6Jx9IWab2wn5g/WYaPCDj1sS2ErtkNwnBQ1hgisjZdBeoQIPWM4VueY3tqwvcQ3yE
y5yuI54Q6Wz5MKAwowHH9EM+vkSycu4PFkbhvBcxirP4jXsIQV4nYTEFVpSp0hSlxps+qW2Rr+80
ASiMnKHNZBp5/6wMBu14Q2Vb9eSrtZko2mq6FORwaU7foviABU+bcNs3aRSDV1QWIqJl09Iz2+t3
iBsIAotCymxjhw/JSWGJhaggH1x8iZ4/WfhhAloxRBjkHlrDDqGUhmwJ4GRmXHThWSTnqzV6kIzJ
YMq6fm2nKB4pZkpO4dHG914Es2bIbP1S0wXC/jIuUhP8NcwDgxdPSTMFmU+XBgU4eVD3nWPrffqI
+64EYQ4KUpDD7scGUe4Fn35bGsGkLcQvKpzNLZubmqKKU/fe4A5h6+CRWAPEfFqNAR28VaXQh7uB
jnk66KI6zb1j4LLzteWWVV19VboCd5Bsf5fDZ778C9WhUn9xEAJXyupAwCBCubG5k0RdAGQscy65
l3JEKf7tVMFTbrD7rumxt8EYkEoZ0GnwzX6xd7M1+72nqnqhKtYRmYBQfWBy7Ck4dH/5oRoTHsY7
2YdRmdIH+jx+VohrIGd2wPg9Dv8U4mpaofVvXQI7uLMgEs2lKV/vZWZwtw8IrCtFmPdQUTkSZH2p
LzZrqgc392lLQl+Vh493fPgsDWPNwnGEtnHvI1Z5crB9HIovizcGZQoN8PSYwuDcleCQQSDwHHT3
ER2CdHRc0XvOxWzv93K+ZoWX+teWNO1usf3Iu5NggJo/Kpvlnnz9wQUqgoLVut7SrB6Ubl7jpHTZ
bN8cqGWfuyincprZ1Vgl+Uj9sL3149MPKjD21/9Qw9ZOIveFJ5reindjfRufhSMdAktm5f/Vbleu
aOHgHljl/Sd0L6KTUhX4S0ptXuRh+B1Xoyyp0wCRhKCSKL5HMgA6WwhdVC8cOT5HChIVvU2JNMDZ
5QdwMpfl4Z8v5pIKvP1GCZjRRyx2CKmk4WxViBALfkMPpzOPks9vvuGL5NVJ5qTp+BNnAGNNM0KZ
kXaVzXTqx6XEIjrcIh+H4ttFzE34Ilqmz5G0So4eHa6ZaSl3/Imuz7pO9z2J4ogyavEEeeekvM3e
Xb3iS6ylMdnF9T2eTNcp8Xkp0dNIDvjsBMrhZzVdE2CT/pIM3Hnv1xJNpUaTRuggsx6UxMZ2+wmk
SnBHX7jfh1fc/2/l+XXSan6RhGRfIqKWlGa7K555fIGHYjhmPzyjyh4SQNR8n8ffdmZmiQQOOT3y
lSl8rtVnNsLwyvFf3iX2h9KbJfcTv4y+O7nltHRBrOL7997Q+T9nKNKTQoNC+sPbmwstjtIp9qRb
NLADMUKIeBCRaHLTDD2i7HrkbEou8diYXJdWCICEv8ohTMwzBAhOuWhMeNsFjJggDOOEPabtGEUl
zJRlf1WIHaq8/UY+MjNF8MTB8ZiOoLCACari1WpDcyK/NlTtrVxwAIySc2AlfMvdUDq2Ncjx3qDG
065yBO2k8HB9O+dPeW2KNbvrxfITNj5GQCsO/UJOlipSq6Y8IkhEVvlqph5l7CEW3lr6dCuh8/x6
fF2XTXyjJZIHP2U2isMNUx7YCpHK7qgxmNmT0P0bd7FDl+W1qB13JuGXlon8yiWKmZVOrwx2fHVH
Apm9u8qdTmFU/NM3bd0wRsOi4WljNlTTAFVCWNzlqYyZZxc9YRmBYVKQ70VQOjRcxltRDilAye2N
xQ2JKyfzuMgciRpCsnyjJXZ32/UlL6WQYhV4UG3mRJCJizQJpWz/3SbyAudo4LsIlWkC0xI2zp5Z
aMMNLlhZ7r/Dr+pEFHW3VgTT7Uq7tPuSVGbvAUqrb0tHaYmL6adbT9mjVrZDOW5cDnNBHvYt1q+d
wUEmtW0DbJKzpzzUAh5IB+FHxb2yMBl3U1ZklbcgyK43MPkzks8Yqfh9cUVyfwb+jYXCLE1d4Wcz
wv35KvURmDq6syNsbnz4OhvAUHMyYwXjLaM2DA0Mtey8GPVURCbNRDkWlDhnoo8zPzkFUgrzMxhS
bZ27fuVcAFSl6bFscEWeb9+KCqHeoAQ/IRfWWt0BiR3b3Lco8LXkiZXqWPspvEJbBubJfM5C1Cyy
Sgt+L2j3Vpe2Cl6b0wd7JgQ6HByPYiH3KuTmJdHeqfuwvmVqZFtcA1TiTJRubRtCPD3Fo0VrSg+y
SugjbfJQWwh8B+piH+xUirtpYwq43BaDKwKsTXebC2kODxLAwGvH6tui7p/DsZYTO8fUYdVlgC9V
hhlfOw0KwjTPvQri/i0gQO5VzkaIzyE/8PKtKDeG7GuHDl5b2461WEHIKDo+i0E/M4q2awehGk1S
7FjwBrODyv7vUftlFoZsNHBirH3Z1UQpzaPzn6yihO1vRXbsuRdR+2cjJAbmdaGN92Vr8wgDaey7
nbc+dkkiPzIA7GCWj0QLs4bkNoeGEXxVNSki2g3FFZAVX68a2x+9lLbMiwqaecC/OkxYnSRD4sb3
hTbQY+PhRTUf6ObeWDWTjFpYZGyobOhZVXo0LvEZkJEk6Y9xfKZ0jmi0t21mkfoxrjru2LXQgQoH
MDffJ3IuayZBjmjM35vjRZNXQeQk5xR4SEolTtj4hEJGSlR0rAaG+moi/DdBJliiu1m2DgP+KdVa
Rj8Rf+W8svxgorOuDlMAV7Si7He/O5ud2o3OuCh1MYNiFQ1vFw6Le0L3l1K2jn1wgp2T7totU05/
H/s/C91RB+0bYFRvVQW4U1YUes77+xe5V6zytuFFf+eq4nQEkL9er56ls3FaJtIih3ADu1pIYqHT
oPqERrVfcQbWFjLPEBwiTWsezG/Pgj+DN1do/f4Npm19JB3oRbOlGDmev6T+Z49SdzkrLcRzc+VW
f7Qe5yzPqALgiCWlalfV+ax50Eul9qQaJ4j0xM9SB8t7uniryAd7n9th0yGZ/vPUa4i/ZYRYIb1G
LSyq5C4QHKMT3JqiZlr8DxzT0NgCsV1VZ+KR5McfrAW21oO7SM3pdMD6kc0TfM89qeLvgMCnkTHG
tJyLr3voVDaOuXBaqhG9zFvAllrv7dcLg5RAvBuHo/dBZapbZFz+MV09lMv+Y7NIpecxBMPCX6HF
3qo/0qUsEkXebD1oj7QfViUg+lfW2zLEgdkpz2m76XVFYa1SRxP6MiueB/hb+bEmAaxRP/XHFV76
4dU/1MdjWxPQUj01VZQrzFdUYEqBYGwhOlq7Jz+qVKHPoDUnsOZW0Ekpr7j/c82SDnd1gGE8wYYv
5306T6x3TSdbO4MwI6VIa1QfochKx9u0sDjwgbTsogDCtb02qJPywejecUakK99MwXyqxl5ggqGQ
bPw3Gw91xYZ2dRE2DoYdWCglCd+eSpaaHCbgYb5AkyftkR4WYRmL432QwHX5fT+Pebkq1Qwx2nVH
4M0lDZ53piUCLPPyAdmPSP9141D0BCCiPIA6LUTGoVFh38AH//5Hum8KCPQ7AnmlTQRNgix50+2I
ycA00Lnj/suVGMlt3JfR4PE3N7+jQQv3GFODlDVhbv6cWr+7HDJ2OrUZgJTAQdO/2HCLVSXwscMT
oJyZWmNtyu55GavSg+ZHG4OIaJfTkYKB66snYmE1oaNlRaLDv+UW4h3tVrbhVUhaBC58+AFxQVSz
xaqRiVijRRSBZmZS5XBN38aJJ9wvjWPFsOjxaUouriZeF9W9HcWjJMjbXp/irLnapt/WTfwuzeqy
5WTpTiejmosCAMsWvzlswxv7reQOW+y+uk8qf8LbIZZXuqR5vmg5Rlo5Ni3cwXSICTWzbFzYuzKR
pAxlVPBpKUmhlt8V3GuSR2lGy4S+4JF8Z+hb9z23R6XrtPxrZGSQbCGfNbHCa7L1ZeoDFRku35l/
RgXwIzvXSXkiyYVUnJUiMCa21zIfW5u+ho/DzhF1gL5/2OpfToXOwrYdy1NV06PxSj4elodHSTnT
oOLGAyo2kvqp47a2/coZ+TDW74lTWJxQuVedic/OmIDvqXzobeu5+cCfgxhrSIE+bfzRQqx82ZdL
Du5wMh3Wi0nGuf0tUThxO84zSrqtKvFqJuXVf83O8JR0VHy5ZWLIPbRFzRhV6RKFMs74d4xyloCC
QdaRNNctmQVVjJMB/noJGiHNiCJj0SA0eur0/7edk5GLMLJ5V6E851roVAo0bb7V70j0SHiBQlna
gL39cPqwEcPcceq8xSNMOW8DHBRpN6ISsI+9vDEubBz/lNEFwF1tYaRyaxfyCz2J/8YYqNJUz0hn
R1w/wb/OLjKilb1jS6RaCvQwp77uTGb64WMEk4CDDAhP3Ro8Uqi1RsuI8JI7fmfFU+MGdpg1BPZF
+Z095b7+A4q4VfizljjxmTEPXJtEQlFzImP6C4p2L/Tig/pI0Ft+HGb0ccIgP7DPACJ56QIgwZAP
U3WqXLCr1IxK4cDzqiYlKKKZMoJ7tKH4W3Ql1dikeML/D9kADSZdrQbe/ZWeLziqYL2DCDMSvmA0
gBIOV0ekzjOSHenMGiiGV0n0n+8X5b1L+mhoCoSg4rLc1Q6avkPTmFL5JAdlu/ila6HM/mJkq9dc
xU5okBVYzI4O+NDI5UMq2PX6EtsfLEf0Ejj+MWRaGfuhv40TNweme7EmbwFIm9IPDcR6gUDyAsZr
M8A9vk9ZHKZWxaMyxV2AyzHm3wEewXgCAxIN7YaDMPAsfe1amaAXDO+T57ESpAPCXhjsoILvx28A
kmnFXYdn2Y0doAyU750+z6UiE6i3wBMnfBRBSCaVTVNfI9pX5aKCkOf+cljIyQir3zXXe9grW1/X
HqybPIAKcfWPzrJfIk36NiNt7esLOSgBt9NATIzToNjgkwMxCIWY9/Cli4lenve2nCReoYmRkb/d
L0UXPlUtDzTVOM85WenSRaVQky41jUmVIMsPljR46zTo681M0LIqVZJh2hvSjUEDdAktFTAVEkt3
K5c24bbjH2WAHNy0Gytn54QjhRkYBpSZIiK3LTRxFlcHp5SMe9Cu8p6xOceNB0T0QafHbd19eape
ltUUwiWyuI2CElHnEqNPZIwJcYlgebaFzJ//K9U7ydG7CovisNFxQkhkjf9euQnan/VD9EzPodwa
N+dxPnVxj+FHL9bT+UvGt3UPqBJYP9kVpLcyX31ayohE4wdguXvWzvUTaRB51zywYll8tjAQ3V2w
2SNMHjpvFANu/OoIucx8z91XdnA5P7vciD2dxdlFsqALsf7Tcpisr5ziNgk8aE09vE1PNMs+Dd4I
7R/J6kimkH9uUvRaNsFdttMSJWop2BgHHBnznUwPQeLCG+kFGEHYBbIosF49fCizVBHQIpOmtfEU
0AFEWPVlKrd6frfhLwNOaa/LIxyXU+bsE39XXkfLzHDtIW+z3fdH+tX0g+grz3YAGsSSJttVO0Xo
hXr0ClDHtL2ynunBmaaDIM6qoR8/XIuoBE+6rdBo7a5n6hsLsCQWe5RX1KAavKcKsGYCrOdDs0Rv
6xKbJjPAtnNfrO4/lEZlkW2hAQIsbeO++h3KnFEWBP65IDSuElycL23Eihr2r4xfPX1V6rNtu+fP
KN+xzfrpOgzviD0ZEnSQLZJP3xcD5TclvsnbOxlGZ3iDxS6K6iZ7d859uoCUr2pbtxhk/3n8vrSt
Gx9UyQNRFMui9s6E81sX8CO4Ex3RO1qII4VtTlwJM3vmJZpF1KOvN49Q10VpxK95ARLUorMvtyR2
8cG6IhSS0XEcsx2RLlkEGYh7v8Iox6QB9dTaG/YR6jINrCqxWOVWAJYOaPo1/pSv2zrGOHdji5Ef
EoJK5upujY316SCHbaqd4BnwB7gTRmrZkC+k3chjfvP/AGJqrajVIMn90q2rPSnb7w/hF6uYHnsU
EEjnFpKJ0xx8PKus8C50tnL2+dmYb9uB/Kh5N+XJMZ5iHZPpvNzQ7G0dMqRBMJUGBnZ1SHGtLXWM
h6PuC4yD51hA1IuSqjxm8ZIef3MPF1mpQVib7+L0TAiTwLCSShkb+IoPHWy8DCgEWQ0I90KLwZQd
wqHCDx5nkaHsXA+xFk8Sam7nFZbmrQ4V14C5EFS7srFppgVZfY10Vhczwrsgl5/miiWTQpu0/qzs
MQ6NT5fwyR6NTSvm5irR5rCad/2heOf4i1mwTIb7kiC+sbWt5Vhu0GABPTRfYiDRvH2qgcWUrLJg
4si0naBjL8CjCp/QcQngLvvJ7Psffi4UBPHXb9vYxIhJneFJcmSfSQ8CNBiTC9RPgnSILtq5l1B1
/sqG7S56NaKDh+ev/yivkOfgNGhSPsBya8sbFgMEqvd3Dxe3hpys91FG3kx6SoOunI/nOeY+oc8v
9Q4eIvphM3lVaoXV8Ov2UHg11oYrDQhpl9mbPXngP3sPgfGqgdjKUY5WWsAXFyYt56Rtk8n93+Z7
/LEbQ4GOveOLjondR0qWN+E4cvTdZ+VYByBosjXqNRl8iwXg/PW+lqhyf5h7Rjr44S6UEKzzvNyd
24DjQVrFgtdVVJZ515xo0VbwMGivxFH4WETfB6ATXmvplBlgUXYOBSO7MhIxTn2rxYAn7RY3qjLL
PLeuVD+7CYt2VujBWldiza8pELcnxJWxYJ/RGqQssHKY4jjXZ21YcAtpAz8x0Yjs70X0/wsUW3rD
IKTqRrThey1Sa16Z57uGXpF7QZUbJf4bowr8BJJifuubIOBk+2d++Z9Pl9xey2PFjqaz72zmq+bi
9/BuoojDF31r6KYosR9Hqlre+oSeJrCiS2HH0D+YTp3oB95mTqSnRKeG43vdemsSdH7ngld1yMto
G0UTLgJto8XlgFnzfuczn+ldRHUKrzKUY7aPIh8khLvGq4kiuKjA3P4ktXqOpMI5RwxudzpzIOiy
P3kRR4Qb3rqMTk0QtvwL+oeXwjLUBuU8AFPzDQvUTtQsX5x3BF2OITsLgLVLEgigf2Sw7Q5MofWC
LP6YeMdsfMCtmBL8aVyMfhkVhP4Vwmm5czkQwvm1sMRonQvlPkT6IF+VwiDAMyOrkoGC6BEZS90C
l99B7erGG7WiFx+6viH2ibBtboJ/0TtnJYfxhbP6q8VKwVA+Rnpk2Hr1quLwC52liWTwMNXw6G8r
H5MkvEZPYUi7qTxqT/1z8zxmdMcjzpAfcXX2yPJ4vHBpgnRiKdFU99ATz7q9NLJ6ZrmF606Ei6cy
K33r8qJ6I2bKLioYeUGG9rtkM23FrXn29hg1pyzEC4kp/uMaeGNmTRQWK8W3jrlLXRGokPjx8JTr
Vs8trDzWHYja+DHFD1vM6qkJnNpVujUD5LXYj2UlUBByJwGZvekn2zsWPguoAMiErHlnG/WBeC9F
c57ZuUAnpTYUV5QhWYWZO7EiTjBT1bADrHAF7/Rywz7dKrzHZ+7gri1YPZr0WRuGm68udzKxlnvL
KZ5cy2uAnGAZIvRvssK6Kwawr5eX+YTbO2U4Mn9pj/DSDza3mfKDtRpM2Tsr5zeYpg9RlGr8IIqs
dKKlq1FP/2wwOADQU+StPWK2PHgv8FHMsUEhWnbxc2SaqULJTkr/GQGnIioM8tn13i0py2j/0w92
hUDAY6DOUNMEAT4/yrNE3p9HR4M21nrEegILRW4aGGEV+EdQAK2InHUfqLuUdgURUf2QZd21/p5c
f968+SvnxVTNqq1hkBveiEwSplqCM7yWfI/j/LvkVfCr4BhRrCgTJsHu01783uZqRFSWGT5ATZqW
wht2WLoZpNIe37edSgLojIh/r5UD/z+QtQJORF9EgAgtIe5TIHKKfcDoIfsl/7X9F+f8fwWt2vt2
VSUv9CEdP5OVhAdpyGZPlAZ1uCmPLA3uZy7mLJpVqglXiWtA6p6xw4UFB2QXUuZLzAmrkj3SudVk
3Yu274J+AGbw1lcVqw2RQPgpgAy2nQaUDG+c3GOsxbQ1RXQb9fZs2ml6oC7yH7mmEOZMbD2jv2ph
piAraxN5uwYQpNYGCmSkHUb8UsCFfMRuZOyCi6CpUg2NlMy8opcgJUsOvQmWEZYVYYXP6uxv/3j5
PKt3fhTrukVTgOuzCgrWLYgVhpLOkeRDEreOklvgoVreSw07KVGOlP1fy3znFj5sIpBLFf++GruP
7Ytmq6vYAuTvJlfL7egbo+9KIqIEYqIk7TOua5uPXTW6xKGh4WY1kHcWvk+TTxOX9lfv5prCmYjZ
PzjLuPwGeiLs5eLLHP8+IwWcoaDV3tFhoAlthCMsur4vWF6PI/3J40GY8k7neOjIIIUQa+b6g4Fr
dJ+VVYUylo3fEOYIP8qOpG/P+u1u31JyGa5HX3k48BNJ1MYktg1huelsLlOA3dvJArYjt3gL57hF
Xs/ZxJ8SlfPh8EQFO3bCZCyE4C40LPuhUP3Fb78kdkiWKLzEYvNPw9ppJQXEUZhPRk9ULhLCR5nM
BqZGP19a+6iGNOu5Oq63CVki5b8/14vwsjI5dvGjRP423tln0G4o3DZ8zPKJzbMiotQ+LjxLpjNy
sYTi8KvQQfr6U61cJv+dGvez0b0xtDplWSqZEp+wschTKj5jQMC7ZVVgT6sdvekvBETw7wrjt+OW
+otTVSAeyMuIPn5PFGvTk1StVXSU1d4gfKKP3ZE9lQAM4kwPOWKoLSXBM1f/J7ft9JgaDkF2tK59
S4EpQMvRTr/yUYB3otfvQnvDxXZ/4Rxoybb9zeomfuwX6QvKhpr1C93/mINJEEykpWRPi7RUoCLB
nTelIokUWXAhzpeQCy0L/go+Toznxu+16JKAblzdweuRlue+bRhBHrF3vjf/KWm64ewEZcpHHWI9
ff3gkiwklP4Z1zam2l6ZFKZ1c9ACkm3IUVq58lqb3YdVbpRlA7b+jvn3Jaf3tx4pvIkb14f0SLdl
lVNVu8j/rkCYqSpbmbZwLtm9edbRNUJm7V9WyZ2YY3gnxcd5YS3KzDx6ReXeOV4rTZZzQA06Fgio
4NQBBcV9m4WGbYVG5a9eSE+ObW0rb51i+arJnHsw81ysYrI1W0ez/4YGmAQ94ZTEsJZTg0dJBBjk
KN0iN5IYHDpwAWNqHDO24MdnMfZZhE4iBqLVILKuN8/ZSeOczmXi7MALGfBh69nzGkNuBVZ1KDLR
rfWWKKWRh2rvVHXGn87dOoCBUeFdN2EOIn5h3OuXGcqk1zVDYXJfXdBzzs9KtCnVeMnPhcGLRAkd
G9WnuyWR68thhBFjH/ztpsIErJpT3q39nmXUYJlK0yM8kWDvfHQjtB/7YUzCVvl54DbWD2Hd3YG5
NUJ7pUTJ+Ksn94k7H9FOPymVNMPvR+64PhQzCgG5XR9KGpl0CvyDFnMfs6CNApmtNo1yJiDAgvy8
TeN1F9eFVl+4jG9HtcHpjV1F7qCPkOMzg2aWtq5qYoZ7e1J8BqXWYWKRSm7REAznd47ixaskxbEZ
ZOhe1lA2C8lwAftlt4xBlC4/WoA5xq9Q9RysYM3VfOUD299/kBz7IRHZOxLiNDLuE5VhQGaaRsrt
3COcrkYVFccD0WkpWuphfDF3jBNCstthDSJpz+EZHcCtYpD4Sy5BkhwVtINKn4B6jgg49TQbv+Lg
3FfWDM5RdHtbHkRiZe29120wgch+O/4hKqVpkm85qxHfxxlDNNC407BQOXvgHmn7yCpvrio22qcS
eGwaywZXcXK5rqKWj1Y7UBzhq+LBwjNbEHpzWFmADxTswgU/hIKrNGv+GabOwk8+wOaeH2OBdHvs
aRjjomBPDcvGjMZI9MW36LCpOXgnXW+trE5o8iLpl2Poi1etvfNU6Lw6ASqQd2N6bmxRkIfl2GGD
SltbTU43P8c6x/Wh313+mtY8xPpFeNwk90UJexPG/1zxxis1Jnyrtkr8UNCu70D522WzJGeqdFu2
Es7yhr420u9gDe1of1T+n/oWdq3/e6Lrkk9n9aZT8MpWhqVmt4fuK0s7A/WrkIyrLc5AQINUG95r
MD/aDZugcUcmbx68iQtC4MyZvDJZ3hZOc1E5ZkFJdnkJl1jyNjwdCfd4q6SeP3GsQcC0gZy8ws3J
RxvuPGEIeSH0rPZ9NnSVLpleXo593rNMlVObaiTXBVQ+Ci5aAtKd4hZ71DAtrAeiF/EwaoavBDse
USd13fV8dIpAxVcjHebHXjithyJFVS/ZunPE9hWvi1cgzqosg8JjZShFUTuQH7y/e0mIGVwA4u+W
K6j2czjuUy/jF+MRR31ddJdJZv4H6dGEfoW30BYER6P36gnj1SFDNSRUE9DyEwOPG5OZ3lw+TM28
RFkoVoMCMp9wRq92tcgMdSbuEBGN+nRi/ug/R2Wei4ucLCPcMhm0jMYAO2JjUDoJa5u+1B/0lsOh
MQ8NiQRtuXGTdMlIa+HVIvO3EmTBUVo/GmDSeZV6nL8YN9B+4lRZ+Y/EgykKkpzm5qQ8EER1i5YP
pWChDY8DgwuGxLptuxJI2EkCa8qKkrjBPKA2Ommzr854SejXgxJv0vpBWO386BuNGV5K8NphFQve
w0VHxhZVdPp3cQSA16dMkctcoVfJRYisXBWlsqdKG2XSGFz2vOaVP5ssVrCQ9xAZlU3XxWlc6La0
2gVOD5FdcENjjChmpUyFLAPbDUSzx/I6JdPOyTSXkeR82CHDbNXBXEhwjOUi3RFZobR1DNvpQ+3e
peLHiYFKMEEgDyTx4wsBurc6BdoYEozmUT/K+5bshJN3z/kXe8+Xp2PHNSrYCGNKLcGVH8VE8xS2
gI0UGzjLgYRvKEAtw5/bk2hPEQ4/9GtEOsY1AwoZoXqkQ2oi4slgFG/5uulwwTmsTZNgSjLB4tg3
cQ3VZPwmCKqzjXnqWWfrdFkEiD+hvUw10yiRYEhc2t4PFu2aMNj4D0HAN02TKElPaoaGntS5o/At
NPTV8iHqnP1u79FuNjTMadjVKanAj5KqM/YSA5Hr8n1Aqgzd3b58+Zl3CA5TO1x+rZeX46Ji7KCk
fIo0wUi/jgrcyyBLF0155AZXlMcJACRDDs0DNjOPky6OqERbU5tDNGGA5siKGCrYLlyT3vnIwDpj
IvX64tccseJFrxxd4LAlJ/Cbrpp861pAqFm5/axJH+fSB6X5RbUANGrCmtXDZv5f2eshhMDIZ4VB
DUhkvZ5jH7ANiP3EGV+bQamN9EZZTWcYANHvP+bmrkrvVt7hS/NGwUNKiRXZVJLdszGab2te4Kh7
3U7f5+FS9QgDuZnyK/IZgDMhnJn+59XKw1XbgYj0lYhuDbDUhcrxiGGUcVfAVhCYRpB6dc52+yY+
Obhrzj3Oh0CvhA2MyjCHsJhNFyfdJth/eJarF0jPo3RlR34fjJPi6XeDXv9+iY84UEjiHMl947BI
7nYZW+2Z9A+KctA8DiLHL5XQrVCxbVVuEUd7xS++KKUMjWYAJb4j19fmaw5bY7PSrwbJARR1momI
pfehL3l6JKuAm9um0KU8TPpalt0frIFLf2G5XQ5wGWo+9gvFRwTxstCnWADUbIOcjZdfJBg+2oVT
+QIy3kuq1sPLk/tabAwT16JOfKrwZIituWHuoKlQhpTGsx+zniL3czy0896V1hGCPmevg3GKLMjl
Sx64ZiZyvEXnYipKOrNdHYXf5VbJDHEDqNjjk+LhuFs+uom6HLx+L+50inVH5E6VSK1KFH3hwG70
xAxl5KXgCGYDqS2bzyqLVaCTRBXBoq5C998H3z7tnTq5n2dt03k2nCR946wSkvd4YGKNXZJwiIcf
vMhwb6bIUJo/zyhfhnEGO0s5Q1ydxqta3Og7dBoVd4ARo8Fm8zKhzuCUbAJb8H5dVmvKQLQjzg93
QXAT6d6KQ0kYWqbDdewIHDYfKLCFetcg66OJvwrQg3USmn3eUulkPymg+4gcqAfmd95+qaqRVggU
3CUSGHiDW5gWVyBBaDfL5BMsXCBqrqSCKNI6vRNRuaHTC42jvYKHvtYM5mGhId6h+4u5jfzf7MQ/
xCkTH9GTQEpX9kwawRzhEyAOYP27HPPcRQh6E22DHDxnoIrx/OVOgjd78WTTlnDSSxWMVBujUnPj
a99rxZx2sNPnFjP0qIr2EHMiYzgeM9US6FQFtIql562zkRNYsj76SbAhNkhaELRBL4IcC0qzA7cR
3RRgNTLCxqFrh8nQzLeU2Nzil5AwSSUmfvwskLZvhHY+VgzkLLZHNY5up8eY7DE4DkKTiASIv8BF
gHmLkK+UpMQxPcUhnMfvf3GYJKlzp3LNxGFJriCXND24i2HPHvdOYTwH7ZK1ZdbS2ZwkzfPUpYzo
+COIa1A9vkPSSQmPgXGMYCWIbf9ML1qUcFdN2Q/eVtHXZA2eLWMRXKZEq4YpivLs4jtIlwYIEWRE
zivD+PhUN4qu5Uesypw4vjhAysrA0Mf/cGcdAIghSl6/zmrq7Rwxz7MEOUZ308kzS7SeeLRYTemO
8+2XASXvoNG1j9XbcYYDfhd8LY9emdlsfUbIAbxRnWNkYzXuPyggnWs2I2oxQl/mL4cXRE6duYlb
XnK0eeCKIpylFmXl2Oj2MEVut8IxkJz4bu/zyyYse535+kq6WbKfYaCIncLpxRjV28rWJzeM27R/
nTYsUDDaq+qXOEH1osAD0zYG44M55NI4mxNG5ESrhJV9j3kzbn/iGLlJ7d6EJArS1Z45EWLOAq4R
iueH7rSPg6s08Y721Z0aZdiVZ8kP+Zzf8vOGb1zJTtYrpMpPeVKFMl8hV3SOGkCZT+B6OVRttQIn
LsWWqI5JQeHCsEAFFdurB9miLbHreyfvBseD7xq7QUFAGsFzFcCgrab8EAHF7grdPP5jqE5m0vXN
jRFAnhzkbXf+394fHJXCNqjEwPmCuyy8T5ZT3R7TNxfB5JSX/r6a/rgON7g9iuReOQ8WgpLqdVK/
BBiT6FNwiA2jK2Hsl88+UD/JKxhRPlaj7kP6aAQ8fahd+VbYU4OW1E3+cbqcfIl2gbyMfO1LRsI6
6UynQdkJv3Fx81rKxOmi9R5yVULC8XQ7yUa1LOPPp7DHDEaHFh48zVMzLZ0XqAjjTdWgEgSqMmDM
htLPlQN+IL6xKbRaydcakjODra8MyaWLCEKjtyyVeJRAoP8i0yOKqItHBs4C09asOqAmDxaier06
WF2jZX4PvZ0IX8CVlK1WqlR2Rnuilo1rVxTKDWay3YCKp+j65QwqRqPsncjEPLfZgnHhq5IzdkHm
/dFvHHpxQej4VdDlJYgDS5rwIpwyh3yEibu3D0uBv9ICLudcGFTSg57x15SjzY2+RLEFdQ1ZeLal
eAPsjqExkToa0q2D9LMFFWWHBZDSBwIAYGV3LSNyDO4Q0BwNi+lFeepJ/ciiY/W84pNEMn73AwbJ
GZr4fWIR2pqS5zhnlUjqLnoQAdCcqAKUhwVMWpFzk1AWED4/R8hKtaBsTszwr5wjw+6xnC0VtUCK
64j6Wp7vgR+9+6kt/oLyxc3jSsuzxqU2AVysH08ekCrX1S2WNdUxdTGiDsEmVSA5DNyw+VkFHp+C
EwOSvZAdncW8Hn9+61+OlORcSzOI08p7UGtMn6lbS4XCAq8JPC/VVHgFRUxWb6gVXqQd/SbvyQiQ
7sb4szK9P3LSCHf2vkvhn1xofDddUalI/U0MZyUVBJirHHAmkV35SJ8ak+amrMSkvH3i83Hqmkss
AAV8JRddNxD/NPfYbdKaMxBDVjGtkuUX3geChKViBIrBB6A78SYZD/l9/7Nk54F9nHtWCIcmez+m
hR8QgFJwIP23q9gTXOUn3ql17QEgAxiSnCZSlHO3ag0POWLpGre46jEksokA6abx6zggT/4l0p/8
KGHr34va+DenLJVRbkkLFgtAXRpSYmQcBbGwyB81wCVVg1AzmxdA5bj1mx0EcSMfPKysHUmloulJ
R0WHUULfxz9XJ7T+vvkUpzEbfU0cjOhQJPvZxvuebtHhky1S/WtXAYsbAci/1MXIP43QRxbGFX4H
BruwJ9jGtuB/HBe9BCdHI0ihxt+O1BXuCFhDy8+lIYWEWa26PwYWr24D9Bab61suq8yMM0ZXXhFP
vZQ/LafUZdMHNciRgnysG/4JezpoUsax86zzPJZRLwhpum6T0MeYuqUH4TwDVja8f4Tn4I2Uw8BT
9/z+eLRQ/toYLVa2NcGWnbdP8WPHNgFpr6d24hU106DfPsfrb82ycJU8j/bJRzTM+QAopUGcNPS1
5Hnq8BVNOhQa3uZ7PRlUPKqI0yAbRRpD8gjnRtUgikko7HbxbybeLaQkHYRj0IvOveojCl7uiy/J
SINqcgLD8hAeBvms+2z9E9Zmo7rzMFeyLoEgKVDCtvODClPaEKG6vzTQ1vHCOtcHtBg3jgia3LVB
ZqrVQuTmbOFt/+4XpVeGfQy1nRoxeOgQHXB/3kTm+gY/UuUovpuPyg+vdDS2agnm0kvoYcl2DI0Y
iOJE2vP0OZYmUKdzc4ATJTbipJ+r7qH3eDEhMOusaMSUpo1AKnKKjB4WVYuLhZ61JXMWfxSJ5Zi4
PWLNAulwQN9uoV1scXYAjqpPcKq2SQblYv90wTdWzPw6X8n79l3wcC/tUhFrDiMhC03/s3LgDdWc
77sn87qcvYyAknqUxbLw0RpaY5a6V22tuCXIYjaI3mvG1Fmt2b+Ku2hCna+NUVBBYNnfQiPCL5Jl
NekLtGrfl4FqJ22KBniVAxAfULQ8hA6h2doFxVgH6KzRPWhraMQICzc5Kwll0ssUeywJ5oSs8ter
DNmNtGLLpcRG/YzYkilfiCI30U1Ramw5V1v/hAiEHOE3yHWrFP17fFbw8CltlJh361uVnfcHrOO5
q2fWIuy9KqSCaOWp5Mg6dVFJsYzqTmQhgNkT2BFtIKZkb4+1rCJwoQDew4BWYI6sf9lqkbfy/vsV
xwI/w/9oyECHAc0Rel55TayAO1tQ4uToShF0jCE/qe9m8sjwk5MKTcTUM4stpBlwhceOcnw4UpY0
rePSF0u8kH+hmudgyRrQ8DJBKue2hGF8y6B/HzHM4v8LfUs3ko5RJGUzo9k2OIwXbocqYLxfSEi6
LFFK0pqZh53VGqqK5r96Ov3mOM46kxpyn+wJM2Eo5ndqtazHVqbgt2lt07VVmWaFYZDvLZHlAc/h
EIlaEsaVJaVlEohTQNNxmhxK+rVVoLEuxedLwZK1bJUIjxQdr1Qf1fG/RS+Ccu5wvHukybJaLYGY
5fgOVmpEYq0b0dFoFCYuGBOTc61n1Zp6OzB5aKu4KbW36ieKdJN4ETtFkrDm/CfEilwrijF7QQYg
DL098JxEv1dOewzK/QCtPndtlJKU3AlCNWxXoIfBN5bgo6fLvQ9+mq/FySskvDEkbNmB++AoXVci
N2vNopEE+16zKt+kqOxV+K9ndHGxifqKfj0XFmJShaw3U97Ca5Kp0WUspBQvAadiU3KKny1VYsCq
fko9etKYqA852ue9v7ViM3GnVapgXQAfMqFCF2XEO5L/FLekGkufCJS3CQ12ik8zMuceeQyrN/pQ
KVu/bn/Te/3ReI7yvpywCPqAzzUIy8FkOCWW1AbrOs3oT1ZRWdQP8UcLehCZUdCJ3Uu2swHOxBQb
KWX0ClY8HiqBi0qzbMUaTYNXGSTtQUMhXTxUAep7VPImqtr0cIkHjbyynpEjup2htluQNBcsxJBq
06JQMsunH38doE2VHyJRT5ODxAdx05HDAjiW+1Oq3w1pyYjmJTFCfyL7kDoMHvs39T5x3go4byKW
yuXBtE0GXDoME+XRqe+LMSrodEHcaK5vVdcja/CwvL4IM6a8Povz4FQIWXgs8cPdRp78xmLPNw3k
/PDKo3CwWFJcNGWphnjudcA1XRmyHA576YdHJCVP2BDk54MAIDSpplzUoPYm8l5Yb4q6yR6qr+ud
fLvD8mROkxAOkLBqv/cCQMGFiaGpmgURM0MX6YaFJUMNWHS7G+k7l+892Plh2kxHRENEAiYrVNwu
fzWF9awXujh4qsKVY5HEerD7cXAEJVFIWu3H9oPyLxej05h96IIs+ARTzCDmlo04Etf9BGej+HoX
qjrfrPqfyGfHY89U9Qyjr9IFuGeaS9lqaSK0DJVuWdeuPm7oD7+LSrH8UFzjc/VBRIhEKjYArTbH
PY0WRGlA0J4g8SrgxzLtp7BXfNar2i+MJgt6Y0SeNWL3nEsFd5cJ8XogUr19ISF+dvMPXzPIXjaz
eICeyU3C2qNTVO6CfjIFkt7zQ64hcNBd27V3HXbrR8/5Mhwh0VKMNqk2p7Z/n/DweXaxBSuvdzd/
Kxg9lC+P3i96VgxIvI9MjNRDsX62OdTJJikkxyJugq3JgnrGpnJJNhtlmCGb44MB+7JC9WsC1Pc2
STXaNL7qU6C+JOVmla+DH6rcwrJZiDB7qYSZjdR/NuGXjvMN/hsRRCTr9uI4YaH+b8lMi17tAlq5
K1EJvcHjFLcKmyeS+sbm7589NDkJ2Pd3tIlxE/tac+F2e7g+W9NMmQriDFAwskFz0ENx45LrGTZ6
DjF89ab+xKhXfsP/ZwoY9fDkL8dCDPdX3wiPW/0LWEq2aJRXgLcau1rUhD/O1WRLqMO7JApajLLU
e60TUtd1lfwvSXHAbLi8U38o0s/WA1dMEA/DQ3g1SPTJcEmP7S+V+x1NEQBz52xRrXcaH6Zcn1wq
hCoOhIf8vTCvLOL2wAmP1A1U27uAKWjyc0XFv17XcFDVdoRPAXwEK8S8HoXu6bOSe3dHRgLSGt8a
bvxnadazP33n9IVbYJz/nOE+Xn9Mwy6bj1mR1vg8+LxCiHLYlx38P8/ybpkKSxiD8x0s+mh/Pdfb
CSKlnHrywr48m3O2LLXhne20otSYhCvD2cISgNaWUW1zqlDtJIQTSOzwCVO7aCIIZb07qheE4V70
8sQGiHE+23uV6f4SrmXFYHz+znlNul4po79V4Idln1lXuaglkDeP1b+YGJypeCgeFgGdA6UeeOfT
Zn617h/NH6Dcv4tGIDue44cn6I9gv8zU2Y2ws0rJyFMfbaWqpqpI8dpWT0Ly5qoHERw/8s8QHdkC
eaFQCyLWOpMB49UfVN7HK0QQRz1e+5rPzNzSMjqm+hiaiRd01LU1ssVGcgiXqV9Z3+BQM/IjBrGR
Uu7OJ5PqjE29/Qbb1zN/lAfIqkBoQEDP/54whGMWRug1c4N9qv6ORAVCqpqE6Cl7pJRw7gSh1gWl
WhBDEyjpZaN2NyuHM/2uwq5EaBvgLvxxlEbegMrN/OIwGz9edyjlrceONKM+Sh6keOSW/i0G++IV
9v6/hr0TzOh8cw9VmAkCXKTpdXKkS/CbvqticP+6ChxDWJphlnaVN/461p421slXrGWQcU5+qLWs
EUK3swQ20PlHr6iXlYOItEZS2DvGa5jjZl6mfRbCDp9fxOuv2oabbz7HpB4wD9MUqr7hRnsuNST3
076gTtzYwVZWBgk3upfGHjgQcwbHx1SUVSIvjf78yTv0CnAqDHDZuROoDZn7rkZv04r0T2Rg+5o7
WyxgDMSsZ5bn17sK/zaLILn503h+HK5ZlUl6zYfvssvvyZz4M2mQXy6afrzO25RlgKR3Zgwl4V7E
n9AfoYZ9oC1CZanMvL0rp7uKmv3j83gA6NqQCZ0DivDyuvS+4pHbaUUSjd7LAEHtGA3cDnMTn0uY
J444x5a+F81/yjWd7GB+d6az57U5lXiyWsm6hAvaJEOjykFfm2MBBajDaE1NNEvhX/ULqkC2df5Q
tTn5gBJtKosA3UhDkPurAaSWcRB7iBhaQvcz7JqlADwoDBkuDWUNVwXXqQ70MICSpnVgi66UYMAV
pgIDYEXcMCGM+i+7fapFQMrgUysTSRTNezen1W6Ydu1WBZr3x7RoNbnxNzkJQ27jUUb7r8kBO0MX
MPK5ki/bZQUGkEKqod2oyyHPH7+1YFd/Js7ZMDvWJ1/O1Ezk18arlh2+xtjDwG+Gr3kouNONJqCZ
O8Ij8TklX10AO7E1H4e9PsR65w7B1z4fcmv5fP0MW3uUvBN/aB52Tsbsn3FqcH8MFsHhQMvUbPFL
F3HQawGJQzpoECBwWrp3ZCvmvQ4nhkkTJVZQCV8uHa3o9azeATEgy6eaZFqjQE4bsK0X2fmOq5Sj
bUBtfa2hnTpubN8joqMe/g06WheCXZ0MF7GODbUxkyDdb2pEvTYkNBPf6d2P7c3dezeYAf18OcEJ
helVh+EUJCI066arPYNsM4+6AKJKhqKg3LF3UEZzp6R7PX8CBBI0C3cfvwFNdhct/Nad7qymqNvA
3s2Iory79L60tFFBmh6LSr7Vxn8TnNDK6oK3fJl+kN2+7PE1q6mOb3lCud2EpwZ1fY75EzNDUg4r
36McSIqeqm59WX3jnyg5Tx3/4pqEHxW+kVHJEEns/yPnB+DNy8V3xtu7aOpKRTgWiv21VHS4h4XE
S/NH9DCsNddmsjJ7NZskKTytp+1j6MAnCFlNo1mbMoL3d4mLbYo2rlO8uogSLMXTX8k8s7g62SjG
pbjtFO3O7C0fkOu+i51ptCnSgcQekZi1JSmprZ81h6UtQdntbFWr5Z6hNYEQt8cl7GAejewza868
aBP00V0RaEikDDinzqCyV9gDjzHdI5mjuEfig7ZkaLcb8/W2Z/1buZkoP8w933qyGRlbzFDD3zbt
xtllw03Tiv8URuy0m/9KR6chO4i9Vt0YlshdRZ8yOtMAPke+buy0RkkApqObtcTmyjKrip0kGcUO
9V/CY+go35rggIY9zRWbzkdqDZ/5SWYq5yLJPVj0zURjdQJpflcMFWzTGdAGM1QY56ejo7zEqf0Q
KxAxk5F8GlNc4I1/mr0YNPCeLvdYZfjHuceT0l9VrCpgbZg///kh/3S6wAtapC/paU5YF9gOY2pV
/xxkhiQTwPYEO7sgS+PvgBN8nnaiidy/7WrwbIcE+LnXwDNCvWvzpEHhHmyZNaeN9eRtqnFfpppT
SXtPP9YHW4RUoN1T41+crl8ovc6KGijwyg8fckhXlSdw6zwiZHraq/WFG9JsB93YI8Q4A4o08AeO
rtkLufxnSCR1A5eF2uBe8q9byuLNt6EJe/JD/wwcxFQ9+tF3BqbrhSDv6MoH5OI+991RNMvgJ0gl
hveu19qscTPB35CdTl5idVnn3J9zuPm92EOY9GzvqrTNpb2OEKWoZwv4YBaSneAr7yDIi5GUefnN
RNA7XW4csUevZi+Y8qCO9bZ2y983so8iuOjdFJMEoUp1r9CL7rrMZYqZ9sRscLGInfXz8EKoPW1/
bwnbuqrpvpOiJOnOeQspGSRB6zTMB14V3z/S/7nVMDDrezWjZlO4RjkPAa31e+nfJwy4ESqNCzhY
XDJRq4za8TpT1ZRlLTRuFjo6AKJ0QQpnanCdS8nE2/5S68yrsdZcZehc/+vigGACJcyOt1oRGu3T
njObJ4LI7HU+6sgnSQrP5x7aWgP9SaSZm5a8fc9DeWywtb0x7eYx92nxOrsE2WHF78FahxG3bkpf
p+7sxzXJXnlefhaeV4ZPpsc3fbeYPNJVl6A/iSdHY1pIudIJOPEhcFvP1xNw+fYNXRcaBoUT9As4
nrAyq1MEM/K5Kl3Ty++jDOTY8hE4FAqRw9/0+4n8TNqt2GM3GccOF4WLzCGLeQcRxI4d48C8lU3J
PCyfTs0fAhpVlZ0H+1RaL/k3kG+BQRfqGBJ/h7G557INQ2/6gyci6prwFMdyFYq/eZ/s+9N8rOgr
uHwBW/Uq1XoLyHg1nmYy1txbxiU0a50MnPuGAUBC0cGNLXnp2y5i/Dylg+YI/D/T4dJZsw/+JZWs
BtkkOD6du7+/UyxmyYDfzUSo89cKHxViwgtEWX7iMjTrPM07i8Y0DFPnqUZQW5/mhtrIvj0okCYW
zyyGen0dINjLgTtbROH2uw2qw8l+jo2aEiXH+QgRkbFQiJ2CxViS+gEeb/ciCADkaXUd6MlwAoh9
4MbDWyHeREkoRmiYP7VuVDXhmGGux1yvWazu0S5tJMZx2hjE2e/tsLdujUFvLwSotZEkM+6Pk8hP
Ifnx/gpMvoCyQNDaykU7r8nsQX1yOfJf8oIQTlQWDTUfrztiT6iMSngQdoBZfw3UOOpIKLXBuqiR
iglHbZlwNl4qkbKiwefkRYD16tsyjqy03GUg0FmGZXWmSPfCTXfkZX3rKLV9M1tv+V1QBD1x2lzq
jFHLNGC2cW05CfKxNNlB80FLTdOR1RVWvzsv4xoDIalDag/7OnrHIbgpQ509NaiqPT7QwZvszYuz
7oAUxm7RyHxzgj4+kBF7A92MSrIwQZgeQzr6LjrB4Y/SqGXrZqZp+/4BzFpmHo/dI20b3JNfgiBI
O9tYgjDq/EBrwxaK5HSJHZ16vHl88u2FMjjY3M1sMoGbsCHeY1lsFm9o5UYvIUZrobpehoZPHZM4
GDW9wlwuAFsF7UbjxomIX3jTewBbGnlcFWSaRPTXKb5EzKIHa2kAxjRToTA/7KGLEwqmfrV3XrYb
TsCr12ccIj/YYTxUDoQCnjcZDW3VLaUwGVNtfT80qHNcT/TERUiWogH82MasNnTvkbJH4/yuvmSt
bTTZmN/n0LgThzBZ1+97yH9E/IIQD2Uj/pHF51dsutAdK73MedmyYq0VW3vNQjtBB/o/MhHlKkKN
Ewb17Zv3gRjL/3DNDpFQmggNaATuYHDVh6edJDb8StkxT1Kj5XNz9XHuUgWucSnaHpzQiykGyzV6
kSrPc1FriwgN2o7hzgvwFDp32Uldo8K2HJzz/2ZHeUa39sYIRraTb7ohbMML9mjdWtVNUI0i7AZ9
+3vsK7nMrVrJuByzgl/vHVijDpUMVoWamz6iLpeW1W8mUS+uEdeXGdoIDnoBuygdvIUT+Zal5eiZ
M75rEibtxMKX3HJS189434yjGN/78Hb8WQyBu0tHfQYhpHvzofCmAYf7rCOsE6s14PIBIeYcuydk
W+4MehfE8glGSiq/ipqXw8fJ1yu1cwwoocbyFoUd9dA56GR5njH4WfPGBJJUC84+TKqkE4bjlR1q
l9F6u7nPgVlyN5dzPEt3U84q8P9BuhBGljk53ubsxUyYsMKhpQc6+6hVWmyUAL1w/ZVO30bDVmls
44fC7ZjasEvEb2kCTmb22oZ7cymH8Q3w7ibkx/lkjxlEqEPTaQoWvi5T5+/IcQO3cFxx6fxr/+3U
76A8BDN4d9RgPvjFEZvZOalk47VFUPnDX5V56jXJ/JjdWUQj5NforKQq7XWnma99BrbA46G3xPMT
mT+5u4YDz9k7SfberKBBbQcWW6Bd3JhtZo7K8aVfnHeX8iuc0aOVDSla9ul/T/5uMq97oAPA8zbK
pDOg8Ih5GYTeNpaxGrJFhGHR7dYhhfFnnsgLWlkqTap3deuzlpPd4JB6RIhxKshnpWTc0zJCb68x
/r1k0T/ZAaxCLx5F2Ua1KJJ5a1iV6+nJx/Baerd3GwZOp5+xrd6jGVqzmVSimmcAePYdxFUgA66d
x7I3gAB1MKSp1Cx57MBmsrTDVxGSE4CeMNU4TWkQFT34Zjbl68ebPLZKltEx7TwvKxfVeS2s56pr
nBE+BIv7+OAeeFaeJmnZP0QrNwpFRrb4wSwriBQvBj2s8TueTqpuktdgItrR1TZKDaKs1ndheuNu
y0iJw5Wg0WoZCH6YEzp3Qcn35Dpi4p0AElpsnQdgtOU7dvLZHZLu1T/uKpvc5+RG0+yJUhbPalYT
IR/T8R8cGpArk5/+MT/RDyQn1FbbzIITtCSKWPH2G2rFeBSL4At3tj34Yg6lhOzU5C+oA/Xm4kBH
IVp34vG1xJwimLI9QqAOQrhMEKEA3j9V1+yXsjq1AQhRZKkI6Eqr0DVrjDb4jnbsBjJKAjyp1+fT
8Ex6fj1RW1bUq57qPp8ggBbxAItVadn8XBAhXjGEMJ9k9o03IWaQtQdZx9E1hVjGTyM1u+ZHodQT
ZGKcydxZEoV9Ww8gExySOV2LpgD65O4N1Lj++7C4/HiKwEDak5A8AgTv03gB86xZUNK83rfj5Gfj
6I8XcQkI0ZcAYWqAzVXtgn1bQAfogALOG1IFji2Ejifz/MMK/TjxEbp6YiQlR4jZnPr8rvtlBKSA
uzUZ5huMhaNpfQFZLkMgnabyA6RDw4G/TqHpxXl4K/LGfT+HbnvzNqFABlIqzTqSJ2lLXIZkbNrx
392Xf3KY1RohiW1sUZMU0lN8v4pDTTwWGPxoAyYnwtTOigzcb87p+gx510j5QsIuD9FBmdHNgCLM
8k7qW7ourGMlXV5GwCTXnjyd94Y48/vrNFKTJi3O/zlO2Ho5fYX/CbtmOlzNmz57oiJfdLl2tPgv
vwD+UukwpXydZvT9owIXk1zuN4S2laLigReaSLanLE6mA2Ei4tasvYxkwmKETMz7RDfxic0uqP66
rVEgrcL3QY4SokWd1/mqxOfUX9ETOCOYfx47zNfciFyz2hkIKrrRYezNQ24GNXcRGkyheZ4GcLNu
HOo5Z/cgDZF46g2YEGYVxxuYrcpFHAX+4wr147Pr+Trp3C16hK0Fzytp5chiwsUtuhCw6fN3Ooph
DjBV8Iw6OPBNZlmZ00XKNCwm9708665z7Wzr8ts5MQ6ZmzxFOll7LMf8LlVLj2VEASrOQZuremSN
VqJJf6hsZyqU8WNw7wDyF2l3Z6F0Il/wtgGzxTtcWULgLVfBmiG+2AtxxDhtyLaPIpBhx53fWpBM
EWsGDZx4zkxv9iFk1wm7JsPa2RgEt0CixEKtNHSyhBTxMRaGy4Li80OPr1yzt9B7LyuB2QMqJxow
byPFSJMT5uA/ZGF2DRI2XgKlL9zrD+SKP5g45rMeukxfFB9gr9X/P6Tu+3SMwkpuQsihfljihWO8
uZQtdd0ULkOM71chmmRjyEEiazVjBzduVmo5jPQRGFcNEbTaeSbBtA5ZOydyBE5iX/Q8fWIKkwDb
/2i/Bxf8lyxxmy8/+kb1IGelW3TOlaKl7U7pvDTtPKO7iXiKfZNNRV8nOPTUoGAKF8OUeo6L6SOd
+lFyI/58jDtqyJHEw7o8wezuDNgK9/99qaRl2wHIveqQOdhSf5U4xeod1dWXNq+lST1KjxxsfmrY
+a4kGLe5ce6vJAl8JOkA9N3DCLS/hPPtdoCf3LQHazFnvlQ5AuRjC8hcGWMkp9d4n9YG5v4HPjH7
ZvzhQ2xVqG4OSHAtyiWJr4A75FIzp3ugJk4wOvVCws7CZNFm2DsE54PYvshdg68cBX0qyuzzZZI8
Gdzuj1x78Fva83ZWCExOuMhcrUF1WQ/hLGDKdcN299MaYkw/eK5LbjyRPYOzaq/9NZ2ABSVXbsmp
l7ZShxBPqevI6A1K9WajsNX8C/zptxuhA5MZVm3uzBicybGDK6dy09kKKZ0qOdrokMC7bLKljiMr
4C8Brs1MZDQmHVF2mREAFUadF4NjoCeWbXhcQ5ffnKwH6bPKr7cbmynr4ycQRmtPmXZWce/5eAus
aRbckscSBpo1LrpdNdO+xCQ8p8SXAnB2trNL3qgJKqsQf4V4tEnf4C9xBa1i+doZ1YPhkdXvxs9a
OdAySz6hpZG6VRnF3PFayobc+8znVivbMilIAmOMW3d6vo3PVFtKhfBUHesdcgG07G+Bsj+t31qo
Ukywzh3vP61eaFCgEDE+dTyBSBqtG4A3Y/5mQPo5P4ZYuTrUjwNj0B9H76bIV3rv+zGx9GbTLoVs
JsEMc4vqUeXBgS0B/brbffnHzUvjnRraykaNpmoChAkBHdGc6/+cNi96HHMorXkLFEJ1gxQl95X8
s57BZ/Gfb+sbxZPx5RdOBgbAGYeo6EJNiM4jRefC05h9DhR7A2GJbX4WTpEbf0aE8Gsw+L7vtnPm
YuWNfEpIOKLMuFTyTS9b7ZfYuwgSYAOu8yaY2Wo2+T+h0WIQZKm7ZEZQko7El9SWCxUm77T0luWC
eLtO+IJwY6u8jv466zR93cjibiWgPM3xWKN5V6qc6W2PyZ+iLFX9xIQklT8pLl2iJ2Rn1ZXnnTHm
0XSgTplVVSjLDW/3KzFmpjqYThR6khJ/QKO7hI9gUh3/DjDDKlWtLPdrHLFn6DfUFE9Y/k5m5y/f
X9a49vnQwBMcpTRkXQU76LOq6El4Qa4S13GF9LiAHvXHCEwinqZHwz8T5t5FylW65tzJhrNwBIxt
YGXlVSzTjC3BijyLHTuQIvpjuq3UVnK4sh/FzPcEXXs2I5rdzVd1sKg6JOjAVY6aFJs1W+hNds55
987+aTnzVIwiy1IFanVM6dn666+cBiYii0syCyMsZibQoETl+kpg8z5kF218EzZFD3cIuMw/gz6x
11HJBNPLHBzr6xwKASYW1CDAHSa0p9fF5yCSxiKpTfnB2fVSxT7G4Q7qlAx3FrNhWsVWXaz22dZD
cXrgzjFOhvNY/jIXUmTQTr9f42qyKolqQmd0PPgwhHkAzrMgSz/grJ78Y9/D16q41E+6Vu9xMU+W
HqoocRZVxSK7rDQqM84nYYCBeuJXgkeYf4EWxzCKmB05ST+sWdNIUqeO1glVU1WVfJd9lPrFf5g6
9G61SgTriUFJyCm1OObfmHdo67R2UAB/dTKyEbGpZMI2PF4FZI1XcxTrz5MUSpGQUpM78bgg73KS
/Re6utJRO6lrbjxJg1zReidPh8Dsl0R8AA9vmf3YhwOMhk0nanWsRAMFdQ/LIaSGTZ/cSOOhXi2F
5s811M/4dz5cOiwjB+N8H9BUTA0NzfwMq12zCN0DnHOiAQu1JrW4TpHBFD4p5Xxn98j4Gv4n7Bda
zaT5KDNmdHhKts+Qiav5QWUCAhuCYv8g31ZFchlQhMYC9r5yxwSbF4FI2f3WjAbEiruuBTXQkTJ+
hTLd3wfiaZUZQyI13D0ys0qNJ0tHfBkk0hLtsUttC2P8O0wtGIGIyqAEw31a6dS0gGLkLqJg/BlB
l8ehp6DAdjgNjb1cOj/HbwiaxgNiQgoDWWl7gjSYc1CxoqnzNpAZB5usf9809QxJyCJQPuw4o4Y5
SydBDwkBPKksgTpTZXsOJPuzTp32snIKavPEtVuUZuG4BXzO2/KcjpNi2k+ZHFRxRMQumvMGm20T
OQoSLBhWlUZnBjQw9tREjOqIswmI+21av4oBm/40d0kK43N38X0K/ulRQPV2E4irRdE7vw0eNF2d
Xat56eLk0TaxUAcOzrRCnksFqWuqTXxJkN/pFTe++IyiBYSTfDpTXb4WFONA3AAxtLqYVvLtljX4
/+ytr92dk9VoIZ/y6spacpdnwN5AnVS2WSa+9c4SCaYIfhWKuDdhu/5gxuNIppilrYF12K3EUiXD
Jv9rx8oKwLIGC/X1SJTrbZFMyZ6lx7J6pGrRXhDrFx3im9/TXILAAdeuPggVAnx5Ycq7QULip3hR
pGatQ+qkg9fL3gvnOqo9OaTf1pYUxIFI54aSmhQOyGNG3Hwt0RJe3+T37UIbvR/vzWzRXtOZHHni
DeP6x4Pqi82fc+9lpz8DL4lYSpSiAhDOGKcmkrog81Tr1ShDxR2/4OO4WGJfCys3hYvAWOICXP0I
0w15+cHiPD/4UR6W3XHcq+z3Q9XYaTQq0Q7qzwjIM0qKuD96LcSdWU80hfI6GZ+9PjeLuZetoupY
o6x4z7shXA7BfVvF+0eEOECYjrSl5YPi7kPkAUKyMYT8n/EVSyKLBP6t+LMgvGHhYb+bKaDUU3V/
IHT3Cx8T528IER+HjWi8qycIw1vtWaroZLHn6bHtXFzJeMx9tUBT4I7Twq42zGNO0z5oM/p0VqJu
dpG+ln5XvwayI6uJtgCn6Smeklp1YmNuFOyndfHyN21kpCGm682xI4j/KCo6JYPXQ5YSfrffR3Ta
dAgOHwQ+CJABajCdEmYbkp2y7bbxeh0y3cJobBa3HD1TRCyeqkeN+YL3onGEcBuqL54QlPl7TN7K
c4psE4xn/vv25E8Wihqz96O3wsEVjC2s0TryB9fsyBT9nXmPc5Qjm8YoXFTuDle6aCdF8E0oQa9n
J7T/DGxM9eS+GnmuFZiQFlKcxuH/XzVnZsv48JAoLlEKtU5LS3SfzopSmotiKQ/34EQAJqeY1ZIy
oj/vcvtfnQvICCNovBQymcdnDzXk0iJBV/wrl9FPaYmLc02ncuf9ws78d0959dQiVCFDlBv2l3dK
8tz+uwN+1WZIN286I6HTIVu4+2Cjl5WxI3CrYJvQXadGlcbBA3/D/wVzb2r4Ex5WGKMJ1wiTXk8J
rN4op4rMgjqpGiadIxyZDiMq8YKbJ7C15j95OmMmud0QRiyzF9S85TDI057phoavMMKjHTCgfT1U
N1fhRHNbs5axuZkko8cVgd92Db4ZIdiTN+Em5SX94OkyiB30cVN+SxeEoMqht56IADExlyi+BDYQ
ieXF+hlv/JzzRUi2FckXo6vUlCsx21pE7ehAg7wa6riosx2AbFSx5uqMeU8ALiHO4AdPDpfBjzpg
wFdsnHNSqWELce/VKz31HxR3OQ5NySl83MWCmkrdSFgeeAsWexR17R2d31sQf3RGI/2Ur4SZ/OuK
VADL9De3DmoWl6XiVpXtaua5KDiuy4av37t8vvo9b06i1HNjYDsWn8No8/imCOzVevkBKint56CA
oAqRovOivZhPMLxZ1G96l4eOLj9EnRmlrdl6YDSNPrYqVHcnejeNfb46ttoWCvMOxB+rs0eMulRB
pLVnoE6dwgNgBs/qtNbzfH6TEX3/Glm2Emoi+ZIxzcHf3GpY76ce0QupXyV/HQjAOgxHvA5LKOlN
9M14OiGDuDCnzyaul0BqAJynkffAXwKe1eBxjhj+SGvK3ByjXZIDk74SrXGOXxzl74QWEx6MbTHr
/JSQc+ucqD2RmZ/jojUw3HK131eKpUVFLOOQqN3vHeL4rkLsVevpv0Ch8ekBXGnHyIRP8Gh40+P5
Whv9v3azR0Uu/ItjWGlifkKIusbyjZXf+GHfc5ywJ3FrpkBDLHoch2pPEu9erJT5uZjjdPhbFI0M
j3oGCqfhXs//nqoEG/wucqr1nEgLAGRWjem4XLmed6kwBRJ8dCWhRELZrHFTWW3de4jqy57uyNSv
QS/XpDc/yt+dL5OOef7UcwVJRoGBPaJA9IXhm8uO3B45FgMdQesSO9vx3Myi3kDoilda8Jnh7hFK
1YSDJtxnrA1xJ2b576G7k2SHjoExNmHantKTqn95qx1aciH23fHEcAbdAoyWzAAi+SanxD52+Zl4
QAV0lp+64XnvkRm00MfKtnZkkMPTvNtjRWRXdyluyB1zx9QkPnMJIqQjIHNilq5seBz4qEU6AXui
BaCVoLQYNUpX2SZYzYSe3SDWYLMSm9zwDLsLZrU9hVJfPUPStRTZLd4LVrUY3AU7pE018szlJvOI
E9m8r5GTKRP2t09qDeRKaUdbt2dQ4MbYsv40aVTNabIjAY0P7TnnzWK+uMD+w5Wz+pcjfJj+Ropi
i9ze68GDZmasPvj0djrk+LTQJkbeD1kr4CrQnz7I3FcHBySiaEI52R/LlRMSwG1mtfTa7aB3AA9C
z2oaV3aaUa4FiRqYZg8BHmbgjlEZKGLJCBpzPSeGunquMhhk3C6PNCGrSDOgzmELkPW2pMBiM2qi
sQfGYU5+WL8IZZGJ0ofsEtJ4uijsf+cIwbdt8zsWYUVyokl5bmwTzdzID70enmBOarThBuWPbNnf
3+tJGBnVKHfJpsPB+6VhRkiGh/XljZQLk44wDXzS01LunMSGqqve9d+RxoU8DhkdgEClGZjijJwY
zfHCZDymv68rX9qPl4RWvGX/hTL0x8jMHiiDW+zrIzZn8BbAWdQpS/oEPhWzQmYcM5L8zg38AHzt
qg8xDvizet9nYy047YVjZbISHEdepJGGYznhJZj8dGjbQ0gCkhKufNBfdwDgoeDBe8cV8uPhW2OX
/iqNrdebI/tPV805zj496pNIdmDcY3Wyqqhol8ZH2HFiQn/AauT+Cyi3dWn//nsE/gltAFBHa/Oh
Ij+ahzkAwi1KoMN9mBspWJTY7LDK1NKsuU/MQBdBhM0Mu++vsxOZLxTstH1gzz7hi9Vq7PofURO3
oU5kJ/3R4eoy9VfPPw/hQlXtj2s0FhBoufmDrMohYWGi+8VSZ6Mdg7S3vrSSyQhfE+rYoh2x0UNh
uUnA7ekqFBCLo+KeoBiHKImmUctC2oa4gL1/Zd4q6zeSF37h7ZNwtAAghllVfHs5melRAagZu48Y
m3wn9ZZepr5OG2yCGcVkGVqKVTZmC6OjK7roCYyhVJrN3fPgkbvjT6ODV8xva+R0F7vxRG48NhfK
ItA7F8O4Jq8hvC+Ex6Sq3IN4Fwu9ykj/GkF9UbARgCG/xRVZo7rk2iCa6XTruVGvfb1yYUHDjdrk
sO0L+awgtU4jpm7ZP5bR6jRpWXUR23E8oEdXxIHy38A6vY4pT9NLK2nFjT1ISqsBsvJ95hWt3U/h
muc0/D7Zffg8qBTVfTkF9K4fLt4Czaa4bUI6VyD0Rn7eCpCvV74mEJVS0SlbYQFh0YRdFj0RZwv0
2mblKh1RuLv3Ws+0J+faR3KLsa4HCfdeZEopKml6v4plMEEeSxu+zaZqPwpTw4g4u4FU1rqHhxLr
qF5dFxSkSI9hZ0QJTyNHtd1ZNtFGxVziswz5EALforSjqEbWQSlbfcjdfnlmqjmjx5JUIVKqF0Au
uSmYr/vtkNWg2my8SV3fF69T2HHg5oNJ1JDM1RyC8BmCX/NkGQXuON+jVk0ld6HUciG0YTw/IABG
zI8Ui0DYQKi29u/wDm8z5/P605EVRBotMIVoLemp+HnzZfC7XQFREaT5kiA31MUMbhTlZSCtG7Qf
CGniFPdyOzAOKOfSfeJJKRO9JFRI8bRbv1WtTP5w8Anj1nS4kFXsAIYKqrb8I0vMGGwN34t2D6sI
e2gXI58051gUkBGQbth9WmJp18m09MIKaGxkLpWv2kuZQzLBqnRnDDisontH/i3McRlzl5DfQLi1
pqIYQ6naX1nw7RpGIw4yPZyt6mgy6QXB7x7jgfdbSdaQSUCUuaYItfGFYxPum+Af3V/DUyWI8CUE
saG2TkfE4NPLBxlTeisjAXHJwtWKpEVFpk5e5pXtITJ5Yglh68qmzXgErozTag2HjctBv4BIdEJL
egl4jiVF/NftuVvG2a0xsdaOqxceJ8sJdo8s9dxGalRSLqc3Ev/tfMwKyuFqARHCj7baF6SALhUa
ZW2d0bkZF3u9+DUmvUjIZrVpMIPRzIQJzv9K7ytFhXOSXnLGOrzqDhyVzq7zlzADFBb+GiUu3pMs
CddFsHtFhpVuiZx7ycznkzsJ6gUfG1j1NYKVE8ib7HpCuj8qKPfNUPrVWDpK9xxRcS9t+LLwb+Bf
hmKzIgz55bPssYBMIKiIVzTWCNxVFCu8WiRWD3GiwkV2ZJQ8HeI0vHlMuo9hnSFTsPU1jjkenbHg
ZP+aQKVdDhSuTaarOwdrNBB2S5RtZMSw7/cvJGAaidcNYxKjbSMDKHmzq1IsnJoPv+zwTlb7Qhb/
i7WjP809fqqWKSC2pdnE9I/6/F6PYKWGFzk4yeaHJKPbFEsFkTT2B8K2/+Z3vOsfwTA61A5tjN6f
qQidWI7lf7GZWqPu8msxylmTLjeJNl4oU7qEuskB3NyWgV4x23qYk6Ax+V/HclBg+DsSicKB8exD
cN1Y8QENohEUGpLfQJ1lNA5xAKZ68Nflx1VK2z3FifRAv0HDXHeFzC7p+LEWETlA8o+qoBnEw92i
nIaTSbnoceQqND/aQidxgMiQhe4fd649XOBk+5ijXPXKSoLF/sekotib4aeSTD4ZlNZ2MeYJ9rpC
RvksVfSW2WMuJuU8LAxQBT2/4XPHOU8I1xkawUGme8klemF6k6/oiyx2y/4uL4YPoiFq1d6SJtnZ
qaFd3V/5mAqRUx31Rodlb8LqVLTw5EzF4LDNVqIeOOuhpHv8OM8jcwfBxNGRZXjQHxvjJNdl8CCC
XAZg02QFW4TvUujF81bDiKQsDJsC4BIh6VJeeym/U8bQgqwO0Of1Ut7zlwy2zhQFTSo3gZuCl77Y
i0zB3xS03DuPeSqx0DiQ+mY7uSFD1rXzU82NlVX7VhwYYH0qnCF1Mi+1vDYdCRjn0vR1nzHhmjV9
ytQlQRYHZCqAxbU9x+PO6Lbv3MAAb6U2CT9g24AbWnNJnDoxnCGN7nQtSM428RYlcoR0uouFsmNY
1NN6Fd17qR1/wU1kiDu9lKtOTop45zaPruAKGsaFHKyjTHAxrNZSKzIWbhq3OAFMyosl+xjkzs/G
K9V4BkpbTYWszHujGKAyOCdQ4VPdeiBV4XW4LSs+yWXsVETnuyP0KcMtP4c00Kc4ysJm6rNBtbXx
RXOwQN1SDcXR15GB7nVZpuiROQUSqEOzQSF2U8AYi7jCUTeZD5YBjbKwYOv7PDZOAsKwOpojOT/N
BtzBqUfQcJ1xASj4qgGTrbeqv6pnLcJTwh2vT3TUDyzGCTabb1jHn4Vt9s6EnGNL0vmSjq0mSY3W
9+urD8rppnRz1tChXvuYsPoZiS6DMTe3zJQ/y+HFGCmSdDD6+UbEtg2t54A/sy1aTyFoySak1miP
TmEGVuEWoC6G48xjK6j8TevVcBCAsWRYZzHxTXDt+A0YUIclud7cAJo6poCRKZCs7kNABFCibSEu
S20Mpy/QxeWT69TI94/mi/lmGSla44Mnk1W3cU2Mw1lkwYNmwgaP+UqhiG5+Bg2I5zWwvUQqQ5wb
RrJ7Lf+NVjwLhtHb44s6Doif0rZz/7FVfOjqbPapc6jhLPwI4zCH30nykPocbgaH2BMSmn6aQDVH
xQI1XwdZA+okVxPUM6cxg4GJJic8fthXefTKHFa/GyYEMeBck9tuCbNjRfe1Hs18ZwCgjBB3/HbX
WHVMEUJ5ec6D9kX9BSKMZWFsat8UdGq0K3YREEglHotIlxDJX+IfJKT9uNrlEvEirWOjwtT75sLf
i8MkY8jNJ797OoWiGoHgjLgaMKsqaETVgvnAEhL1L8STJ60I6RUaBV1YxiCw3pOObhwS89nQMb8Y
f4BaDCu4X695KEMtCipT5pWeFDX/7YGNAwBl7mcIFKbcHg1yFG6ZfmdwTfaEHNFZ0R5Ho3mhh7Ks
djAStNH4KYryaWSFcCnImsWyksTEGYQEwGoThaFOOgETouz3ON2p+eY5FQNGC4+lQLNG1silmymG
YEcUWGAiaJmVBL4UMpmacestPCRO8NSS0vhJkx3YmvBHMfKWAtK6HgSO6KoNdqJZICMMU7jv/Si0
u19R0onJjjl5I0vCq6fqYzxftgpL2xsn2WZQfDCHf44bRCtbsmms3Qzk11Ey9jaM5zTrx/kNdyKr
bR0zhO0JtZwhgBDeMVGJzCdWQionC+XdvdtO1rtb2VA75g5Jw0x0fnPKwrbArDJjXf7DffWGdrP1
+1Az7Nmi7bwZBmiB5oJgNV91pmz+a2mRyKdYi9uWXkNvTgiH/16qIy/JBxs9Noj2J5/HIDI+UUzM
C7nFwEmEJewicC16Js2vA7kOvSjJTEC/U+7mtQU1+c/MN/ykzU0Z9DnRCxTjbaYdu2KNlAbDjWTj
C0LmrLsq4nIo/4dLPr+EVsf319LS4MZp40Yb+X4qIo6U/Z3DRBsOkmqYYJWYQpyj09fJSwNJFNbf
8dP9LmMibyU8goHctv4QXAI8uIf3JRr7Ub2RoD/phDR6auU94HL4FzxfYlBQj7Ytr0/637wA6jx0
yoI3jlTyq1wB16Mj46QzDrLojajkpEfJ/ss2kTX4vs32dRQj0/GGIsKUzFtpCo/MaAb0NDC47pRG
MlM2QxBtlk2AapndLdy4Aq1SSJDGoiC9vy4GGSgi7LRoD0H9C4KU5+FownsztjF6KWqgMog1sTHe
t+w5OR9YbfZ/VBxmMe3X7xJ2Uq5JgX4Dq/hBWvN1npeHLraDfj678h5K2jkpotp6x4Lo5ONlTsw4
EJZmnh4wa1dH+mSioAxoFzu4lMmY4QX92odbi1TfGnFi4cHhA/JrY5GRVBkBgM/Ljlv0LRHZ/X3+
KjGeWT8d9Dd1XCUItb1+RkgkYLGOxe3D2YGHelk80X8MEUccT156dAdLmomDqz9I5oqfX/sSGDKj
yW4hOwmTvFWFky5eFHbXG1BQR8SLrTi+tcAZ41w4Aywc41LiHACLYgHFVHV7JHW8IZITXPBan0Ep
6n4jNqmx4I8BZ0TMVirQFs3sBq2QMHb24uUODIOlsfCOBMhYtm6o7ipMiHh/AJNSjObxVKL3AVy+
Gx7TZYDXnHzuHjXwXyq/ZpFZ+LhunbEnzUtX5xiJ7vkf+zGvBEc8S4w3XIWp5paqlgAObbCwNKDT
mtA2xK2rjSf2jJ1laFpfSK6RUia04JqxDcsAlU6gQVAlpnYpAHxxXZsrF60oCpxFMsrdYhUdsbKv
1l4TgFKz+NT1QpGRg162Y7g10aPoiDeyEPkU5L6BoAYZ9FKL5VX/NZNYz/8qTOb/ZVxn9BswwDcz
PdrGY6idpmNrHCkxk1OxPS5mxZyd45+yJuyLpQPzshMOKoT0brfZLBZupDs0swlcSOKgc2EMdsJs
gFlTJXBq0nVUIc0TTmuA4mj3k/TfG11Hd5uJpVbkaHrMp3l1QRXU0D8a07qylnrDUUi9x/A4b5vz
V3xsMDZVNimWGAAfVKuefxoA19GYq2z9+HR9TVeQr8fAVr/omQISnjYGQMR96Cgiay2Plh0vu+tG
1CBsWug/BmjwraMx9MJ9aeBNFwusfSLXfkl82JgDmAaJG60wJK1IWoKhF8G78g/dAqvfDk+qxGt6
UeXpxnCc967mdRFrPixf6bWZ3gJOXODOLevXuAgp414KnRNT+5rausiT9Fz1P9FoEmAidiVr1/92
EVSNVRw5dIJ4jX7FajoNQp7d3qIevPrgTToTnyBNefiqfnfUrJCpeUkIUvJ1Uvi3uiqkgeK/PmHq
qxeE8R+l3TXN1u3gz72MSwLJJ7KV6/GbIhRCHCYJ49htuFrCO/crQGV3N7a18wbFv2AtiGF3TJed
MtRqY8Qyt8h/6PFgQQ239+Mw2g1o/yLT6WHAlBES6wDO3Y5jeI6LPJg6jks1pHu4k9KoisnFtoS3
um4cO/2ORiXVE+8pSsRKysulI3t6CkfGKN9ZwKvHH1/nMteNxdPsG2rwl7EzMjud+5fx5n2eqOJU
qRlYTOb7jcGEs3zXAy1OPlEsNxEkzzIM9QMX61YQXuY3Crfu/g7M1pGar4+mwkIzVKsB4yJrFIEU
M5fMXlEWOWpXhKqkwnQo23+idkqhXyVwOyXmfk3RJ8JP4h/5R1j951Bqvrx9Fzrj0r+lnWRgWml4
/6uV/rBBJpRyqjGs7hlMSVE8WoKdY+mA9CiqlQmP7vt/4kDwfEF+WQA1oaiyU90Lb1cJFeXruAqQ
wJyKCaiaDNF9wdZNnrrdcDRTNcmHocxx0U9yBjVWHRu0yudEnc6+FrVZCaLmjtICeoZUSmzyhL3f
vN3Jo/GeHn6qM2Rf82J9HEjNAPJEQPDC4WshyyPzf9cv4Hs4LxhugvRfucMlMYNxEMimO0WhzFI1
DwXAlETBrP98p73kw02uJdToc1ucvo4f31di5QyyHNcbFkMzgN9l7KI0jxoIqqcFL+RfDU/htQQd
wSsz7o9QMZxk9S2kXiv6FCmTf4ydfCW5+bEMcQwGzt5aNK+zZPrU6d7n0nNEcs3VWBFKPnRb2hZk
YkSM9s2yMy4LMeszs81LRNyNzXqbauF3VvBNDf/wzteZWYdlHUq8z2Vz2jhQnVtJmhgZ8h7dZhPn
zHUyGTGaiD24igYj4D/mUEJJFv8B3G7azh0SXrVqdOHqj7cDmU5H0mGJtp8pqmmuuzW29WYbK6EU
KzHoOvDf6H+vGcAbah9lN7AFcss5uUUW3sSI73dFLhqiFN6Ef8hjhEjsL027LBBNrq+hJsIIXs3k
YCX7HbsdeA5Zzz9DazEeJPRtyqiiREcau5yqLBToudBYsu7QcTjR01Jy97JPbr4cSnfWFpJLsBlb
dX3RBUUm8zgLsaX098y3ad1vd7MF+zrxeUPzfuTc1kuvhsuI0gieuwbt5BzK0lbA4t6GY2VvH0KL
Z8MQX4O31t/pbbDZw/M6n+1iM2G2nY6ztOfDQSvCqxPRJwtNUFImgYmoYQXXvqnLGOT5FIJ35ARE
1XVN6K4RoORd9xC1eNf7vCMBeGFWYLWZMvah9Y9OSkwXffYl0ct5FEsnTrb5mUqifhdfT19w+XiM
Sfp/kjjSaM9G+BLM0nXWa43hpUVBXwYBoov90ijpKFoVcTU0pxoe+fcwTLcOz/MaDzb7UnrPbjl1
mncXdrQ0Uab1wjtYfsc30kRgqV7klAG9E6gXwJh/ih92VHqj1Y6wu7/lodiBBy+pyBaxDFGxqpPJ
TJWwsQ1ZcMxq9V1qufDMFlOkYwdbs7YOy1lhIXIJ4VYH21qvNFGrNZjT3XyFU3OkoTnLpUCSemhh
oPnRmNynvBJp/pVxS8zFTPMSjcra/CZIIEwdOPAUfWk6H1Lr95tvEDj38t57/vmzfWez0PqlotBC
MhVGHj0iRDQ9PbTOEZGQwKr4+QMEK8LnfdBW456e4DMwZpbdjzd1VRFWXjBXB2u0Pr1pB8Pr/t6A
yaC3ujdKWNvd4r4rBEdfKAY+c9llg/BgcZrsgupHoXtj7fVeedF/9ibmYu45Uv8fSbYp2zz7CHDt
5cs3tAJMgraPJkBPYmpH2ItxbZFnThekYf/qBGbHPpNcNkjrYRpR2qUdUy0FsNovOrSyRxMm3Cfr
KRhQeVU31Gl7IbtIGhYo2BIfjs/ZbMFGZQjCzYcViCA+Mh/lEV0oFOzSQxT50GlM0rK6mVCc/wEv
+zrC8Gugq1ErO6LMAq2+MEX2TvJ0jJCr7tboo81EnA/sWTv+TPvWWcJYA23ZsHhTy6qsODKrA+vJ
uNqPC+4NDBTM3ykRGm+iAYB+71GPy/f8Oop8yCclqNL8cus0pqSyBryYJqVxg84CbVe9xPbLJkS/
hZJpb5M29rQgjtZB0VMvTE9ZH4cr3ApnI1bwHRuo16nBuY1zoJylwgOjptT+0CjYM1/+iVRyggnL
jhIAmjyFoeZNt4zPsFb+OW1G1uZWX6DDjkK72ilhaRiUy9QWmvcrt5hGnJdvc5TBExsGP6qMqDm3
qCawhq/iadDxlbtu59AYGPiq8kcfdpRraSKnsaMAFPw+Okc2E3zqG1xIE1q7wFu8uOQchaYYxVwM
+2Sp4oeQ7D0rsARJI6oTOuxkEHQL5v5QM12ogvYGLAWVKv1sf3Ks9xD2VNPKmiLxyG0BZPE6VmLu
pTjishJNOiIPNmevM+6GoGJQD03Sk4yIqyBTbld+4nJo/46dPORU+kQIek+1M0Ta8B0Nn/mOVTm4
efzy44RGC22xrt7AUaA9vcNZ1hATEyp+DEqf0pTwa98oD3/mDdMToHz1zPW2QQ31oKqyyLYQ9x6L
RZ9A3WHANDKt+8VLCgsG4woUaaTkPWW2IHoeA7SGpoc9tCcXL4R1XABXhhYFtoogJob/lc/6+DeE
NEG5kTikey4slHtqKxaGLvPx/lNasnOheuas1WGovihHyC/ZnikxhZSpNb3bT3rl2lxMXMfflx3q
OFn1Dj9GMeRO/MGNa/bMYOuZv6gQhoZJFFT9mDVGi+xyHr5mrIKp+C0lXB2wnMXJ4cq7K5Xq0Obu
ZcHnX0wT5xciDuMP5f7EEFq4rs7Rf3qeMo5XjVO6C16SWUiNciZZ723LXYUqBns2t85lFsDnuhYm
YczWom9WAc7yRz3Oxc1bzYK0590GPe5EN1GZqF3ZFrtKD0EbBw7lEOOwG124/1B2dJUpONExq83q
t33OKBLFGPsKoPlosaLsba3slOUtuPXfJVuomsT3zeHq291ygdDgBPoiA2fX4jH83yozhgQ2p+9R
5pmAUrtks/3gHexrxhxfmBhvPyqAxEzDXUOTPOgI3+2B6wzUwgAjQfKL7JaaRMJ3wx9iF8mEEnX5
yoMJg6o/nPdvRJGpJJt3BjIuT3GZNvsU10Ed5CyDQMgHhmnGh6SKK+gYvPJL8JglXbKqizfcZjdC
oLDXbbNONaKvJO36GXrHouEvWJaVqd96RMvCXx4hcPnVzNaMz7tXT+KLTvYpgMhbcF56VSx7jXyj
M0/fbkSwanZZVUxS5WtMf6jFA639rwph69kbK4Rqun/4++G+UkwuBk1DZp/jJMlQUmN8TFMkg+zC
WDZ4Tq2M+SYikDJgHtoZzNxKx41Mp2Q6A2RZu8YmT40FzFWUvjrUTfHS/jUGgg5jYc48ZJMpKyHx
bmEkkOqjVzWaF6rQnlroXZBubrTzBz2xfMtu07gTMrCj6vzEtnjYjf5GPJR0L1117lAMGe7FXoGa
VP/mUnYPffaMV4sG3XDDulAY885123SXvun/08/gh92eL017d1uKEU9bfGMhmIJT0t1eJ5ChDKe+
8yJMc8hG2hC0hzomZgi2ILwAn/coYshvQGdLZW/LCC5Ae7Y1xFWSl/Y1ubstHXj51/Ecbx4nFvRj
lyZkn42yBEHKpgTw5iDVhWvh6jwEkSuYtHAedMy9SeeScBPrmGyjfJuKwWOTYn07iHy+0aQ0QTrw
C5ZKpOlqNer2Va/IucSnuDNcEUnt1g3Z7zWIqH6h2ni32M27QAM8B0wPTpNt9vtYaAVa/sgS8Ozc
aB5cqcZ/wBL/YLcb+jjwvFqx5SgJeevsB9Hf32jeTvs+U76SLwKVUker8g2PRrEbYoeOc2euJCde
r03zz97cLlx+k7j1GAP1OpGT0HxvlYYt10581OmnB+vRghhl0/8HC02v3z7JCMikag2VYn/oCZxi
Ny5X0WCHMbbPNmdBuhRFPeXuo0doBFbgJC+TrnDFf/RarmW6pnGWd81Dk2tBShWhXFZyofHbcr2U
Uh7jvtJzsmr0ANYS1B1A1jC9UuDqgEDnrVPEM8jPyHVqvPPPZOTT+gmPAjZdeoZrNkEuBSqza9i0
PZZWmyWVsL5watoJQnhi0/mh1Jl7wKKAIUgn9cdreQb8tCSXks/MQvoni/QIn0mHrGyqxoDXo8IR
5/hgpJEwc0mjnBH2Z45atT0hvDQfe6QTw9xYc75LRtVnV3SkP6oq8cDOS/BFINcUkU0T4TZXslTl
ebO6eYaCTfUFnfr8XGjzuBaa/NjcY749GLE+Zl71EMeFB/E4dKyRDX7tYeh7U3dROQdnTd7jN627
Eu7orwUS5xiOAfGG2Tci0Lq8Ec7e5WIZ9nPVZqYqaZiIimosKNxLcou4ZColceRcWifXd7ktpqRj
TdsG32StAAlP8lq4eBLsfYKHPdkVp0YSA3ZPKYP18aIMeH82RBXEHgin7pZPwI07bykJoLXhYVjT
AtLO0bqnASGob/9uKY6HIoz+LB8aWC5Q6gJxcBuTxlOOyVnOFl5pABrC0NlooLD9tZt6qj5jJG6M
4Q36xWcIWRgxSdHK76cWvK97NGQj51p6GxXg2yj7X7yP0xGxbLW+NWdZiBtBqxJEasNJLduhwdCr
KBFUduZRgcRnfi/6S2hmiGUiZF2GLmlJUmxZPGpqKOzfSAUVmZ8RdKITYAaHm9qdUMCurXPNPebk
h9UlRcctNGpHEgjKFmrdowt+zRKXuXxnOkymH5YzrVokLxjLfBwHGbiEGk515nNt+GsYQpQTQlVR
sPN0QbiFHBZ6U2fyVzop+0iJQoDkwKtqN44M9pRb5q+z1A9f0u5Hs26OkHPdofefxjW0Ogi+ThWT
e++cC1DSLvLXpq1EX9ZarAPEbD4X3he7Pp/8/30ziOJzi12UqQDIobQb/OSikVjG0C/9QWDaw43g
/Lji2+/2V5CzzVj/R2K2XQWQAo2dlpwOOq4+UASn/quxiPdStJC7QTjCigG9ZWa+6E0t+/fsHqGN
PBT3BjK/fXQOOr7sejfrJK+wS9I1MiMvOU88Q/0007dECq0BmE+8CcySzDj9Zi6xwYV+5TZJ3HGO
fn9Ln/9tFsDa7IGW21WZneNIdzqL+MIRx4AO85txOtMnwtFlsZHDoqqyYAUx/YQTU/XR0EvKVxDC
Srcyatkbmo0okYzeRcbezt6XkM3ei5CU1Q0q1vxPizhrIVsG1hPgNuLix6AJ9dzs0eawFBhW8E29
K94bNeu8Cvfjt6Y0XZrpPkeSTC1CGdCpQJsntoPFzVvkGGH7SfmcPiexr/AoVxJMuu2ey9gij+8R
zRSDoqYrNKBnmN7+E44AaI6Htg+sgtExqtjCL2p0y1SRp5UqO5KAA8FwXMSpIp0dKUTgBwqEBSEq
Rt8CbGlfIjmO3br8lMOsrMjo6CYuOAAKsq509qmsGKaLqmJ0m9KHdXNaeNuLWyYqhJ1Yqy4YwNpg
jkh1queJNzER6f6UqqOIHdnlw0cQMjLKoTw0Wv1WabV6Nm/JUO9rRkAylucr0wc9Av4UBT9QE5Ie
cSo9gYqAaCZYHioMkwvqVrWoUOflydTs4vkN2hN+wCx9F/MWZIdu7DWKc+Y3cTnkrCNIHq4sEKFh
C6nPuyWjrsghFLS4R9SmVF3/Ad0szu0fNdsL95V6tF3rhzno/0Ac3dQOD/ALg5k6X64jDM1h+ppU
KnBUO1Z+rpZuZRSK8TgRMy0VpiXJqYldD23+wHzLiyJuIoQ4dxT/L9smg/IeoZaOyCCdKchp0a60
+jyqWl7IE4JSEQZF2hP65cZpnDoe7wRTyC9uFSqkMkAtJ1gnpfJ72o6gIL/8IVfjNybGLsl7ZWlz
QxEwNjwzHZM/SVRyupy5MZLXx4QDQdd3doGEtsTXR5SxEWodvN3VAaX1mK1h8iaiQuce+OhTAi8v
L4uBHXGi2IbPCawoiaKh67s+NFPKJ4uL3JwQJat32hRMz3nx7xZ5uEv9J8uJRHL8dJj5/Efiu1GZ
CevYxnm2IPMdpmyrsLDfj1Qddc8L+hGu6RfyPG53c/1cnQwoRZcVoqJmr6TX94XzATu6AmuJHvTR
z1OyDvHOQ59tax069B164+TGaEynWqPex+XtMgvcKMSR8Ntw8M7iDmk+oIo5CWSKBlCOe101fYCd
ViOJ/+B9XY5Oa9qnZZeg2MB8Ta/PIMmiefm+QVzNqaD4/fXFjavSJPA3G+hqb75kR2WqiFrnF7B/
wH6s7an96yhNAXk6J5oPHJj5sbpFnGBvEB1ZyI2Te1UlWG8ZZogsqdc9y3drmC9UjSJA65Tyh7fB
s9FDWto24SJL/FFWCbwmrbeJaqtmRA3CEN20HnoVWSXrwkM4WkudrawCYdKea0Av+DWFUCgPVjqq
hzRLx+xvpRCfxN4zYxQsKzBjpG2FbMlQ67LhQGVcCgh8eTpHEmHJ37yjk8Pq+cjz56tMhGEMNI1M
6qFEbp7L09nwhYr9k3YGPXr61M6vLBj+U3UhJFFFgnCKiKR4FiQqjLRUdmLg+S2GaHEuAMFbAN+F
zFD0ePA/XIy8H/c0pUjbWeZP+8kEQ3qhbSNQrap1+BJ8KQJib13+vlHq0ac5kWE1qFmr7F5X/6VY
qsKV7+j03KvYcerYUjJZR7ggXf1/de1eTGQmGcy+Tjs3Bcx1LcRGqraBFe7hvdlJguWLDBlT9SnJ
WOHiG303UF9VDkeJy7cjsjFppn3sJsFnVS3Qd9I/EuZoEDoaSTeoI0RTPeD+n2rG5y3p0j8E2JSf
D2K45/gjb/5hAE9yTaB4vH71fPmUNzzrtEpPY2F8bPR6DOFisdCI8z31ucdfoeRZ6H0rKKZlo7LR
UPAOtqoizm/Kucvfb9XeLCPjLQNXXHoZ6Iz5yZvnppp3yvMzZkqa78s5mTCYF1GFVhOL6UTGcB6M
1v7yenuQOT84pAB3jAcOMtgOP87lVxPsTw/gncHPQoKm8Xg/o8mlwKSTBTswSe9vGE6aKmB1ZW2k
vWz9c/nMGKpycBdI7+2rVfoNEQRCrptKAQrJsDuNItxtnuVJAIZgDlFA8nfhA3VjLXSe7cQb9EhX
griv3rzaCvnxHlJaUu6dCHVhh662ReCJeu8OkQVKNNqejlFYoBemcsPqKJTppN8V+MeTa+c9CBol
CgiYanaoEUYJiNEk96WxMYa0YOTwXz+yIhPyqRY8KEfD61Ki8RrvsqhBFkBDykM3U2SW7I8tZWto
1rD38XbaTJ2QDViXSDaEEUBVcSnUxuXQOpjK8++9b2RecqRPnuoXPn84OWo2XU6seMOJO22v18vy
/JBiuoYewq/Qn9WwsmO7H+nIRo+PDd/U2PKQ2Jdo7wL8nMmmcEaOVZZJ+sJo2wFAX6aPSWEVeiyd
1GuqlkdJ/WiEePG2cACfsYuM0Q31TO65qiNjT2pDtec3hw6+wp1W/9jDCWPVsyOsriGUTwnxedz9
pQOeEBxrOZjvIdX+8C1hvPrJnHLl/ZKK8K/PunwF0hz+F2w+Up1PfLlMaPjwyzSaf21Xe+hRt9Zf
ss70JrqBuXG+gHppA/3TNdt0L3fWUlj0PI8OxXzoQ+xXEAHE1lEfl1Ds0iOPEWC68wmM34zfvBc+
GivTRfYXO0yRa9T5/Ucet9lNezUhdHeNSkqNKdOldqHuzxiriX49FKKJAViUlDraO2pD3LwYTofl
18YqNEGUlSCRsfYJ7GJfPCCSX7s3s4vk7V57HlQUG9u7Ct1zEY+mlB5GTY+6OLedHyfA/oqYTSnQ
h2N6YwoMQM6odggbWMVwuKnRse99sMbJREpYr5xqB1N1niMlcpIef+MFYKIrMeSHCCHcWmFdAxf5
2euBF8Cqa8pmoQ2Hmha7SFIP4geuZKdc7g6mAD7XX1hpvyuLL2+BOlKBK6idtjZtR93GSVj5wnDF
i0tbBsiEvu2zzX5GxcUG2f9xPql0W7c7ABb6eC3VmLaXOYA9jL78OceRJ0ZjO5/lXaVqZL26AjzS
g2gtyY9KEhKdjetN6rquMTBaGjMkhneqkM12FwMxqwyeGCIU1kSK0fzFCqeiewEc/avEe/km3i2k
tmjJpmJVQDzpd/JjlLeYaaPlcgxZIVwRwhAF4wR9Mn/lPrNSFfTohLIUHCKbJN86jzUpBCuQ6tmU
V2ysSbbHXyLxhO/DIpC5tdHYrMZ46qK6sPQ6fVSyP5HSNCsOjPOrqeYtGjGFqoQKFDyw8JnW7UMI
IJuIxw214y1ACDKIxTKYbh8TsVHYtMWWmtBqd/PsBARrGR51nxVJ1ppsBEvEQEKtScgvkeqGquTY
AfTBUUU8mWNRHfm9kJHPo2DWJxtrU3X0E+J8+PmwsTHVRQqKVUtb0Bhv4Vl5BIFCZiWOeUrnNTQe
5UuRj3Gq2QAVwt8/RuKSw/f/IwtCcfRWZfgfnWVsZS87ywiZ/qPaNLflNeFfAjw67ASGykkWhehg
a8mhGxKWWQc16o3+tP+x6ClRURfudK7evsFR3NmtSKAHzGT2TApqWyc2lgsQoqCJYYLO9Yb8g6TI
aQJIQUTLsxBoP5iRGh88FQM9+n8RR+UVfU1jlp+QZ6AuBQmkw4/VousETVfuPC5zxP0GdhTLtAW0
kT8ZIaKlwDyfrRXJpcZDgVQSQtKqMawJ39xtTto8u+rQe7x46GT2XjxW5x5M+WfZeGysuX4jbVDu
ZfJlK1xBJPJLrChu7Gv9fd8o3vRcp5VLyXzbeuB6EN3gDulGZ0dKb8ZpMrmncBIAnUlksY7rkAyS
Xf0usnAQ/lM1YjWITHI+SxtmoGcL+WxvYGuUfGZ4SAEkS4dDeq7HEWUdA7XUMcsoVrpKsgmTlUjR
w8peAhQfe644MsWuY0UZGWO8z9hFKr58spT+rTNxX1uDs6siVAn/AUeGgcaBy9sSOzIZIa7BruYY
gqkudVvtSJu+2FUtB//Pu6DDtcT6MfFJ/tRjfVuQLvImvIyc23YLMm4hJzck01NE/9o0y/ezbbLW
HlAiEpZRi02dA2pA/WH6BpLTxCi3p5ZyiSVhrSXgV5hCBc9naInHN9IOI5/0jckYdG+yO/kmAiP4
8qvVezxQxZ9NwlVx04kMSiZzeO0cqh2mNCcMCK1Up//QPjhy65H+Dvcj95BpyvGMQIhfMFfy8bzL
b4p87xlEWKKpGdl2pwQ0czuMgtT1b7Ae8xdPxcRC2pHQ82r8rpbfv/JvQU3iV6Bu8eBcEvzIeReL
xl33PmwSbITk9WpCyqe9YUxThHzD1DdavYa1yiJRTfdRwDcFpFuhULWpy+x/0U+PnfnRyJL6WMpR
7x3Gy/oPpD5qQf+zL2Hapr9dUfZ7T31uS0oJCM5WG4Xuqo2I6A29WsitwpcJh0rxl9/bPHZmyERv
AxaeVh/vSAHYlLZEEYTzBNVXzq+fN6FuS8ZBIXDdSkHPbOGrmz5buB43gz/vFVqlGZfV27tuqW1Y
TiHa5cShK+i1+lxaG5XfkOqE41/fmaYbuAO5FKYgNjRsKxfn4aUW6QiBHafJJ/FpvbRPBBablgoN
Y9g/OZ3QPskNmkIIOIlfQFxqJUHEotEj0IB3zzTLpLqe1L/Gxn3wXSXHn0oQWtwwFiyNdJLB6NO+
R+58JyNgqbk1oltWH6v6z1Jq0vEMgpolQ+RoKHtmuT/3VZqaDIBPdeS56GTwbk7l0FByix/EQcAn
I2PNkFBMEOrZNXw4V2rGOO+NzjLrvqcdNpowKfM8jgHHAKdmhnSI1oILE/r6vNiCZNObGKQIROtY
aZ3o5yhYujcP7xpFUlE/TvAR7sq85/k2KmiUvZrkFcvHLRyzs4pscv5aD2kc1uAr44hlpbYTBf7z
Mcs276/wcpTMTypVTUsuQ3BLUNBXA5wIT+8b2zn6KyVlB5mt1hJspahHdEmdU2hhsBLx4IblUBoz
TrmVxUlZW6qy51tP95z32bCbXsaBYlwWDy7P1xnUoPb+KlaWQA9KPkHhS42U9nwmtpXpOAXW6bhQ
UK7xSdtG/tNRgf9OxHjaFYRV6LpKH2KoZOw8+0XS/qKDMaCTu7fJ+/KkUnQzaP88GwZ+n3LYT0QV
JrxW3GaBxj7EM/CcB+lVwBeyWYkrZRxi2Xd9Y+T0asmtvNM8mNDTFWElecQYGagqewaKfWT/iJld
Z3BuHLmqrPa8T8vlm8Qq+MrG8/zSCJjV15Gh3NrVvnYP8v5eIWPZ4xJKoPEy+7RfCuKIopZADEKX
LGuH4I1hTCVDU1J6si2ycWmkyMTTe6EQztA9Y4NGQ2EVII0pzQzE7Pn+JIn7DI4C1+yQjcDw3aLJ
XGqudsOi4PeeauZpwiC7dGPs/DvLIn0PNDfGq50qjTUFp2p+NoQLVYqmCOxrh3nyAe7TJvOXWEol
OuUGXwj3glpjs9AUjrRUgWFJsx8yUIKu8GMky9884DYg3upZpbCPjQOcgWFi9kBS9yBQDdvEC8DE
7+f0349hRqduzLLLsjFijgzfdoGkl1JHwIn18xwqsedM90fjvSwZE0xIqrBtORXu7jPLPRi+iNps
UnejuNgGsICCViQfeck2+zuG7lRH9C3ux+yJrvN2p6Ryw+JqPNRQGlM57B+UElrKnhJOzja8O8yF
meHe+gpiDleBLB28Sc15C7EUDreYUAQQ6+4SNHjMlp5Cfl/BaiHUw+d8Quvh4C0uIa8MF9faRLxm
i2SaXvONZshlPSJWBqx/9M7n8ih4jHCcBxEe0llKNl9uhoNVScjg1RmVVvUjA2DVkG/7TUMbk8XQ
X5GW/ZubKmuilF2AFC9L6fcWI+QctRBlg+9LeDnFBu/StkQNtB7JzSIdaR2+DpG+g7QfhAiJsO6F
hqHAnAtcyasv+bFHV8l2y1zaGnSRxgLzwls273D8EzbSi4SeOkwWluxaZln2KzxIrFpsSxYFHzcL
ISfYY0zgXd3M8pakGxrp2xnj+bgc7R1WaCffoa9hi7lOD+CdV3ipQIy7j5gNZCZ9dQqkRetNYNK1
Ucq4XUaKwl/JVIrZ623m6HAUTikEFs5K+qX8lg8on7zv2VV/w8j+mloZSQWzTl9yXQ6A4KeVeNF7
hWU6ikAS92sMC7MS210zVM/V+qkxths5BOgLw65B0OvH9k4uXxCdU+toe3wi4z2ooyFMISaFHMo6
+cGkcJ9/Lt+sR4X+6urZwHfYzReFsAxFDBguMmdZMy6F5ktvOpQyMpcC7MVzITOsTF4jVsneF4cZ
Nlb7yXhkNcPsS6riBl4ca85ws2FMatJLM/A8ZI9OqyzPcjzqKK3DkFfBQ6rhPWqKNxNj0Kj2MqT7
zThRZiJZWNjRFyUQEIjqrXObXVKn62oKRE/f4ixfOpK9sl8EZkCjzAEnwle5kGu998jtKKkaYXeW
MOlZXtVLxj8sufAhUabC/eOvDZ0u8xqekNt9zUnje0vV2WhUMbvwbDHKnRwV3F3kZMRyES8IXSso
Q+8fUsB86aJYMdvgGmdITPi4liizZdiTu4N3yvSiYO8ENUPbXjFaw+mjqdygx3gHapIB6Hkz181N
wa05I/Xr6Y6Zo23gs9pDCX4DIrqwpIKybKAVzQogMJeDsQL6tL6aUoCbwSTDL0qDOGbMqR3erDxd
X8MrVx8SxTbjIlUjrUF6D/WFxLmtSMpK2KgsgO8EC9wgDUt8+Rf4rGqbbFNz4/CRMXjrtN9xBCHB
qM0MNh9c5ZHCqRFuBSDSh6oZUVCmNd2GZv1PNFOE7XkslQIPClWbEAEV0oUNdByu0+LWrMKGD7s4
5uW+92hrzThxE9PUphs3pHCaDd5zS/l95Yn7JiphvvwYNmr0p95CKLtXk36DKItgk6Ch0qBDA76S
ku6lMAfijbOEPKyWQcZINMluER6PStr94GTGIBtixPr94HV1AxPKpKLmVtiiArAgk5QG04KW/5rQ
+LnBhBXcCdYhoPtf7AuyrqFZ42E2Btflh/0WWKue0KHVW20sNY47491Byto8ceAU5b3YIoDyEYY7
gsaKnEFYTl5pLd9Sdz+Hytv5KKypluUdXMvrshsb0ah9AdPEiWo0zyC7axcIPMY3NykbebE8ol0c
PsD7ltHETyii7ZgRQp4ytpwD0lQt09sIH1/7+sNOgOgO11IJ+k2otPf6gamzR19c+WZhYRQV3C/A
3jkvHrBDZxu2chqqIG0CZoI3VMxOsgpx2IDm3STvSqIDpRrFM0JV2uFQ86/JwJHkaaEpPfDjUQC5
lewgjXPCQV2atcsB67klg/43z0xyKg/69LBYcbmcdHDEw6u2yidmqR5BJxoEvq4CaNBFfNCC8fWc
ulffkU7oEXdLWnUBN+Mq+mK+TdJko+Q8kJs9uf61CebebJBUJjgMDYsMouPIRgv7pN0dCjnjfUzq
KFlGQ0yPt9Km8tqHtr0R4Z1bLjj/efa+2HyeLgL/YK3vN2dr6C2hNGScZ7l8D+JdD852w/VV58sH
hBfsZZBRLdgNy7MhzZtFw2TFBPK1c0CIcqrifOx+IGv+SbhaWkIFP1CbNM9VRTu4sWqge6Iuj7mk
TCbkcHLsiqmrrIzD6/tmAJ1vzc31HzT95kLVAitXuRXO9Xb2PGoqs44Wa7RLOJa6JuhDNq8BDqNJ
g7hr4/4h7RIuY8SMrbLmXy5tqk37V259Dq1sV561La5V3GddGQcQPickpwtKgbLUqo18pilWDI6S
NgbxY7MPgkvRByJzvde6uNABVlfvIHJrgyS+2LV4oqvWRo5Yb8rn1k+yTfvfoxvNN1SMXPJHzZY/
NUw4Gnl6eMoetM6zYxQeJ+oWP3lHPRqirw8h4n6/sauRRn2wFQvqWvd551/FCXYJ+jiUELMj8POp
g8YoD3wjjqM52nF54qQjc+uO7QG4yMqX3ZmqS8diCpHcWhjQJ2NzYEyb8uJY0u0o+tJNkOjxay98
owOATz11wBAilrGhhWYD3FQr0ISl5kxT8J1o4aw5HCTT2UTjnWtMwws0tZuayex4HyC1W3CVs4b5
BIkTILKLLbDt5UGuZ44BaAfD3rfb8lmKs42m0wDuaZ5Pf1JO+2AiSY9QWxkHDLlocVVHfG4dk/qp
amFjFqROPFo/BEXwuMKZiDXcia7Q67Qru46zuPKSSae9BXIf7sHMbZTxDEW81CjLoPoNIQ+2rE8L
XMVLZJ9P/HiUSit6aTZ55zgFcahuo1AJtlQc56Yy2VkuPAUprYSGcB2+RpiqXSIgCQe92WARAJeE
CK+Wgfq9gkNV2SjRBE04W1EPNAehCX8n5tLZI+1wPp9WC9LMquckhg+W15lVzxGG7OTq0inmk5Wj
D+6KHbNP8ZCjpIHw7/ZRuXrI/cV0Sp2ZjYNrnkSWZTVbYXs1ZBBn+oIVs9npKTYo0FmFPAqhfvoB
eOO0KbB7Do30vKGs5HV33Jz5T6oDv4+trdUunQicYLt6eL3Y/kMcl+YxJPTbZ03ca6izLScEmpD2
5q6DYxaUZN+AQNyqj1+A3ikalGfKllUu70ntFetEAfpaCpCChh6dt9agEokRRY6URYgSIKt5J0Gy
ndj3+D7pOIIaTSbjnB0pPZfvf/85Buv4WEALrrnvTmEDXme/NUNPNhOmTkFJdmQeCO8b20wa3s5t
zivpddBE8Zq2AJU7LHWHefsUuJHxCuC7ghFVSi37AGPhu8vejqHmeCoi5Fq184gsarg3kiGaV79H
TZ2ZxBuw1nICLjBrBbxpmVf6x7ZWH5qaVTEFUOtJcU+SeunbEmTd+q1xbgAZzb8f5q34MVTuJQAN
bbX0/OECqyOsOxF5gg1gXHnzrpjwX8KRt1Nos/edHRNzfzW828V3pR/+KvIRJrOISFFFjl/jTLqR
rzSFOmsmx+m31rR1AVvS2gEdYaKdWThR7+cQh0hZckcWclIQ3koTD6kR7YMxwHCXcmAaPzuTBsjx
axjeQATqCp2NqN5Q1YXSw31xHbD5kEXapSxlZGZetiHBE7ixlHEUpzQ+wkGTVQAPsQ0DrSVY18Rs
TeBZTcAPZJh96Rr/WUmkuPOthm4c15dfilrVJmK9+iw5lMjSj1SEfezN9OFCUhFEEi7yA7C8Mesy
6sdv4aDlPhrApa6rND1Ayt5jHutypgdWYRUA8jOeZMAoi3A+7C669XDCO5Y4vsmg3U4DdVAvevT+
66FIJ82Cyo7SzwteyIKqvwMG1wt7Zw9iCutzpE5vTivdtPMN+iXJSPy68/s4Wxam66oJKeR4EG33
VT7+ISbLscwO1cCXL8tWUSPkIYoAiX4xRvB35P6WgDtebmizC1iDrLrxIKpbmD+WWigxvEZgS3f6
ph6Xy0UvYRTxOkqKZfIA8F/g9//HenmDuyRNcJw/9Kqrtf6CE0M+28veFevYIhBjO1QEoeTEbpzg
9ffZCECuyyVo6Ut7FGiec83RZ2/Xa5zSoo6I/WgkituuiPlLaioCIJyUPpwfkDx8fjQQinZlKJ3c
XCJ/0uM+JKHs/4Yq89R0/ypBRrPnE4pNPyPoN3IQYk+1KnFHvdwquTkV9lu/VCZHlepkxKQInNjQ
Ar0HEybA27UV7UdgMHdiNbT1IoV2hT162oMobzVAMnXgtuzMhZjn95+Qzzm44nCjZnWDRo/Dedc3
Lu87K96PuD2KjW2CdA9RbacQaRnk76czWOTxsETdq2oJEmNAmpYGNQTBsvESw0vg2rG6L7zYnhsh
kLSaQcJT6uXIfX0PqOkytddZfzbA7Jy7EoJcIgIInYNl7s2yw4DerAP6WreYqvk91I7W9sVsZLUJ
6hGI2BSzkVak6scPzaaVQzr+Ui6wsR1yWvVpbtYDm4pDEBVbiR3MyqK5Sd/I8P5y4qoNeItI3k4q
2OZOo5QTZdrx3gHmmw7jRN6NJvFf0pb/dhKXkcMA/vEEO/aMC6W1CIurFZrJL7+UbNGKekrjrnVp
eHLCvqgvy00XOMzJmI+4spdVDYAwAU60FMfjXf5Gd48DScQ71+Z+TMPYu0+f7zBfERcZ/Maxl97u
ZQBBcNG9TW6qbP+Q0x1n39PXdN6s7WOI1QEgv/9urN7Wdp6Yeg9kpUI3jfcVBs67OamfTF0odVxP
US54OSu55du0SUqxKe/Inq7DU6DT6OkMjapJvL0r46L4yL6u/yP4fwYUYD5mfKZhZGqxQrMDJ+9P
qcqRf7M2JmkGmZF9xkdSG68IxIZHhbBkEySCDAd7x+7y56u1rv3yGNmolRzOf5yGxhhOIkanjmVO
LQH+DRw92/5vhMFXZqfzQ4+8kX+0BkfFbOh/fYCWo0CG7j/H/Dw8fBUNsl2jjKrgcvHORHibBjjt
QqzLpJ4tNAb1Fp0YQDf6qGbulY7B3nkj4ExU7MK+ck9RnfC8JkdBdbxDvUf/qVvn0j8lGd+wgAtX
UATEvZLnnUTNaZz6ZygZTjZxDi2Vfp1Ss/r51LH+22AIiPZ0s0gLrsSxXLR7J7v1pGM8qBbvw9v1
RXozRxAZEv9rYM6ZPXIWzu7KD4TIniOKOUWABB4IbkaEOwzPCJ9jJTkBZsMg/dvhwkO/GQmZyNL0
+GreB5TsRjHO4IYQ8/qClktLgmK6d9cqBSD4NbbJWn5eHM9Uj52DNLWw7hg3JZASPhKC3KHZBoua
IALNEntWXRHdUkGIHkpfbQG4ykMSJG255146x6zH4lNMbLAuz3A2vrR3qVjUoI2ZXJfV/aWbL1pQ
jD0ZhFxKjMy/Yr0S5leftURv+zpyZMnLgRrfh3KJRu3W+4ts0koXH6EtlEBJiQ4dweGcOUL5SuXA
cglX+B5de4Xbw6deDwXTdI9MSsV0KDMutmAmbSsMIdCBVlYm3FUaBtHFQsRrYWCyvDbd8Ka3zn70
Tq1Gr3QsLomng6TdoyfFvQjgbPDWXamp7Epmuu2PWspI7vtkX3I7tgs2dFFR1vqKOz6eiLN8fPbz
0NfGElUGsBo3euiZhgj66xVG1OKOmrYtYz1jH3HuocuJRX4Y2vd1ubWYH9dfMaswQXNR1gUtFuPe
6QM8QR+/d+mtVniRKfdif0vXccgdoBvkJ5fwqlBSlBrvKpX1MTlK/Eqr9YC57fSZt3IqAiXScneV
wwfBvTmLZQASwzBsSG2FznUWoxSikcBIm/uPaAjCmwar0x9eeFbYxj2WejLnKl+vWedvd5/QRCHO
aXFM99SOOf+8pd3qKqop2RoTfQYhIZn9wQX4aDJyzxvC51hZVivwlllxt+eKUg0C1L2clWPKdZu5
ZVs7t+MLC0/JnoWT9OpJBFIemjyiPmv/cQV7qVs8aDPUm+g7KbVTbL4KXqVT5CKryKDyNhOoeHUg
WYGjon28gdlfgjPgLb2qOyxWI0Ho7QU5MYSneaMTT6qHQ/e/zfvUKzU5u+GkPwn8eFWK5czpgDXp
ItmuDXDGUT/fUZkVW6RoWUS1tUD5fblaZApGwxapkYePZTZ8yTN6nApSl3XX2QbKixlM7+8aQO6d
Wi9TuKwR9MgTc108iuxVfDCR4fnlcCmosNm/xHpk1Y1UY1NgGzpeQvsRp4Q3Hb5mt//tvG2cgL4K
i/jmsxQ6cofWFc7NeTE/LGbafXhqOsj24jFypOeLVeij6IKr/2ZdFKin4jAo9Ri/WE1UoQinx713
sRvOEaGvo07n4h73zUrTzXGn1bI2xoPMIdKLZJS/oQIU5ub97aLm9dZoq5HCbIOVfOF37VVRoXMC
gd0eig/iOtyDE7CroG1F3dTEn5QCZXVMgvOGfRPa4uBXm5YTk+3sop0g7FY8Ztw4e9b7cCPI2Lc5
GoLlu/Fld45Esab+yWTV7t27q7s4Xc4c0Y9K7kse26wBl/xKnrb12/HZrKfPexxjLP0aSj+3F4Um
jOYCpfbtwDE495M3PBrJzMnA36fOAGSGznr0szl/kFyx5ul9+afap39BCb4WvgBgKnAWc5W8hQTH
QqpH4Po6eShqACNWlcVpK5n50uM6d61lNVgdv2eqh0fw3ajVnqz/idyf1eeODXFC6WNfIdmGk+Tw
XyXMeDVYjfaNmx46cIqXXdVu7jUqZaqlFUlIhVy61/a9t76XdonBv6jhHCifAUt/6RVyhY+xVM8Y
qjUd9fK39tvHTan4F8aOEEtFgseSw6/MxJn1QtoL2eK4TeKmf8kkp+FPNVC4JZblQt0WgZ0Pni/D
SBm76QxSD2TEPH3zDuTPa2F/AehIHQdpcPj2fZ/TyvibRPqDTz1g1qYtQJnr+K+RxX0g+RCL5VmM
oCfirBHCowSF/R1S0+ajyy6nJT43mKRdrOj0EGNv3epMctrMItR0akubt+8h50ObvhNY+WujXetn
VUswkeCQ4wNLGkjvabzvNPyLBhxq7WK9NZPYzpU40zgfZ2qNODlkn+auCCjDd067lrDPQTi3Y7aQ
YzxH9+3Rk2YysoFwMlEup6VA9bnWqGE8D/LBMPBSabLl0s7f4kP2RCNwoppQ9WgRo/BWNDmBn6zm
acAsfcu5X42IF0a0sIqXb2rMYVd3GCNV3dc+6jS2WTh6P/JQ4XtEFerWGhnAjMWvHiUJZb0yCpj1
iFtyOiO23e9t0sTKFdckmA+ztm9R27RUvgIoJvkJVAoDP7dRM1S00XGRq9sZ6WjrPOayDrHAYkmZ
EDmU8mB5Qsfuyu7+MbzsnxsGKldQ/wi0bdUyDnLbpY8E2j+CMddMYNfVLzfySbzu28ZAca/rr4Vz
0Jr7JeDEXtrGJYmAO7rF5/Z+jQtifwgtYq/ZzKle7UOMdH0BSTbO40wgc1gIKY/qLnefESFRvNag
vbUkG1gfIDgzAwxw3DXkfkm9NwcyXj3JgZgITMOsrm5Nt2kL+tmQo3gSuBjyPswXTzt10ByeGbX8
8C4RS5fkKcIp0RDY5dPzjuT2AWRl2kW1sX3/HH5bkjUVFUobOc8QpLiZfzkAaHrxW/3j4ty3Lxw8
shNZqYIB7GdWdeLK1USvZ4oE4SHPjDaMHljCdFaNck/5ohFwdHMe+335/3/XkEpqlzYPw//gpcIJ
jXO51BW3oCAsmW2DIGfAMnlNHGInRYjLQfEDC1INQV+kfHXVl1mGlqylApQDxcoNGy3m/WW0U73o
IFgUpf6UjO9QULZEhKeW6N9sc8h5Mku/3DcEPVxIKWQ1jHxu8CNokW3UQPZZ2iBrezZJW8xuNIFY
8/Cm3xyz4XwkokvIAnk2HUiLhbbt9rY+a8bdDLhKJqkoRA2y7txm19FtUsGxjO9HzvXfMJILcFPv
PcsSjQxN354C8jJbEGktLyXBcpuMgJCl00JQRL03bUWjN0SdPplTVLK8KqFVqv1fH14DwE5iIN0c
2Oo204mf0y87sR1oxbHddJmq48c/JaZp6rCLOg5WJz3pS38trVbqz+g1RJioZW5VlNfy6djbAsoJ
CGaiYsP0/dzaK4ck+3FSUejX3HdMtCxmXY7ml/CZxjIn3qP2AXMaZ6dC9RM2xZsG+Ps0JugM2CZ5
VFeK8lyqcvcoQ1047CLvLcoQxEar9w/6uRIXo6wG3Ha3yz2kx3luCmWtBW3pSh9goA11Pzvvn+md
KvmaeIecFGL061lno9nSj9EgAhJH73x949Euunbo7MQMYPLbQIjUSG230kIsNSUxNSUplj6wPu/x
k1wPWNXDCI4WBkTNES9ZoFaHHv0uTQ8DLN8cfzEpeiOZlgNbaNntnQKb2pUuNoLLXZIpMZdmEzY9
0Co/5C1zy5qU27URRTdcNBodjYFJwlUU1+zW1G5/hSRKohaSV3nQDVVQ7PJw6xyWm9489Q4j/0rR
BA258sYH4cEQNZfsOPZK9cCV13HtC6ZhIg13dxjhqZXV080nMOlOf3Lk0tm45YVIzE0fcP2t8T+W
efBlecXmQp0Uf9+Ugq9fOA+F6UoZwYGQZjFyGqm648o9KJEmQETL8Toi3kMU3sTI3NSwN7sdOQen
5JYBd7DN5/0bdj379mpagRyoGZTecVtM3ecf5J5aeP6rNh5QDfyjxoegJI/wbz4PO1G6nVL02lyf
POM9JM83wVK0N/VNvu/530FIoCnQPwJodWGiEfcFhHv667QY6EsaSUUoy0gwk58B1SUO7Em6bQi+
CC9slQDDOGmIGQUShgNJYLWRwvB6Jv4TAtaW6i72M9nq5OxaNOHG2DKC43CLbTW5f5qlVXWOrw0F
x9lTgCVjulRQuXnKWeexneknxMypXN3xiSRaNvVbVUUhWJfKVgXTf65RsRgxoWpQ+PK4sa43Semd
4S/4Zno/6lv+QZHw2ZY4JCqrU40K0tqohSacbVRGYm/ZjOE4vJv6CTIPYtP4jvRzb0DgjOl07SfE
89+Zrb4y0/nT3RGPitSbEp0bh8GqqwEbTIpPwCjVjomOolt9ypREz9ZoDju5azU5FLaqHkP5gzZz
XPxxbWNQ1W+3xuIuiKAwQfqtC0NXIjCBBhNuk3CsZet3GXCSpm9Gjcu2KVdHJxoDgFmJ6iPeGH0c
UgH5TOE5K/AfFdqO51VQTWOPWQzrBBs9OjgKJSmoLDOErjsYNfNqTi7PtFNfvuOX1wURbJ/ZWEWR
/gIwHbnZb3diKhjZIfXMSTobJaUbRAh89GcMGxlLvLNpo2L7EhvanANlEDUI1IOl5T9uzl/F4HQY
E016AD4Mx8lf+otN9qxDs4O0i54kyZqU98fl87ppxytAaoUNNH267V10uA8sMThd73tK+MekIA1G
wvL/ESPnovYchjMkfwzOEdFZAbZX+eszSl9xNk5zyhWg/Ir1Cn2H4fgDMtVsDn38snNqsd/2Bbky
l4yYyF1pMDEjBrjk5jCEszlKw9raCz9WNQ6ICPI3bpJ2rJQY9eXQy2jpnTff+m9hCncP860gZEsw
re9y/WZ1ahDBHlyS4GIYbyMyC1yy12tu9zVFqcN+ERHTtljrbGK7C+h5ZkSqG82Lz7SksRMPvx4g
EKxkHwYuLzJ6DZoGLmQKfoqc80ZwNSMK9CJcj5loyyxuOvIktSl4VSyvQL8hreLYnpyD4SUYDFKj
0GeoqFEzt2JgepjHz6HcblrbV9B45eGOiEbxxi5Q/2Yw7FwqmgC2Agbni/4FwW12avnT93wxj2az
HEx/hcFNOqSHHAEXDP0cEdtG3oLPdez/Onl/kPy4/r6Hw8SnZnonB2HHQvLKcEk27716zaDzX5PV
I1dRXrL9h11UR2b0SRRo866sq/pNLsW8zYcKobBgsiEELXg1UmbEw4xg2q6eKhu2gS90prBMo5D4
xXsC7y0j995bCspugbn9TR+Gmzzsm16vHsIIeIkYRo5kRsCPn6nqKFQxrOwTLkIWVehpihpAfJvC
o0sHLrEBZbhMK/iP3BYVCMqW9nj+tSqDH+Ec4FeziIRuvt48Fge2Ye2raKs4RHIA8dXnG+gX3m5Y
hKRgfn4JQENlTvpVqTctBvqEyw2kI0I5RsUP3lpxwTaEFq9G8fkZm6qJiwdVAb6zcA8wBKrsAK5t
oBmdNZaAdN/AsqYCidXc95EJe1awFRfGYsS6dC4bk8DlBVrYrXZzIMWn+wQ9U9pXQmp2l6FRLYdA
LyfYuIPBd1Hte3WPpzdMUkGVs5JANL/BOGhkiujB+mzUykCB03WeJ6fQjCEeh/KyP/JbAn6qxekn
srbaBkM0Aad9jVK1ir+fMsr9EDBGDnMy/laDciDKonQZ/i6nFCHt+/jmhss5Wdcc1QQ+wGI27jk4
e8pbok4EGzzOEf8YKLd1SUcLPUMbDWVUe4uy6Kqjo92jrTA1W2BEnGgSwH5Ks5DZgPQUICg9qfxN
iJSzInJ8gC6dq1JqhxSiZk9nWT/3zg2KOkl67/0sTsuTZR1l7qLz/vvzbi4WdJ91QW2uJX8LhELg
aANbBhgsqFE3PFDq6nQgzE6BsMut3m2nwLvy8rfoGB8nBaCCf+dvHPBX0V0bWIh0TlreMYs1aqtm
AA1NT2G2ZnCwQoKQeEuk6T0kZIpZSFD9Kfd0dCyxxVezKfC3LploajdYm1lpraMTjqM8qjAalMQH
NTTQPTJe4uQ4xmlAZKUFiocMvhcDqiuDjp10vuD5TRjpnhVTRtq+ohg9qS38niVU/8i8CF1t79f2
2uyY0IwO+iRSZ4+IHsgnXeZGxRf2nP6hTk9An/6/IoILb4rVAGJ3nTNdyquV7Irpnj/GRhU3jNxr
mKCqLvFtQV4WNKEUekeBntb43mhl5EL9SGUddUbz8wpzjjUNNZSEAQ4pcpLJSElPyQQPuzqME+1n
tHNxsDBjyXM97gLBVk5qR2K/jMVFtMvDyXfIFo3CzrcCYTvUOgpqlJTtZu1eXWT6jHLT6WVYYzdK
u9B/4IlEwKJ9BIGYlwXPxs0C6dhB17z3eX5JDPBkrEywFrIYzroRO+ZpPpnJJn/PStbCpC4OTHoz
YqbQvzCtDUhI++n+e2B45bNiSJ6/CbXJ+pe+u3tVBAIQ7/Dm71cYiZUJlsILakK3qqre+7iqRuW6
khBeceBcvi8ZpViMjVuD58VSKiIRFC5jU0jA2cDcI3nu3uz1Lepgpf56oHQNNny7H09yqFB8p+J3
wIlOcJtkeUoqecqsPAd4OONxSIKKn3S+bzrvbaPoqOA3lrDwsxiOqFVoSSkJ38HN7dxSQ9L4ux5l
Isi8T0H39r6iivWtebzn9lpKkRV95bRXTJFABAxz1HkZOykMw2AvqppP7dJZ/doOI4WSa2F/HhJc
jFHiwQzdNoe03n/gTPM9DsxelrtfqT1MtRIt44aHyUDbELj4YbqGiDwLN7SptLPVoVrPYwyxLvIg
/NcU+6CFoetgOpNiqp5Ivqfjaky4fvziLuBcHaYeYhjcODn+cQG4p8c4ltUDFDVjmq8/QXR5eWdQ
mB3Y3jfOc4BjvbmxOua7wI+h/d6lsxfa+UtGYLs3KIadsuwgsjHn+losQ7EcgM8lx3g1EviTHIUq
TKclB3rK3zgl7kPaedzD8IF4CF9tv816bZuscV5mlnGPu1TXLzWF8WE1226Y1LKNQKMhiDVDzT9n
SlxgWfvqGcxAdlKUD6KVdYwetsxXLrbGYu4jn35jcUNou4LmouLVjFnzeEA+5tN4ZyVLs1jJgi0D
efIezCCPsoIFZYwO2wRmO1jXnYnipqcTqAihQjmPa9CNoPltU8KyCnbGuispCv/GNrPbs3hK4N0Z
LulXUpPk/dUlrXBAjAOQjmFP61EaugIo1UbKSLAlOdGhKV+b2Q5wvNV7CguLrqWFHVzivxNZWMkI
EXCX1oSKfTmnBOc/bzPMySRvxbG6Vvr1HowlLoaiFF/WyGXAnJ0O9V3t1oMwLHgon1B2B51w8JHe
tT0PdFvE9kN9olVnCEaZlDyYPLN/WmbNNkNnUMfY8zZMyS/vHZ2hiGQQ+pQg5GFa7deJzHiXC5ij
rIpaL1664SvJ94q93Jkxht60BXgwhL17oMtsMb68twuWIrfSF0ioTDnq33lILs6ih/tNc7eeP8Rj
Mf/WKC8Gvmy6s3DU/pTwAsh6p2XbGO8IOEMDvq6WBInpeb/fAm2wTs/yGWD9BGRmuSQK92OjRyfD
VUtsSKjFfblspkfUX4RwItJfIvZUSErMW44h6sDfwNK8MtHlw2vu3iYqGD0PFL9Oi0ftDZBDJt2b
fm3sIgDCv5WpgRTLr+CDuwwNShiNkqDfJwno8p4YzpL3bqL0R4FH1R3V2ci4jxCWHUVPQIKUtt0m
n9KEQrlRhc19J4cCCCm5sfgiTigl/WpC3N6NIscSLSCSu7HYUIQdK5N05dJgGyKe90WEvNOk1GqQ
t/z9XEzYv5KkJ8lNMZf0H10GWdF/SQ6At1SoBwBmp8eAtCAlS/bHR8Ai/suMmE9TB0tn9gPdlW8B
q8wC+h151PcnQ4oBmPgCU3zvoIh/ucnk5XkaowkNmDYV2+GKND8lfWRwaT9ygOT817dzbR6jH+5N
V4kFcDfMODR7gUNPVNmOtZKHu/e+o5Cm19jxJ1lutUVQPkV2cAJDg1LuaLJkc/UcsEoZLy0Hixhd
Vmkuv93KgDQbXOY/8d1zFA4W55hEy9f5F0LYA4L+zoo5alDIHrG6PIFtxp/o+IpFA3z4B47rRK+F
pPsK3vYONd8xyCutdB1bUQSOPZEhqOt2wdcZdwAa2H4fPw/losPWKsIQthSqW3NiM1Aq83NtUue0
hcbN3ruC2eDzEePx4KUlAtsbRENPmYy1OdWhGFKBuOZ3JgzJ3/1wBM7sbqTqtWf/lFpCsJhBz/dG
V8LS4mRKdqgebP04MFDgxywmAz5HeTjAmYLWkoEW800pRETPbUwq2lggxcQqaYK7a4vaZyMYl6Ny
BH/37tMS3wNRQZAbGNyv/qi1YU06Nb0xub3hRfb5IbS5TZfE6QFHmgeKUY7yt7B1+XXoYEoqOhkA
8SjWMpjkQy8pQRD2RIbjh8Yoi8G78dINPbeQU85mKNu6irYXSt88lVV5PGaMP5hm4NMWw/bapERE
QyeskB31iuVixVIUv2jgUBDwCxawOMSuLUIum4Z13TkSjl34e+V+HPtKIX98lSLyTsrjc6rtaWvh
qQlc9nxGEEMQDOn7+zu6ANj/6tylEikOIIAvAS/Qx0Ny4NBP1EoneYt03OcPq5Jr2DpuL5Ewmpl+
yWngyoPBKmByei7s/APvZ148z4wNwXgMZ5nmTlBE0qAMwzW8HBBWYWc+JXKIwt3hDi6hBJe5XE1e
I038jRVlxsp5Un9/f3r2dqRbv9GxXqjxFIBCqXLRYrUNH7X3byzo9uE9J8cll8V1ZFtvdog1bk60
wOFHsDBJcYRsqoPecUp+AdqKbJfXLgI07E1wZeAx72ztLkGBCslPozDOcfheDUJZdxdfHw7dvDiB
+w/woEqVFXyF175sezkPqKMMwmi/3bu+o3iAL3J+qKid7mpvjr12QjpPgiOj7FQ3R73zksVrH/53
o7ISVrY5OaBWAglWRHcIxDBAlXqhH0J87wSkH2n/DwyYfPIK7tQGzbA7WMhQrhLga9wOJhnpStX8
8BF0sqq2Z+yqbYQn0IEwp7CcYgJ51wsNNieNaSErtKORbO1fsq8B9IXhZ3gYpiPgu9PlO1j7AysH
5L2w+EhXm7rDxVk40uUNYrcbdp7y9Y8t2l7vPykowD+V1VQxgjIz2wXNd8osDGHx7OCWV3bnq7Vx
iGPJmYu9rlVmItNLT/GjIG1sbSthA8TPT8p2JbhgmHL9FIi0BfbiwW10UH8LNr2SvS/yCymb7e3j
CaW8fTCLVFg/GMu0fdPC6Do+llSXJ6n1hhgkT6T8uYDkscawPaiYgh8Rzr+YoyzPzROJ4iIQijns
sMnCvJEJgwr1peIIE43/U4e8yPFFg2qFueR/e1W+11ym7Cfv1UEfD1SXxykKZDxIWCYQWx+ckSnH
QwnYC9V9+DYuAp9Kzh3UvVjbdA4dJzk5eN1LoFDUhkm+l+3vDAZULWqYQsS9x3LX9C9hrBWZOjNf
y2WQqsFxOKQha5h0u37T2IhsHxEwnpwSiN3cSYhbHlVqpva2vUTfZPf3kGbGPJgjE6pVOTR4dqPF
eFLdnzja7/x0yiDG00jQCIEaSc1phNnBxPl7fFqKMKdgSsdqMmwM0p/bDvOtrd3iHnxnN0Cq64Kg
QksgPA9wEGUOoR7TYN44xmcaQJagkJUM5F/QPWNT7U1wH5A2hUD6MNUTGpnRutHb0uHg26xnfclv
9WDtseKANywoZvPdfWRkIDX2lVZbt34rSF5jVfl0ktVWSCNdc2n4inII9FlYQipQB9yWz42IYAyw
1pgt2YLyfWT1ySdBa+8h4coKL38/zXF8qi9hiE3reSA/Op4iKrWL7oXMPslNWBcpVnoMr5UpLrq/
FHVrHLeJyqGr2PxLZT6YcNl8kpdnbppthkmAn8Sc06/5qdiX8v8u80xc/QxzaNr9SAXCQV+gIh6R
qWnWAdaApNOF8cKLb3/YvSTIOSTz75ITkZP9vNcDqhnBZYKak4bJiqLCtZHvq6WNPLK5HQczL61Q
MSR3bN47wBcFzUuDKGsslcu/Su8sqMWh2oWZkynnOhAWGq11PgxyYcS1pBZtb4Fybvik1kTbPjfl
lx3aUoX1SEG+hr0dYnIWt2CGUy+VJrIIREgvB9W8Wo2t0AW9gTqs02eg4kBqzJ24KhHFXtWVZ+7o
TgeR9orMGFgE3hvgroWZWZcP+eitnPy6JHZnmKYm6IG8GiYDZamV6JYCf95mBFLc2hMNW6yLTyMg
RdwygngPkNSJd53fUASUaBBe0R7EBJi+s4XOgf4VtF/GhYtgDOHr1vOogeQ6C+7XAySQfZUIueYN
UFuZrmBz4kr76cfKNwj1Rv120QMHC8OBpc89Wv8dkqNqwo2BTRAB9k73f8LkXxYx6mbcPjnKbqjv
ZUdN5k1r1C5U3E9Zfp4x/u+XTQCpfJnfo+7o4hDjseu1XMOLIZ0KTdveLV7BA7zGyIsi6vzRvSlL
tKO9PlE6FRd5T1TLRFwJ3bc2W+Gn3Nr1ZL03xnBzP62fQ7EYiQuxW9KCsglx1lWwUy7N9hYSVNCN
ySsHViwtmxE3tKi8vSYExfHMTmCv8SCC52PylHy7iU5HlYXySVPkgxfvKD9tzv3m2gMzdR6oH1iR
lGnXH/aK3WgLqyzdD2UWnSZYcrmQ8Gs3fmX1WwDKbbpZqonHUfLwc4uMAXALsMcnm/Fkda2baM6V
96UeNtnSqtz7os8FGzhkfn3Kr32h9oLk7VijGIEV/UavB6IHzvBN+ZA9pKV5fsufUrE+dR+dkIiT
UTGwPE1kuiq16wxV33sRkWr0aAwShgqrX5zVyvskIATw2fRPbXD+UK56SSE3u3PvAKb/sDJpLlz1
XlAcgZui1iRCFLZigePZiPv+w8lFu1aa29m0ZYBTlZ/ymSeWCBmjzoOLu9yzJN3xlcJBH0y7vuaQ
nOgrR5/pou9/pTIVxuiiS4SVes9sQ6aZjoDC7HYid7Ft55K/MYGxdwNfoVgKTBpgtEA/UmUXieQ9
HMHnyC2WWmQaeFtIVddAbRaGrcCH9KTfD/nFZbSmSkzTg337HHmr703JyvNpxHQ8FeW/zgVMg1h/
C/5CyYd8CJinzdOYBzGWq3WzE4O6fKX9h9FvPsACUIGRYd5zsR2RjMPkW1llOGwiGFn1FmaB5dP5
ut7rBbo0ENdc83Yz7qB02ioON61mygHoQiR4AIaCn2xUEHE19CHCS/obsXHb3GZya5L47CasjgdT
QFBKPJ3a34MxRhc3/MnmUFJnph/7/dc1dWl56cZEwEd/xves6gv1lcZWm0b5IjjmEqmsdAYxpWGV
kfAAOHvGiRE1yMqh3qGSdozse6/I4MVVc+GDSGq16XY6IwgdTnb0gbULzeN1dXykC5rFdK8fX6kM
9jdb1vmqtsO3UABmQ0p7w1tObVCcIklfF6/98MtCdT4iP+B/OjHM4AyUiQ+OgV0o71pOJiUb+f7F
BQzlK5n4H65TbEenUuHbDfyUzhHE6DDr2DtFcTtRSMmIMyKIVrslVRT2Y66Ldtea6Bqya6w63z4T
SdIeA6TLo3OgY9f6HiTwekhHcAho6fu9ScU58nMoN5frySNfsZNA6j/ZLB/wQpg9G3CR1bt7iXaN
w+WM1EuwEEi9vuMb2sw6qXvTM1Dtsotut+LZi7Dr3QRqZteXnF8oie4NaKYMbkBkxUglNDShlwPT
wta6hBlXRUOXNwl+5zsmI5GxCg6EiKb0spkELhwInQisBikGgzRUazAJZDCSsUiDe0IwhYWR8kij
tO9b4n0TGh6d2mgsYc4sSW3if8IhunQDHOsRoB2ndleEsxEU2Cq5PlzQoK/bIhEr2nEgdjQlxKlH
Us8ZOUMsNZb/oUaezrT3jQDilv/opbCFZbEjQZ1bcD1TmDXnUuOiFT3aJYszXj90i/JaeQYsHERa
lQx4HLR/YNqKdvZMRdzsTEpExJkyOdEQBi59/0zeh8MBywOUIpd0hD2PgI1ruu1ZmJVEbH2fe6wB
bBmSQqGT0C02+I9aYz23YBZoghQh78V68C8H4mal9fx/FRlXAdv6y8nSDEP2op9pP7kEJdEXki9G
57Mad5P2NN7+EhTjIzHtp2wYfGHz7rD5f9dnXhxu/QwPrBqRF860wSIzB/n813APWJJ47RnmnhFI
wk828l6DOw8olfy16G9im3T6F3LI4lg4AI3Dde8C15s5M8Wd3BEg39HPTKLxAh3J9WqC04/U0Qx7
MuLZ2DpLMwfDiMyfzfq+jv3yNpDEmLmEg7r7lZHmZDbj2qrb0DSX9RMeSpAdFZoF7yq+zmHS8Pmh
XHJR6A3UuUOTaKCv/fjvVDU9fRZqTCxJRSiZaSaKs4f4VEj9ovx7q+3kb/w34ExgiTcbKXBiOUZ2
hra4xW4v/mcS9pdA0DsAsZJySm2qFmqjZpOMpqjtEpHsvLoCcrnP1SIBtsAHAL3SK0+Ed7XyRmUU
z52GTFxPBA5yvi/s0kM/n3q3whOVJQRIWcVyc4VFkhKbHBfsdsp32zX2wEucskw+BwTJIPvNUClJ
SVGL+UnOwPN0Ws5GRS4AUKLfTnLh2Vze8bffnl4a3Bxm4mzUAuqBEpYP+hwQnO/Kkt+uo7/WcGkE
n8VgL03vqXjrhlicorroGBYUj+SP7CgHLR3y7soqLIoahnClLH5EyYKJaBe3XhVVF6D7ZiPu9OXw
fljUXpn/2ZRWXGiQfmICSUsETDiOGlBLllRNxLkqHR5Os9P0LRWilUlVQOOC+O4YabNrjdS6b3vF
RED5v8P+2csv2DKORXMpz0gWLNxYp6FRIyft9cuK96WzgT8xKzMMnkX60YIzGnUvJUhJ3kyO+Aa5
xA5GZURI0IXIpV1V7OxcAcbGtL4GWW+fbeYVobdAfS8rPZBuSrAfB+45686bNspvQvtiTKgBHg5M
bTHxIp4x+R6jKw/dLTYElxu82yYM/v2wgzHy87PkL8qyrKTos9D7auzLj0TjtJiCVHw+nFuHzLO8
qJh1qyGMXFkKOm9853JDvIrUxbV3S004RFu59V5PAVSMVIssDpUDqNKeNxs6d9mFh2hVog6Na+BZ
3SPxedN2fASbJJ2hM4UbcFE574chFrCFs4xu7Th0e9esL41sL8BOzN0feAgCDSMXv8I3Jh9oGQWe
lmWgEM/XJGghSs166b1WOBDM8HGg8nWIbpLKkhIqBew0aGmAsmFvOKGrtM4B3ZLIkPmM4Yz1lKRJ
zJPciN01CxFcJsvfxTLlDMzbBfNtqB6GfVrMb/sLtpzd7xJBIM1kqJKxHZXTm9RuyVIrAj/ukr1i
/a0oOHlejNHXL8GiZY0zMVPT1hokgxirmb1aylC8670WkTVUfbAKIXUI0acq5JGpigEACBaepcPU
211VP0ZpJNfWVCmYGcB/xj+q32nyWpGnXL725CdsH6sm+rFgBne58nWpxZPuS5N6uKOiHrG+U74b
ibs21rE1YqmsI5LCgkIJTITj3BR7ZQwXkQksBgF8+7IgazRF39DXnsjJEaT3FQyvfCoO7pqNuIQf
R/91zz+8YlzJs9Lsnvc2iCdlyqCeNmw0XkiK8Bb/I7P7TF9l6UJVdg4vzlyBXRhZKezQN8DXx0W4
ETD4fOS0cYdom+ayZrFhZO6VsKELiqKm4b3kjfDANBbdGZvyLCci2jChqNeRTdR3NJ/M6+rmuXaw
p7oFBEpORqV9L/w5oqp/gNvV+oY1H8ABINCmTH4QDUjGIDHvarU1YSYnoxYa8H+epWa+30WSy80z
CREYOmybKXV8Bse5+XTqY6YTceahhPdyDStiSn61DzGBrlR+Jb39lsiiUgIz1fGHtvHqVhqsJLw2
59TKtBeWeYqXlTipVB03qfrYBPNf3jxnxIf8FEa31Lae9Hg9xFHRFB7OnGuMBj8YmgKs63pPNAKg
VaLPbP65eAtSZztk1AIaw7YZnVzLx6FcwuA8qVPyl4GqEPiP1rFvqfVIFhO7a1nFzIs1B+NJMr8u
yF95H7I3hmvpm32/IAoaQq76GLXJ1o1Xc7e2KGCXznZQUcAoAJdOEKr4j+lyxABY/LOCfnEtj4SP
WwDC+xw6NFco4K5/mF/u1BJjAYNZrCOZT08vZld2ywJJ7TFb6USOQpLFPE5lLZRAJH+8u9FhmipQ
fEq4E0VxbKH3PE2dD9T0zpa0YgQisoaqKJ+RcDMgmYohM0+iQvHr3k9icykOkqmBBBoKtalhfcJx
WEE48LFujZY/lMh9gJJZA+QHhaOFVGLIM/97o2GPfGXrJhXSBRovUrQ4v41dI+xPygMovzdkFEbo
GQjwsYR5FmcTgU1I2jyb7dQk4ZZnPYgZh6/QbMM+Z7TGzIdeQyAb2VYemafIB0X2ofzdjUGTA9Ju
W72eU2F3PFioxzx8i2YzEy3gXssTCrlVGJD8L5VxPgGh+30DFjzZtGhtSSuuXwBqbTr/Ul54i2/w
wSYR5WGGsh6LqQO/f4/FWUva6RC08B7ZmfYAKGEBuz2JgYOybOVZBwywtgpa21E+AInEdo9dfgC7
QltGSTYyfQ959Ey86k7nWnaBCfXeml9jGaxxHDJsK3G7UcS5Ebu34vCeKR5w3HRcVjppFMwQFmqf
Iy20q1FJVRFme9gz7miJNg/SmvDtmyFzC88VLHqLlCE38CuXa1RE4z6PjKbaomdN3QBG8NJAEBBk
uvl31ES0i6Zw3U5FLpHo+SEYbkPJs3y85eI2WPeXo+wDby7FEsohgZgVGFLU5x+BlQOAZaikY5WB
ZQRUc7v9TdrblCXX5+9GPh9XdP0d4JjkBUgndP6G3AM0eCwHjBd9mGi2Y+Vvb4Yrz4NR4bmxRVGi
95uGlRu3Q//0g45/cC5tcUctdQCwhv883ZGmnaK3GoaDjdR+ZcgtN9p6LMn4W+jz5fNRnKPBmHpF
WPGrv01WxOJG5KS2wdpi5Sh/gT7i7AhgF+5mSUTcZ89+mloiOietNRKNN1RnVkaWeBQ8rL+/2ZKY
RimmxXr1s8SgsQ7eZg9Ykk4pdNfzh+7I7emGZ9u6RZlocLWiio/UKuGiAp1KLPcDnKRndEEwNGXr
OG8qml/AzuNBBIbB3rFt9znB8RBzCxgcX6K9MBE0Pnwn6g/Z2USf+ujUdzbmlhjnea+rbObbDFU1
XqopsdFkJONAwNTLHj4593b4Tb1xfu7iEHDJ4Jk/JAX2oDn+YAZiMtRZTctSnWmmmI3KV3sfIHBM
124s5cb+nMdk4/oSq+mld5usYl8ejpDtYB0S0ZrGkg3wWwuQxkoGDJAYHKb0HS/YO2sv3A3ZwpIT
I9yKMjIVxVuFo169qGC1SuzSfeAGFtfwm+Gv7EjTAE4V3314QGGLePwo4THuxKNxtKPir7Rmp8KX
vHBHm4PP3bBmkvIMZstp+NJhXxFsA08p4fm52IX2UH1TDD+k90hbjlQqMw1DWNpfWvF1RVvAAICf
luXyC9yq6IMKvTX1FhkchW+NJTc7bM00DNT4q8xja5o6AYZsDzh4uRA6uPT2eIQSoVeLluRPRPuz
ci4UZb8WhyqEr6HnQCmjBwCMDV7l3uhOnLcYjW6e0US0s10HPNEDucCg3198+GWBxOIHGpr49IzO
5w2kZdnuXerw+Re9ZWT55ryxNIY7zBvyc/7wPiDH+4UPGI75lxREjIvf4UYUH9yVdhEruJtNjEan
RE9eQ6xDowKNMk5x0aBqVASFhcxVekAYNJKalkJlIaeI9469h17+F4x3JfQNhOzE/fGq/+JRi0Mx
nPoGWNIhlwgDmXH197SaT5Fef1KFvv5J+JoIUS5fdAa8TYnbe2VaPRq4saqyBBOJA1p1qslspOJj
m0xK/9Q9aJ++PhZwVj6ttv0kj4r/ulyUpyc/0wzXbvNBkpIHeOyzWw19FcOHMylmaJXkstsrLlZv
KmJdpLJMvvWwlBSiuuxLOUBxVC8TYErGCatNIQ0LMAXs1lZxdiJvZHJJ8KfaRiP8uwlCBxFcueqj
MQsy3D7om5afAggcJEeaXiZeIti9oHWNugz1+oQLwMhrqSF1Dc4QBWgnAUOH2YeJyAuyshs9onhX
Yt5OOVCwwQTV2OYFC51SfxE8WT1qcB1MiGF5RlCOOuMt1N6Y/B+pB8q7hD5AJ/NnusG1fLbQfi/o
5T22O9Lvzb8O758MAxue7wUsucv6mjv/kYZNRanrNlOhDxTDcZy4EQXxh/vCR4IyM+9y6ENcTFsm
Iz8xnb5NCggOYvW7cB9aQfidRMFOKCCX3jwJCVkYcxopltGZDqfO7+Is50SSmhirVu7S+5oYJDXr
bjzUIx9KLXIofzfc4pg2OgXx4iD0i9aHMDxpKQcWm+6oiimSrLK5P0TXtt3sQoWKnXzYx2QtP1Nk
8RYlAgswWqYYP3f7gRWBE+WNbvOGTG0DEilMook7H5a/MPhC9KEiiB4y5b1qZeY4A4JxjPGDQND2
OUrEquN2yobs9Md4r4bepGPnTp7YgPCGVhEdsPJaFhlUC00YXg9iD8trqrfn0MwFOp7heUjE6WjE
Qr76ALNg6NSWuSEfjVtSSNCzbs1IcTMJLJAxV6mcmaHhE9xOCLmMJlWSue/8LdUV4eo5W8Kx1cgF
u00byugW4EDo8UMytWXHol8Y6Nq09CIPVt8tKoJ7BSAgr4VzMStrNjSV8dvdaT+mPA2ngyZvpenX
sXFY7ELrHzIlFKEnM1S5UaXPWfCj23HU7UO7VDwWxxmjAwcwymPO48B0Cm27psPIfvz0pH7uH1xF
RYfWtmy4306hs6B744WmRZRgEsfP8Qp+km7NbkO1gDA92sS6CRggVV+0YwXPFXkn5VGZD17+/BWA
EBhrOxqXEEHGsY+Upv8xFql45Xoda25t5cmP8ym5c+Arb0FrKluq2ChGz3Nm/cByosLqJTyhTfDZ
8ioY8yzFWnQpZsQ+fxDXvggy+VfHIQLI16OwyutP0WSgAWKKu2SxfP/VqcLOypxVI01Li1XVG8YV
t5njemwhvDM3/HMSO67K9+5tRs0I8+/Mae9EKz5hrAotZyHP/AekdJDTKKaU3BgzshAK7U8uFaWG
8EMXzjMxd6PeQKlsXm8gWIip2/TORdcOgOwLZH+OLfArjLGRIfYg7WleHmvsv+nmMyEJ6gFRwvi6
5aHE5U0v24ZCwYuMePFMMMAsyOOf7b98lVnz9+JHr7iEwJbJIKvVlg2qPfEZU8HGbfGClqq9LUGu
/6r0hZJlftMoOahCchC7on9tM4CemapFGxHpWdhTAUcRIgMMn90LKw2P09RKVG1d20zZkpkdUnhO
GK1VZm/zyix2a86pkDH7xc7zTKG57k7Gy271q5sg0j/8vzzKwpmir010ik6oSe8Tp9tVffbH9Yig
xIETxLYMzpcgsI/oV31VjXSvKcE+pd3MFYsB9OP09FNydJFE8KrrxovOfDdK4p/iUkV/esFvbYzS
8IpH4vmAMFBGmUslog05EZ1Y52mxMl9+EviSiuwFHTQ0M2HjS9qEgRJwxxaF34JHBaFkSaImF0iy
amQv6fwvryznXIWm5U3p3X3BOS6OOKwp3eMa7oq4Kqyws9eSsIvS1qJtJ+UZhbjqkdyRcK7ap5SC
qX72iHwKLLAZa6H/dIpz7CLrWMYnjWprWdo46KZfivXan4MlnpJAlul3SdvZhxOSc5cw2hB3ZpXy
Tp1Qyoj0J0NZqp55EeO3YsbCQFWcg6SKhbXyB85PLsPugNobVHiHZaOJtFMe4uX4SCw0omlkDJ2X
YGFZLKy0B+rlMFKx6QYVon1xQvQaBr0sHu1Dncyw2nV/+wW7tlbPDC3khLLDlQYk1J6e7PNOT/3H
fSKSCU8MS87VZuJUUV6OqTcwayX6LRdBaK6WrTLz6nxQJaGJBHm9j5C8rTa0/n+Ig9DRZTdqI8je
Lw0pE+SZpSqZk12L9WEZbfrpFpS6m9JWN1X9iM8zPDtPSot89AfZzW8y7aIs3QpLLIlB/RnNl7Iy
oOj7mvZH8tdSKNCUvzyQT0BsTY/LfxIM6MIYnPkj7YUDSFfLWRdu87jDL8D0W0p3rFtGL9336eg8
75a4QWMAGzCM/rgIqC7W9dZPmDGtfVn0824duYa1G9LeyhsN4QpQESrdL/8sYy2x05kSqaMCApF4
B5XlP62FocDC7MPh+J2YWsmhOFOaVLOXTCnv35H4o8OOiKfULbEEiO6I5uz1fvyjqaaLnGSDZHsk
grzJS4zWJwKvArv9MW1G1OCgqLBTY7qYBa2urmgq04c0Q18MQwEbfZVIf91Cx9uBjTxa36K/TOSd
EXS/PRgi1IiK9pxkwfjbm0WVfntxPy9CfzsXp7+IoQL3kPB4fYhle6rZCKJrtUD2CEi7I2Bbbmdn
JfVuYmOhKbfHygLlCw2JMZJ2B1AjvbWHTUDiG2ZVFobKGDXTs2p0440cGgvfJ9Wgj6wEHxSgMCZN
j82n665j7KQ0Xb5ZhRopmujStwMHLDOhUUKy9+Bmj2fl0sBxZEXnVmQPG3E6pbvXmmOTPDJrMT/q
zsJRfzmrv+yNJzytvSnmFzd8mhQALMleaXIYOFNzCVszxxXNhhz8o6TF1u6PznlxSyz7btaGDxeT
iZ5lxYE89Dr+XGKjv+TWz/IXLqqJd3O17SwMjl6Sn5as32+t6KredP0L9u3EDjsvF3n/gZHsi0RZ
NHGX25FnsrMD67cYaY2X5mAjpqgA7kg5E77c33gmtt2dCPG4tYuYFg6+4j24pCmel2JQRw/T9+c5
ImCm0ldOe6uIq+cg6DNaddtN8Y/OtC5nUfUbLJ2YCZxMAGq03KRwLEZ+c1baLHYdiR/uFBb16iKv
/RmeXWvYxXRofD6LDK/zIKICaDEoId2tGIz4kmsUpNT/BWHFqQS0mRovqXkLcmoe3Zu+W8IM9XjM
ISUx/ss4hWU4dfmLzrmkq2FczmOJXlM0Uo6DFnFddnKzL0uCUnb+HP+xT1wgUCDeX7gZUkjss4sv
8GskYFXVWl3RI8Ym5hFiP4XCCK75Q3dlesMApJ+J7IJLQOAofK8V18uxGIbVFxou18Ha7GJ+agvD
ss90f4qpQhcDJmN0Wut1vAE8zYj1sHuOhnR0pnrIAPP3D5EBulfyKX4paXdoAKgJEg/cz0C2skBP
RRkzEWXrkWXaE3NM9Gv9BtzfWllrJD+W0BUCwT5WCw49QLCc4/VwYCpaVRc/Aiaat/5ILdXlQhv1
FfIMiqb1C7d6vjzuM1nRYHgYlV+GHdTQ0gewGoOd1DmlpjRJN+WOC8Sr+rC3eA2noKzuvdDQR9FI
ckpR+EiNWxX6Wynt7V2g1s/9HVdO13KG0Lgy8CDBiJZeNxexk4qcgdeO0HgCpa6YePF9+/G01KSb
Hun3gsAMGIZmn0icmpbrBdiZZuIL+HK6QY+5wiCOf3kglYtJsh0ZWPtJPHOGT6OIBZOdpjQtorUI
UmFwzduumX03mSQPEE63Ov45iHlFpv90nUsDPD9pteT7s3fXKbtbacjKxJauW8ltMHOuj20IT+ah
mOPoG9i/3UMOdnRAr9TpHUWbjOnBfpeP6iMzL1MrAf+dyZVVVIVdXVNSLY1ir8ASNhxBjC63zu88
hXFprJnBbuEwfydhFo5NYUqf1ggNuFxPdqEx5ypVxFyErncleizWOWCTKQR0ot6ygfeTIwYGbqlw
WM52tC152KIRwVQ4t9aovB05sQwOreusVBdYk1sXU4+t3jBN0aWyQess3RH+70hOqdZ7zgfQBoOo
70fCDSJoGqVJPFFvfeU5H9chhY5HCm9wiQGbMXVs1mQHBGA41yCjLD2IA5T2cxpSqg6FB05Eqwo0
Mie2hYVQb9zEaPa0f+nQmAPQ6dmETklS5zyyNMRWPbY9xEu3Hjh7qxqApFbuVq9Kn4aUtxyJRyGu
qk5TmDxF/Rj53T8p9v/+YzKBWl5XEE52O3asigMKMR07yi16wmbQgekfF/w3j/ah6l7IHdo9HpmE
B2epC9xPQQLCIYMOq4nZGtMJXBt+AzShLKiWVWdSxXr60eOpjbTtJVnZ9bys1xytdUlhJXAdzWWB
rAIFzApYikTA/vXSW5r/BHeqH8yZu1ZBWv8kG183tYVptfbVgody/Mp9hDjKZ9jAkvb7sD2CL/fC
VPnxbVh9k/HFmVKMK3tIhIcBeseI3yfPtqL0UXp71Rif3W6T7cV09lvdQlV8PiuKO0yEG/F9BeUZ
AuagDOyjnIvHrZKRvGwlrh6EEIqcYgva6wRWxB4NGB8SygiJ3PjjL4A8VExi3y2Yj3PSKcc2snJb
6z5mgqx8C60M2kKI70+y5RpEQUY4gLdUZAGnTMHIUQkN+Dknjo0vTNOvob44bcuLB7wEhetMf2J3
KgBKiQjL6oKZfigvtdQXxE4F6MiagLuTWlrF7DpU35O9lJ6P/XeWJpVG9lp8edrs2ycJ1M0DVRrt
1K6sh3jwePe6LzyenE2sxmJEh2RShp9vMtCoY99oWADok4VsI90TvQX24NEJYemMZ/PVLh5UTYA5
IYAn0l0ocLfqkRW2m4ner8SsP67psNqdq8iRVRtIEGfn2V/VQdqm5ueqDyn/t5lBme0El9f0hWJn
y14es5jdmgTECtC1yJda45RaIMbqH7DcK5y4RPemDH8qOliuwAaR2FUqBMxjazsMfF5GM6gDcI6E
9DapGHaddx0/aZL9jiY+fXDYGmyyMEGsUfxw+/Gb9nehFMjK5MVmN5o6zGP+7iqmmSlzisMyrsJ5
8pcxarAH6Wiqy1ZvvN7WlkM6ikxEhL4ejZsMh/3PAiYR4tTMw8uHd0zwm9bX4cKNs4f25iCdtuCn
e3B74Ys+MiVxqBIWqdUPnvdmEyqM2+lE97ZbB1zWfXnPhu6EOcNbTpQP1OSf1+m44oh+pVzvlVkN
46F3/A8fUoBPjiKfWaVdQI3bIqZFOPEa7So7Qur8D8EHneOZxYbqgdRcXfcIKbud2WGPB3o7QnoM
17unCoUTxiEGynqGocX0fpsRh7ShvGgmjiQfIFPJp5iLCo9tQjAbYAxI07Tvu0ib3t/BC9iu47wO
m8LN8N6Jtv4kVDpU89jHsc4gjbzwgQZRwoUKGQ7NhMJJUKTeWCdQXAKsJeKYVloT5Occi2Y5L1cq
Ns6WLL3ngwUyzy727WWfqSzs83DkQlqk52hPZvDO1tEpUKROQwnobmlP//GqkExW8fsGutRwcutF
N0NwHfcUCHPO0H70UjjlXSAu0Nl7ZKgRE7IG4vx0g1ui5JHyKMUUcfWbX3Oq49kfmCafgvx6FLWD
nf/2shkR/oiBXGDhMw0ub87NJOaf4Vzfp8rFLBEhewVfkDCZrplQSYTKZVZxm1xwgxsM9Ts0Ze5w
zgWQcw8YCo7zvwiuS6wSjzGBPOp/E2mCgVR8wnDi1GkI6GOEg9GKAPSqFwTHSjP+StmOQaLjEpuz
ct0BGJHD48SgH61+ydjNK2mpzpqdLEFuFMqvUJ20C7D5qT35uxT1OdOOxrv9TR6fMAljkl0+4hD5
Wgzy9XTaTIdjrrBB4URYrM0+p/cSSGwMXVVCWkH7HHy4fhv4QQTT4uuxD7pnHrhegi6vq8m2B+X/
sISdgiOGgLpzi93AGy8La4IHNJLddIDULrLPRMFg/B2P1+KXs9COwDgEnPdWp5CZK/D2QUD6/vt/
Z1B49zFw5xzV/jy84KxUlDoRZv4yiD6shRxKigyUxqi9AK7L8iJcLzIPP9gy3PN7B1CxDasiQpXP
awMjSIU7iztvCtDWh+B5RIb2uNEadcrI9qoALXFL4Su1lNDVE6+IFvQXBKe+8MKOtPHRfKE+VgMc
3HSayGZyE1m7XgPBJ848hz0LJ7TsHw/nL00IFQsHcl+J3LgQNKMp2Oi+PBEZPvK2xJVuobkH3zLQ
gcl4iKinzafcIai5RYqNNz/jlXQxtJuV3Bzppe4T9xRzzABjBgOOHTMYL54fuC3GhBjnKz1EGKOZ
lhi239lEFwu9qRtySEw3lf9NP2JTSQGdcI7w5/RZYchBQ0TgaVrjfaS7QpVAhk2z7MbmkdKFqfj/
Cpuxp6Dq++5IpeMyYkN9mj38RnjPKyRd7S5Na6rZO/KsKz9O5RPmoENnhwNIgnFiZEZiGOlXj0y+
6ZM9IMOoU7lOaxXMMRK7wrMMnZd8pZ1k/jsdI4F6XOgwqBkrjtQIK+BCvfBh9TezrFJKxJJ4M6Y6
9UzJOluPQpxScAj62HyXiwTJVGEXqFUhDgqXo4AlfBGZU94+9J8uxbzhg7Izc+bzLDbbhU/TmkG7
qj3zL1bdP/mbY1BuZsx0kze7Gal1cwm8gEFJnhLbvr4IWIIYdd48YXKz/H5kkQ1qdZAOZxcRV2OT
MBIjtFk0k0VaFAPjPU7LcmaLG0D7T+WJwC+AgUKFzL7ucVgHBnfkBKIWoZ+1F6pqH+cYb2is0qTl
L65/o7Au3x/UTLO/fTFbxiFDYSU0lxb5XPiId3KY2U7HaaGw0Q9wyc3hJuoE79rv+SgCpHGdcil1
TWwAJIR7FWSzcQ+Q26fpMkBih1vE6m/cCvCGO9CUaJ3mpUV6zSHmWfb3Q4k/lK7njbL8bUJP5VWh
JMLGLfBkBrlpqSVqVQ3EgFZZq1Hti5KnByROFYPqYpIypcY7nTGHOEBkgTO7r+z5poEAlccJGDGn
NTk5PICdoyAxzYiE43BCWaU8Ug1gtaf6w/AgRzxWKIfNmDqj8oVa18l9VqeVFMAKYArN2IIcml8O
OJXAA9rtmEvNXAXa/7tXGZ8nwqBSYv17aSqo1mdY4hImLkbfYzsH6qTnh06GPqVl+Cpzr1jyy3hL
/CJ7apkdT9o4vCsti1kqVqGdxM0yWZ9ccu60nIReLK/CMr4aTiOIYnGApq703zirNMiNBeF4fTbe
5TZL/qqkegp9p9BBh8hd0qWj3vgi1iadZAfQj1I+vo3pdZzQSCXNMrvnHt09jz23FyZWTzFCvMLc
ZeSs+117ydIM01oaEIaKTEDnOQrycR8UoByFMPAJlfOucqVwSRyZdshOzcL45R36n0hnRX12I3HJ
1rc12RG8+XLeqcTrHkoVaIgNnyDJ3WJsUUkIQWiz4bRNiIJHrWheFdEr4KNocPNPF4Yg/STOOlP1
7oVAdk+0+nMNAQV12buYNP/9IirkAXedHh0D8qLw66ctoXFl8LA9WrKEPegtAWebuwPR5e2FZueK
IZJxsbBtzJcvEHFg9LVnXaivjLY4oWQsoGVmOYOCiRvzJzUEU5zJ3kMuYmcnKoN5DtynD2v0oop/
3oCndOTl/3HnKccJZdSy9rgpWl8yQhpaxrY/rJ+CifNd/J4TNDqvuycOGUSknqsnnEXOFuqVs6Sx
h3CFdci9R1Qcwh/V0+cc7Avs8K1dTFLhJPHxQhTB3Q3mKjlGZ/OFnZdsiJN/roVrIZHYCO+a9KED
60VurWXtuBoEtxceHN0mh7UDGtRdq5FyelKXYwvqiEaZCGUSvcGwh6W1GSA7BqYDf00IeAYABKaS
OVPDhNSGK3j01hw980Hl0wZ4uHpKEkeio1EOOook08dci1FfqIKCVmVNJnzz5SnqCJTxofPEuOLV
CdV5ZDZkdZeVLaDxAW8fsA+QZZIlVtpYDs78lib8oscZf7zfJpiYE1MsS5jztJmdMyMxm5/Ln/oy
y2rlUJZgHhYMckmCu6ibRoJZHAwo0rGpTnUakIiNOzN/YtzRkU/H+O7QCQ8YAdyAK0KcbaL2FhNl
5ocTCJGGkkvuEXY3LiYvNOslZ1lLitQPvd6+bPaxhjKc2e3/nHjYD7pNVPwlO01enuOgGrCPlr/S
iDRvrtsB1Oicq40K5MI7yngEk4VIvoOFIAuwabXr1siVaT9BVxoP7OcWBso6xYshiDf336rbJkYF
4zY6c/qW3nP5lvb7gkL0fpGU6Fjv/AkQA2E8ocXqMsNr9q3t+SaPyTt9ff3ziQ4UcKO/UCGPNQB/
bZ4dEOZ7trOpwKidxgtSE7q4js2MgqB/y8mZAfWXls7jKGrwyuk3+RpzhIa5ZcoHAceSIPi1Fm40
xYwaX2AZVBZ9juUWjXPUi12v7CRbS70XWxMC+oaGP0VCTeAfNphLZWS51xRsi5IGUWLV/6cEHEdX
CWpZcX2JzpJ4HoxKSPeBl+2Io6Am/RA0yqd1IZRJjBzcVvWM5R0Xw3jisa7RsLr5MEoke/DSAdPh
lz2X22FB94RwVQqrJxg7HSaop4S8ucTwZrf6JPN4nKiewvZ0EF0BrHdsQJpqvOubaI/IPrP5S0re
mL8qzRTElmqJR0yzhTTJ5EyN2y5+AACposmrpAtsgAb8nc7IVeTvGg1OkNSe+KUJG1IPjLzzSY8A
4xXzrACJkO6uc8ZV3UkFP/xVzVrTgp0F4Y2oAgk0IbNgR1ciNGVekyjXEz7m6VHxp2UCEeP+E0j9
0qLfIEOVdeutasIqHHVC/eM6CQ3F7qoNjXC90sKqlF9m1nz/EDClwXbLiZwUegl6acsQZ3i+nscS
8+sosRnwCbeLCKhK6UnE2SNifTvMGJOBgWyvZ3oIB3bZjAMN8KnACbcveT10to/sIO8z9Aaskbse
+DpUQ4Ljrt7pxuIG/s3lrR8NPbIWA4VI3T9/AhO+F2FctXJcLFaV/eygnKUvwM9JYn6FM2qE5elf
EQNC8+A3H38szJRThhGtz+brAKl77OGG923LaYxlABMXtKdsaS7Xq94dNBNcj2c9zzhPReVhfroF
ezBOz94+WRVmmW3d1CAuuO0v6/ykxozmeHwGTLNdyQcMgVpW9tS5XeGoIEo3aD+iocx7uUNnnsEA
41lDmBozItP7L/zbMrEfSyHENTG/EfDpjIoIPEs5sKRCLr28qtDIHWc6nOW1ZrGGksIw3smfGd5l
sdWFGvGgcx4jMRE+4yZVienwqZ1dD+if3o49Lx9/VnzwIdWoL35cBE+P6XwNz0ccOT0sDO29/d5M
BHXUtcPz+uTaDP4ZiMZvAiZg2VBRIKxy07bepJrijfsHdP/dNGwvypb5gT12zvlEAnzfMcPy6Puf
Qjbsc4BSqtBo4qesuCe/n3+/9WxP6ttkCaKOrB6j5iitOKFHom0RVQPoXZf8Bbsvembh0i8Kcy56
eagEN9AKWjzKDsBDcTVEQcdYL9pmuOi3Yxuq/Bo+HHUgIR4HrZk2aNuEsdQZqjc4FEHIO+0L0P8i
8zdrIzMj2YUJsyzZG2h1vve9ajRYeo9v5CGBp8tW2Os2rTXCtuZbs4F0T8xEIVlzXZDTaoeYYL+0
ePaJJczCjucw1hIZI/jXy/VW26qQNVRr8Te5hnzH1bomS2qcu7WcYwfHbuCp9d6pqIFyhe/Ge1J7
ppB0ujRWIzSxgjhHuFRuADQSEnW/gIHWnh7Hfifs/kCp9HHV2HVSnl8norhd3ciMRURpSnS15wTe
wpIryUSbsrGHwi9kGwmdANcc2he93G0XoRSne501vkJA7PKUV5WSHJF16klhfWbIK9cbT5TbqJNb
wRJxsT0UF0ezG47lJ+f4TmAXmZZ6zBEm+83sl0xqI2BqUxZueAzUn1fAnIhD1i6G43A+dlnxdNyn
LbJBYgRAFJijLEPFAREo+J+o80RUTuV7oVu8lD/if14O0lI26k7ucHBvwFXhY5eoyEALN7XxmMM9
vrgn4nAgCdtAfGHWwf6SeO6UWC6VC6xh6ChctJ7CYBxTa1kHlBSb9SVLDtFL4PHAGzb2sXc7uEL0
6tMT7IvoPSAhq8JtUojaWanBw2cwy5gIpnIOXTGyCyWM67188xVezOG7OrHxdcGfXhc0aBaajVW2
w5gE+o0lFDAVci2lg1KNA0OQvdsnqioCvs7mJ8H6dQ/Po3yrKh7WR3l5ZYJkMFp/4MB1wfhcGy6U
OHW1gESveqfYiRZL8G2WKn3dhIgoIdAPXKzbYtuM8+GCyPqbz+tpfmNJROrL2bVoYp7jY4MjNih3
tNDr5st5YvzoZxP7M+6oRedm9VdOMNAGjE2cNgvp4O+1ZK5sL7OcHhC9oe2acyyb6bUZLpF+1PkM
UMiQFfXOvZLT26EoWQOcVspc/ka3tkcnmI9zlM/5yFJqlsF7HNB7L1Uv2oUGFu2RGe4V5ucrWJns
VHLYqQ2pnjxVvcqT46/O3jPsZPM1BzfgeKmVBHfPD5Qb2gbDA+9h/uOb48O/UsMe8rX/qPVbIaQz
xI2B5rqM28ia/jxXgqCDg1szfoXcgqlt5rVSof3cNgNzrv/4Lv5zopsDvDYtMpFUYh91HO4mFjc8
5IbNlgKd4r2ulBdozU+ygUewpbgMkKLNN8hNt+069ycQiZkAkQg2Uc8yON9x0q8VTi+oO3Hay40Y
SzK2JVC60UHheoyxSIbgYv1cMI10Oxs9N5HidQza2V9/FfF8nUc3lQ7+oCb+1E9OwFbM4y7WKiJx
BJvQGONUb1fz1gFf01xqtdkKgABx7+gGL576fTEkaRCZSgDLwR9jiyvxV2vfwtNgugwAb9wrwh40
cSUP9C700tnwR2fXXCO7NqnYFgHVKPqH2B3SLGCYuLH/nADXk+nBW9bw2RAoPTsM5jsoM+zgpXKH
FsWBg3/M+hvXMQcqcSOPo8Zu2gIrESNI8Q8A4BFXJaRGvEiH8R/vDvITpiiwkQNVutZScGZ5AiaC
Y9EqQu3qrYZhK0KqzlRZQmXUwT6qNyJVbniXyqTYc4E21uJiRTnLN6hK0TnaZQ4XMuiT097cGvbt
QO1b+FozUidIdbkB4GtfYf4hNlBHtXsufphg5aFxAezLA7vKo6haCOGGpui1we5IGSZRgYUp6IP9
+ACL77gmJcOaYMqBdlElPahlDYsBcPp6mgy6b2lnx8aA45MmOT0+l6e3gvUs8kpubZ9ZB8UJUIG+
8+P9CejLfg775WZT+U/uCGRZpjCNGSKu1dXisuJQQj2pggzSygsOaxa5FG5uCk6xAnKgKEpzAqT6
OhoNju33vKqLh+7SyRu1ybJmTjjkeDa+jgkb2BMTTya8sxtoLM8PefSpl+weEiL4RPX29suarvTe
CAT52LCwmrEXvFFQ9qUDaS42ichJLAqe3uvnCL0TnxBesGtJNoVgqJOYFl/HAHUthzlvX4hkyoVH
pi/nkQSDTnJ/PN8ubmH6WnxaCdYGQkp34jAURKqLhGlqkBzJFVY2/FF2T7rZigFuMX6O1955ohKW
jWs6q2Yw8C2HT1/E7JPqfVJrVH0OOuCXBjlboM4PFvRwYpKakp/MLNe1p+HIFPKud6YqJTnMcIYp
snLbT8yL4ec8XrDRuXzTNvcuVjKOA4u2FVDwHjDd6NuhjOpBN5c3i9adzy0uQJgAlqngR9wqARO2
E08nVPeSoDJVJQZryzUk4Kt+Xnnh1VjzuPJhB9eajYS4xAMOATbjfCWt0u7AMt20hqDARq+1V4Ko
GPHWdrnjXN5x/plOG2nNaJALaggG8zh5Caa3DEN7tcKqowy7pRPlWKbWCdS3JzDi11CTJsPoKVwz
VTcIl5aIBq8HdXMXmiqfVa7vGKppdoVadwHXJGWnjFp78NxGKF1iW3Jhya+k0JjyHBrGrW2K6SkS
G65MRpvODrDxYRnWI4rZKQPEup/x+wetGB/QN8x1MntuFIo0OnmPggPAjFRC3yxIQtvPOHPBIV5l
nC5OzxP5/8ZbcKzwxr8h/1yCteCIEZZyE0rMQXoG+AFHmf0X00rfdj/dT87HA2oTXGfO7XesWR6b
sMtCDD2hfH7Y5/piPv3UqU1waUujK2Ya1SqHUzVmxwE1nKbLG6I3eWPJa8Aw7I5O2Fe6w9Irr0If
uW/1HYPnUot2z5y+TrCKvkCs+vR8pl4COnQirn2NeNryc+PmgRJtjfS9ZqtCHWdjdaqvy2zQARsM
Lvi2IDSx2ycYYkU0wtMSjzBWwORJ6TXavfsJc1q26j5dtdjDMfjxhRT7zR1Emx5aK9J9m5SujTYe
ThK7Z4FnrawU2WFmmBa7FS8bz64DzmElhcChQ+E86522YwlsLjuut82h/3QXEYxPRDwx4KLQ9LH5
7jRolm6afGfC9ykqsA8cLXx5ie3GmJwZ2xgfZxEuR7J9gpmDzcYYqwqoiudmTrC8B5GUtOkhkKRe
3R36IVxjnYYS2S4ovL6Jsyxuh2r8HTmAkhLw+cu//E9dvofrVKDbV251Tca+jh6kWsqespBShfv5
WLt6Ux7pv6qnvVpgBmmLKSNF7MgI9SB/GWgLguC399LNb3X/WRLe0N2RUcCKBPcnK2NwGcePrv3W
78+FGO8X1fzZ8c+nfpDi5W51+LKgOPaW3cT5M9g009t1gVWTRA6dZBWevrn7pqnNfND4aigsNcAu
WzOyhOi0e1xMrvrhNo3qKc1neeEIn+pRSLiUL+5ecniEgvw9M/YNm5mbdXXGv7qw+kl5rCYMu071
/THdR5cODxNu37yfXd3Uq0atsoRHZVZa79gMhGc38U9MmmlH2SO546zk8b8yfkmz0ZN0oVv8Jx4F
ZcPKC9wVUHidlJ2BKwDwGw74Z8D5kfxy1DyMk9fiiV3fJjsfkEi42KqLDIzt/nBEBtjIi+3Ap6sc
B9m8DVVr0CLZDSTMAZVSSh1AJoDRisWk6vwc7VjTCBF7L66lhsHNqme+QhpEYWwrSI6VUtMqWTRj
nwXi95c5sPk4fobsiM+mpB2jrFBJE4ZEM6EMJW4wFR/IN01MygWbUMSzF/p6PY42auGhOrzw8bYt
6GCNnKu6Nd0PQXlFMqBXKjFeJ+Hfk8nlWHOSZo9baIeej3i0z+jpLMm36gjzAHoxJhNAiLeRA5u+
ZC2FEwsTFTBr/OPzMbGEI0yynH7Q2rsbMyFCv2jIUtYHGqCyecT+gRrIbAnFSOM7aeDluC2BSF7B
D1soGEgp4RZyBdB4wK838hfiTHqDYHRPW0vt1OCETedTPW7DQBLe7W0hwHgvF52S7EqbcVUbeV1S
41bwU5+BHrO9F+zpW7IoKYz6pZAAzSEmcGsLBCzUw+uQx7rvMNRULe6ZjIx/Xx+HqLknd7TaZOqp
fzvLZrCPJw3EczEFkHvc+XYTa5iZhAlp4rAOhx9cpO2o1HE2GPqULFThiAW11RlDISUPQt/xZ+lt
hEMRe05zpCzCHtAG0ueSyB6qiy9aEMYInq0kBrGlyU65SW7LQvzCjB+HrWcXC4EH3LpN1ZqQzZ7y
VmvYBAwXNYYInE4Pmxs8bKMGNwAjjRt2XxOgEv0t3Z8Ta0MSz9Vj+5aBr7bzroQX950lky91hji3
GVT6VEApKDWxMb1duePMS1mevBtZ1X+IvA6tOCwId5w5k+pcx8VWSljFed4piIzMW4VM+UaXu08v
p30mgNOspXEfCt8UTgDW6r9SE7lrcjczHb3+KUMPZI8eXaWqiYtxZNbHe3iFJ9joVnvT4NPCJaIJ
RBs+N1Nk4nKdXgSos1azg8jXyz1SmSyd2aIkRunaWJkcQgSNXh2BNGNU7/k9YSOpw7DSwNhnQOxV
tR5gPPlbP1qVwoQn5lqD9od5YwpatPx+II8NBFDoO57BRgVdOCOTKXpXP+t8tQ8am65mgOzwkGTI
jm17iRFL1u5RBWA+qlwSN2KHy+qyVVX8GwntD5jQE15wljJPiob9QHfoywcOaM84p6fDcaQERAY2
A9Xvj48GVAl0PnesjteWyVrluZYkdTsG1hTwixULbuh9j6WxFg5/1Umc/XAe0m587l8w6foQ1KDS
jhXExTI5BClHkFRzN5mGHWpmYEXPl9soCipxkvoN03RrD0oyR5V0L+47uE8qr1aBC1fUbR9/y/kF
wN85HV+hEfDlY0iKOtLdlMvr5SGhFLPg9nZohWCab2TrOuiHPQoeyghcuL4JiVgoiE39W3KFzdnd
UYRRMFc8dyT/ijvqRhuKrwXD2i8hWmC7xVGh5s8YGF5IfSlhDyEpdK9heDRjtlxIyabeNYjqr8dD
Dq8S0kv3z5EgmRRBAqxhZwbZfAY7bpwF9wmyKVh7bXM3UgB5vkRh96YzFibXFNJz++Mxe/9jabXK
Dvbrh887d0nT4hhNKNrYXMbxC/MhFYB8lKJXS4Fbgfze/fzscGA0qRbfoPUCu1sUcMy88HMdh0uD
/O9aabskJpHV5dcoctt8TusEBySVoB03Z9DcITmtnD+YWdsQR/XfTWWlsJdG6eZ+5QF/gmkcrz0e
iI8Gs405uJfm13Kx2hzBT2CzA6YS6RxkAiMlLgmT1abJ/2KpgKmi55Np6RVk7Evs0kScs0MBvwGu
VPOQ/eIg+Qt9xQb0Pdo1n+EU6kf1tBiYhWDfcktq3xqGpkmr8RDeKlun0qNNjgL8p6G8ahKaNhiG
oxzn9Puo7uQtC4XKWYP+rp5pb89SeZKZ59dluf7JIW8t3eG2Cm7dAwVhOCAJ/z3WL2gfQtni8gQS
GJBmYpRWMUJq6CjfoEn4GPZ2Btq7K9AKJ/wiNUbL4wafX27EIIu9OHLzRJ33CHzSzaouF18wvxaP
bsibSykBHBeQij2eBfigIvS0JUPUfm8Q2W60EbTGxVBRU50J0NR2Uo1jwcC7Jog+VDmkcfs9QXuC
sfaivGv+S4flSUaJRPt7jeuEGDcWi31Jp+Oj0vZd1qEzDrHKtCik8Z/Q3LqeczlHJrjOAZU2pev0
PWRGwMXxavYc8dtBYOA7VIH1CYZ6rl2Uy1NyVqR2tIB/WNvKEw/jBZkD40qqWylMhONDWHHioyNj
aE718NjGh+DAFbG4OcvE7LKqOWAlHd4qQmSxJSSvDbJLnafDoKgvAcnWi7mLnXNx8+ZbWQkGXf2s
jBvu5hh199WkcgxYN0fluBb44UdJpTPiB6t+6/pPWAk55csbRdEYOizacp3frnQP9ANWUuuJrto5
WG698jbVIXGo1FjEldEjcLCIzpv6fcyhyZNW9SRa54DEzzC/T84zXP7/CDeLv2oszTHKmLeZYZ9j
+8P4xb/MAxXaCfDuOz8oI40gW+mn/VEUcf842bXU552BiEx//i5hQkjY5WlgvKWBTNv2uL8CAM69
o1MwUWzhef0fWTrYoQuNZAjXPrImiDmE+Vu6pom9tsVKhiwK8n7yga/quxP//D+RMXHQJBgjXOyJ
4EGLV8vkeEULpe5RUCUQFkLFQ/DZYbVsA48/S8wQhjHE1nkOm4ZRWH+s0bPvTDgx3r1jFblQ9z01
MchthXy71+QSk1y6rF8JzqLwTsgtGrFgOJV2U6F6DCQ1bdhblfP2a+jOZcLoD9EjL7+/77PnZH7B
fbzWHmeCQdm+cql1eGNScJQO6A+KR2dVI5srFOl6LZj0wva+F6SGV5VCNvuA1oiBZr1K6LVYSdV/
dCScjcy9jc+Ko/tY/nZUum9l/Ob8Vn+8Ze6gI7Idy83PblPULOxSQIwcAXh82j5UlxCzdPMTiy5a
FwcyBSjo15KEYXwVSnVpd5Adp0yHzR8UVw7ZIPeCu+CWdw3kkG9zheE/YV4tT1I8SMCuezvLwEay
ZEYrFoM6cP2AxbnVZz2dJA5Mgq5mjB9xM7C086XuWbU2lsUY/JmPguwEGGf1ZzodNCysry2MsfVE
s0GgS7nfF/NflaH88eOyka5xmTEYoslMJrkMb4BJfpdXQkx7ya2a8ObUifTTPy0NyTOjOMeSm75a
5X61XG9ZCqqplgWvLiVjzmo9V3PddB1IXS809cTBBLjSTxR4WO0cBU5qpFyK5Te4/ReK5G5tBbzq
Re1vcuR6Q0SQMFula+F4fq2r05g0ifUeWCCoMONHWMzl02gdLtZlaVWecCr6Ch1ofsxT++LWSByk
ub4IHLq66KUaAdAJKv/sa8SNaL2Bk2lLxa7GcELp3MllPZT7AnVNgbkwmCBT6wvitbyUTPEZShNt
lDO3H6kzvYG4AewfNNo5bssAkPwW/CJ0pRTj2yOfjOJ2l3AgEwKX0q05urs4xZwJqb6MlcNwsRPp
3S4hO4mfzHypmbi2LR4P/dyH2LQrLmRoIWqe6U9DdymubQsNmuNAFrT8anhDGCybBY5TsDeEbAhb
xOpOBRY1L9f9jMiU55t4CddE4MCtlFL/O8JxO4xIXtCctppaLwJFwDyAAgSVQAVGqak3CXSMGRKW
kZrvv0uiyomCrOB5cgRIMxSJ7j0j+ZLdKT1Xd2vDTb8X32bpTmkvY+vcBLh8ELT3YttvU3TGDK/m
rB1qUE/g7YNFi9Rtqhlsjb3D/di31CAax9tcXHkBsxkQ8k8GW1BicDvfzFfCmHECdtdymInfIQ28
UPaZo/coiI2Xd6gUTM3T+NJq6ouKpWks1/cwNF2+1SJAO/2Ko6c6UqEubY9CtZiVmr/do3hqOAVc
r2T6Nzj2vZ+OpJrgQjDaI7n7F4OTyDdQfaRQyjhhzb3pTV/pNZqJ4demuUcRIoREVZSOvoRBT5Ls
mzwUIqoCA1STcUFeYE3+Y0cZ9OdAUrk0RRFCFiQHEo5/U9zdKEkE09Upe73Win2I0tdNAf8KbRAY
0q4yKKW3pDKdF5BCRT3tOPhRKf3wqhIEs/liXqLw8RW4BXeagWPWZxo4+efKyno4VqJ6CNYuMyoy
6MutBjbxLx2JY/1HYsEWhmYkmy3Y6tW+WZCoL7ygq3xtp/VChJzWfQ8L7jqvnDrkAUTxG8eEeCKH
gLhHrDYv39Sc7O8cljO71ZCds/Wgt8fgAvRr1PoaQ6ef+t6Hsth47WK50ZlQqT/ANV2DEP2cf08w
5cpjAw5vmnjY/8cWt2c6mUBBLpALBHtnNpSL6InvvIA8Rw2eXnUvJvlzUrbGEklM6fJybC6bkFJV
1OdkbqQ8bPDaGfcoRE9btsL2RlMbI+nsQo1yEqfEYzQ/OS7VknjSI9aD7Qjm/65idxcUxblMEPHM
g4xzeTZ4OfqMXHV9bN2UCCh5itHAjNyoeGlo/KCSG/r7xkvm32GX8OUsY2YiR2dSrYG/euXOohoB
I/yvn9HZZiFqsMNaq53xS+f5m9RzBX9UYAO6cVfwh8sdatMG3fSfJ4IATcezEz1tcsaPxlVsx1fa
R0kJDzntS83LWtmN6LqW+AVSWJZhTNN+Qvx3lJUpquIH8AQRlOkJUwf7DqCJKFPnqKGw9g+O1iqe
J8BJ5ixt031qScAXU/ruO6ZA+F8UzFhJqsOF/WZn0ngN68iP+Ipm2aRoySvmNSTfJ3D5/nUhoBqg
zPn41fhSZGJaE+gOoB4oEs6yMVcrmtjP4GiFHGZ376UkuVXiZ6JFh18Z/BgFDRbN5dtNDNfPbTfj
bes5mkopRED8aXAojjBsh+ofBvEm/jZzqGRG1YeaqxgcgqMj/LDoLPOX39Kt/Lv4A9jf1bIH4DDv
SpA+SC1Hqd2/TGtplBacwx+/NcCoibBYZ8YbyY/mOO89vjqXm3S9Hy4VWGGcBnt2GCVxEx47VdyZ
RnGau0DXaLUeFdKGVeuMkAZDhBi1xpKSVaeqTId9EQvKMAtpx7F1gaSV8q9npSGXlByjBhUFxHpw
inkF22C+ufQlPtiSTIC/WyBCWej9JfmMLXP3b5ad2uQyrEZGfD0hAwLMwq35y8IL6+MlWkmJd7I3
paTjYum3O7ZsdAzCcOEu2V5dw3TGuwpwpuzQHm2iH8CXoZ8S2bZ7wj1dGY5eJUgzJ1NxcmpvGVIL
2f/MFkvBVSRk3KCn3gFWo2olpFa4V3D2QWJ6GwJcvKpPcWHvw9D1BIBdv4ItIzHq0rTc79OOQGhU
Ndz+AjJXch7BHGdgHvjaUZC6Ap0Bz6B7U6wgm+JeV/qRSTKA4LmM3fzwlECLbfR5ididI7Sgh4Nj
fpz1ot3pQFhyrrt507er0ohAoPYJAAVu5+IufM6PIGqFZrrY3EE2QIgZIZ9L8sGcy+r6iNtZ1vx7
U6uVJyL20wT6nnR2RooKqDet7BHiTiOlF0/Tj3ZyK003B5AYjyWT+F6jgR1ySZhYFgGTaYb9moCm
30omEEn4TCRPWNGeEJrO8r9VwX4JwTtVlR8BMH7s9msU5oIt/SrC5uyIYKTt9qHebov96Lztsw6g
WAOZBP6rhiMnWnKu9Q1f3BHo2bIbihFd1HlnEzWLI5HEN965pvqtjmVjZjxUo2svWtrPmjdtCcMJ
9wFhujPki54IrVPjc4cseXLMFuy+pWnsi9PuCK+b7QDOVocYrPpP3T0tl0ucSY4iBR53DrGCh5za
GepySQlb5XYBp3GENIlbJm6pQ6zhIXY0wI7nKJedZP9iFdlqxjftdchhpm4u5eoWO+OEydASW4mI
dG8z/7GU65nB39mfskFWUR2PLpJauS+QW1o4kU8XyTBVXQIFRAnpV2kIBnPqhA/gFeV0TGqTYePu
cpRRQ7mjYVyAgCQc12zMdtHbRr8x9AFZA3ogmybYMpOiVR5B06Y2jXzvdlRaViAwq+657DTm/SeK
BAPq+m512CcRjLioSiPdGRzD1INVOCmJcdp+IkkZfYV/1EQ1iLJABHVY58Cifduc/Mg3OdXzHlAl
TNTOzXpIdKzcp+BFWPrs86arNVHP1Um1v1WSKUBC1YwBlXNhA42VNGKN0JUUISAi7Mv4ojO8XLGw
b+V6ibZSiejRzhziC2VgSpxbBNbdZkCXUKHLD7aUZ4dC7Gmv2JrX7tVgp1TBYG6KzgNi0ZqY5Soe
yoZbDtIdBxjdY4piWrk840O/R1GsMYhGtT25qym/EHYMlhC8i6BJiQacYOyMV4O3GTx60yP6HscC
jZegyUvA+yf1FuWoGLFcqMv8RQA9P8yzdizX5/8Y6n3OhFBLJwMEENA8L0JiDCFnMKcdKCvQECmW
gXAudNEpZNfQjpBPHR6ye607Y08w8oTkfKX5olbPNyoUjM6v7A3yZYSCzIZsnTegOYonVQ+k9BtM
VMUqFTRdlhaD+yMKw6I7D9eQ/1q5iCtwgWQPZpbzmX6UkRwpYzl1TzqQgy8mDLk2xKwpLn74Jnz8
EBk+1XG0tjrhMTiAvuWbR+dSD2HxyAj7QdlfGtWZMek//rJWdIn8V300NlF+t4zTGiG/WDSuCjSy
LBuDHFTzdP72/YYqImcUBtjhMEwWA0J0tjmS5swRmXvaqd1cUvfPQ9jewygTXZGDc5wNOKLyu5yK
AbE8ss7otjCzptJuUotM8eC8LtzsMxN+dX0Hnig4BNqP6mwHh+5ty09u7rpNweaOrxPiRzK/qTxA
QKT7RbwEyHrQxx3tLT+7wEKQCgcBk3bwOTtrcMt7Qkqz6IVaSfwVEoBoKh22IlDh0QyKyLlKbDyl
a+S9ic9NIAFa6kuxr0fw39qEJPiohnCLA9/XNvRGjQgIHrhhScrQxk0dDE3BROC82SWOOuj5veKd
mlk0OPYx0x5pVmaF+5rpAuDwW/qV34ciDeZT1tR9Rk9tFWoahvvqh8vtEYoqGoaoT3mde/3T5hNq
CPqVdjz3EnsjOOPIS9GBC6Mf5V7snK+N4nyWiVFzKuAlqTradwlgJ3IW0Y4p8CFGsFOgtPwwvOKc
pTqqQm1JUaXm1Lhlnsc2v3G9tFJztMtGNi8n+Oi/a+3ziukUsBScopMC+pUONoi2O8r0iW/n0R7W
T3lHhcSsuK4ZlBPe5vGftabCyi7QKoH1DSomUfPCrv2VFYmQu3Vh2L2v1d7cdHONFDM/S+mutodH
akiGpGIJFJfBZhBLO94QAOEC++AxZr2SM0uzjc+Bcks+ZmlNhfKnOf1KlDI2nvba8Xov8wdMk070
thdD23ceZ1TCiLUwGnoqC2io4OzWb+GylTFFdWziAbdf2td/U+5pNVSduA59OOqB0dqykop2ZH9G
//YUPZuEsi4dl1H+tmoAazcoBXi6ISrMAJvYOR1ush4TAyTQYGur/iGuFVmAgFqCxiY9BP86V6yF
t9l0pjianOdVTP1WW2mLn4imG09wb1hb8rANKmZH1HPcLT62wIh0j9331ppUPMak+0gKXuyJdhZ8
wDOyVqcmOvA5k8s9ICErlGkMBCtfCozjgAO50RVBpL3DNfIUlxC66AJ/XIv4ZbBZ3ci/IJDBtttC
cCknz8QGubz24zquve96euJM88mKdpCbVL46xjA1RRzOtY2+fSx18d91vopzDFcxGKB2wpz/muAr
krremD+b3D8nEfflHSH4IQUHAik5ojdyw6OYtK0eZWpYHI4CD62fZQ17vIZCVOV3SVo7qPvWgFZN
mOBmkn1IcYoTCLHPSmhoR8gUCkMVAv11zbRSFx3TgU6W5RTRVzGwPkK9TRwi8ac7eFGSrCrd6P6T
jZV9ttsJYeL9ZBuACxY2V5JHX7QKISC17br9SWlaMFl9FBq/qnFpmGjGx98DLocG7p2jYjx0h6f8
Zg3Gbq44zUJ0INh3uB2MreUrpSS8gVXx5GYZLgL8Mqv1L9wwiOYdz3wftpd4i8wzoRRUYvQGsuoe
yo3hKYGJm28+6QfU/0dARU++2qRB2cLW1Y/Zqkqm5m4ZwKGRNrEOTppD6Ao4tT0UNx+Hxihetbl7
Ea8lQXstyFtT1nonMeQikZ1BjNE3n2Quboe/eWIcmOP8c+wDwWbue6s0WxacNX3A4sj6RFK/gSeo
UYUFY1x5hXJOJ7tv3JmwrGyOWTpcQs1jwT7L6AbWWv2UeMZlgto4K6vxTCRYjUMGVxVqEshJTDD9
o+MKfApq5IdFtwp8+uHsOEvHGiJs5Mg4Dr6xpSIU6kn8OwWHaBRb1/mXQl/RJjK4Qlnuz5dldkyZ
ruQIWnZMmTQkwm12K/6pPOXc7Cb9IPtg3PXqPzuyzYntyf7eoEexfq6nWmw4+nYBILB/b0iveFuu
PRaXwpH/QlOh068OhdESmpLvp3rm+36niOCLJjqQmSLFg49qgpQfzyRywIdRF0GDHJU7UyqwQYBj
nprBlOgTD0XijcpjuallmxcSiNXL1BjaY339s5lTBHQe/sHyHpbFgXTDcYfBddgBDlHNY4/bMW5w
u/NK02KE+IL2VnzdhbTppZjXQzBT89S874PC0pE5qOJkKpdqCue+Fl4KPd9M19qdOS3cqrv64rqh
1QkYwdhjxppoBluapFdqY+UJ3fRKHlLtYGboYej5zLdKgSrdzdDfKwdEVEVMlF8LhJn4Xxhsh/5+
f8lz9biPOSgaDTgQvyVoRcch4LeyX8gHL6C1pVo+L74+GyrZxnxgoIu9qdPTkS7QuKsZGnhTUymq
FZYjQg0iLxTPoLElgCpbZTWRqYERW3m0TxVikP0ymJU793X/Izl38o+Udm8NnMDDzT+IWAuHUImc
1LlFmjmZczCYQHYPmI1x1AKPnCJcmN8VhquDgTDW9uBKlLLTlzNBk31QVekYyz5L19WDUZXUgtkA
ilXLUxNHGoN4YLq9XrBfY3rHDQyzfw3NXkJtGqmT91Unsl6cWjl1O5MvnH64xmOk6cZQ+pUdmopL
g3NsfYCvGl3BfvvT5QdumWFOOUL2qCJbj+akyTy5Ht44UFYUxHmogK9tghz3NYH39X+o8VrT5V5R
ODP6yWqLx+2gPc621Rih8jsQ+DEiIYJJCdgUFqxgnmFiFQhdiSRs4m4SjHP3JelD3n8QZbKwxDtm
T7kOik3V0nF3wFAalHCVSqXngoYZyEl+pjazZoI1Rl6eTk9+uMlaKEJanbx4d3VStCigSocokCwW
7moSEQ4+rl1iZOPaK1qE7eaf5C6Ua7NbKiNOt/NbUi2sQbg6hQb7TFw5S27ofp5dG/Z8DeojAWgv
dsgRtxRNVI60YsrHMgHyXCNjHOSe4k3SiPBPNZEYrUXuxy35noQgRwBubKFC45mXrCaOmpPHMaAg
3/Mre9yzRY3ORi4ZZKLsGnBGHnA6+dDlZuHYlZle74/IH6Qxi7dB8AUrPsBl+s1Oc+UgrlFFDyVz
t6n03ntsAPwvhigIrbcsGoxShE04azXL1OSVm3rXvqP0tuLy/0kO+fciK9PSkudIK4pF4Tl7bLrj
oVo3Gz/xctOoImDmaBYW3y/RsQ77SxAEKTKWyEMAml/omAKfXcf2zeQfz9Etk3mPwj4xtvwOOnVB
gZmWknN9r2G2Onms52Dnn5QFumyX9nEWaJJl+NZDY8DlSrWxbT3wvjelgSqgGQ4UOnLFgriq/iKR
MpGwZRr0PTR80a46NSl+CW58qbzp5w/JA0UijYrA2LOjJ+L07nm+a8/J5V1LUj8lWshVnA4kswdo
uv7Bev6nwmKAJlEA9+Sfa7O19oc5O/RTv0F6mTs5gf11/88YcMdwf1GAS7GAFSaE2eMpV5zf7yMd
zG8GtCOrM5FfXoAW8pentEtTa2Vi/hqxiI+9+sx1/ez/qaGGQ72qSZ9XdULT4+gyXsQH5om8cj7p
UY+YmqCK1zhKZFL9491TJNLS1+ywGaU4CX8p1E9yZ7NZoe5itF6vznP1v80Lm+qwzPHMvQv1WU2S
YEF3B5Jay9zkxH6MYHaJ+GdHkKFaDNw9Dty3++/VQPEfBsdMJyvJJ2+/n6DoiAjD9YqM/suMh4HT
zlhfG/kJYiDxJI/pFNiFISZTrlENSJ8P5oGuff7DdlpqS+cm8SIly5zsJd58pcT9xqcztkiH5Jbr
WN8xxgppAUl1jDIAcUG/EHeKbFiSIvl0XaHptZ3AMN7J9pOvjP86LAI1dFgFW5Xctc/+U25GVFeu
96/YcNHWDk7l3xCubBltXeQij0pDtALqRzI0vvTyQhrfPPk0SJ0Dla6BjPxMEYKlvFaZ4pWq688v
X5nCI+3i0s0F6lBRmXF+uYcPbRSwV9N8T317JZj40eB/sqpZFHMSv5sI74XjcwVZXVa4o1AzgOgh
2mVMgh8k/FZxyOZEuDnY11RlC6f4q10+Eo4w/PVxuWhNH1IXUCrkNOQlrQr4PnVUsClTcepkM0/C
Yh9F4SJtXapIcCPkikoAQOl0mL7FBMgFejnWIbJoeVfwJgz/3sC3LZS7COA+GZqOWQES3BuLES8O
JTCodtxCOgL+dm8wdOeMYZr6nQ13HR4ItfSfBrJDbsyN5ZBZy9fn8zMTa8tpA5nWGFDd9aMJc6ma
xlM850n4yCeec6xyMpw3hQv/j/gWVYBVkFmPUEcFpgsTmz38zJ2e+OjCfBnDYVOTXVd+huYR+d/D
Afai6TDPHhYthdHJoJvA50tVtyLOHkiEliv0aZiO0gagSO+YfqjF9Jw4yx2Q8lAmBzgh/jGT7aJo
uVdHmVoZep6ESoCQeOymgMPZXoU8+8N7YOB7CwmTZjwjDM8QElJHH/QcEAuXxeFr6ClTeGczVXM5
e61Wb21e/JJ4GvfguRGKHYwM7fB3IWkDMxTEDj29XLkFcpi5s0Y3Etka00QTEr1CjDSfcLxU1ENx
lgzBdSz2had6G+nxgzgAtQp15sc1jOrXC7INp0nEy/WOZuyxvbu8arbHKyfkEYKCnNggwvd8ITQv
b64Hs9x4o8vNKAF9PXBhzUBXdd2n5m3S+5uFDBXB3zc5T6f4xX1pbxs8rGjeoh5JQjP24dLJcdgf
1CVIr2UXD+hWZX+psaVZBiMnZsKCwP1wtS6KHYHEDGxrDVuqJiCt5mQAraMtqs6m82GYvxneKhuU
bjVWd/JTCaWEhVXMWA+bQoMyoK8d/FeHe9pFDzcSGyanVtFaNDNRrbr3UWAtaXeZbsrVsWqKOnNo
Z6NbfcOBUWOOAU4hSgxv0KCiRPh22Yxe0qtpoZfDPVDfVoVurEZJlm0xSGUq7kC0mXBUK1Aqy86C
xtLkU4nsA82gmmXXfeFiaysB5EAP0wD8le/ZtSlCWTmjIKexjZOP0XujqQ+eMHNvLPMJywfeI4Fl
PydN8Hd2WGC6ROkiitT3GBEX34B7SdiHjWgZfa5MSeN5t3SeaBeCsUgKdhwb1UE383m8oPTyAivb
kdpqstW0ZuXF38aRUphZdK2M2bMWSfUDZWqjIsjaC0ivpzDbXUaSG5nAbQb4PxvygSUKDK6pJqso
fh4mxuBtNLM2eyrod8ASNKC94ILr+jEmZKBze5JASZU1EqLUlqKRcCkpz4zxCOhfaHmo8VgrYWqf
wwpFktVh3A765k5zNEFtkSI/YKzWHhl0Rn4n8fn6JjeI+uN40RsdSkXXk9hbFgbzdVdCrq6M6bgj
U1MYudiTUBhMKV+qHRC0PiIVi+xFzQ9PoS6syDplaSQEwD18hsXkctg+W9jqKUlkDw7BP6oxe9bD
U5uIsmRJryeh0vPCaEoP6VvrmByIVVOw+Iwx7PAWuM244y8BHehb2cxWmr6KhiEHvHBoPzN8+Z7L
IOi+UsPB0u2vD98rCyUl9neosvDtmC8/n7+dsjaehXk4QkrkoFHWIZeT/WKjpM2MEgKD+CgCqd5E
Go00+uxn9EisWA2sykMUvKuR1XbV4a9taMHreSR9MBZW0k2NBrPlMxn1IXmVVvaTVeGfeATwfnMl
dbGu7z3em5Posgru7L4dhlndj2ZEvUCcA6k4Mn5fpmD4ENplUtcuZo51627PY5q4TjnyPlpiaM9b
Pl+jmZHRQXa9n8oH7qSaQIsOwph1Low1IOYKPni/XKfHmS/eAkGFekWJ4X7jK1HD649okSF4z5HO
5Mg7PbpWx2+G7qo2mEwJffd3nyEMrBO7TxYpkS3qRJTjT1u2JkrgFc7hs7oewohsO8HeeQmwrky8
Ro3APwLh+NQAge1vurnMX8S6lFB8Jb/TTA0xyfPeyZ2Fv6/3zbNjnGcFi26ueFY7NcILzGHFDDPY
PT1dsCJ97hpWburm9iXoDsbSCeZPYMdxJcpwr0NRmzXzFZTwsKkcPcD6pDrocATFgUvR3m1h1HPl
HmYRYF9jrpaYa/YZL5Qy/+DF1ghNaq/l585yi/KQpIBtSfmmWQiUTb+GDVPwk0dD4eNzx5y+K1XI
wT3f0iuF7vjI3E2ZbZXwuPNjqv69ePHzCw50I/x3fHlY3yJvU73hVKiflyWdJb4pL19f/MS2ipDz
FVz+sSvl4ia+P9VaFQb0EdgrQd+5bLQzWXEQnpQRXzt41BWU4tXKzV+0wjCFavSn9p2JMUykKwIE
/novfZ6gUmtAXzNjeiVekaWGx1oWx6S6EWAXqtZMfA6SiRuAzFlew7KLZn9YFjfaLdQBhhfcfaO9
qg5KdZg3db7/2VX0RBZpMm88YRhHb/kGTi8dOFeHsH7DSt4F86CvPHnFRzENfxSTkP6kXoRfosqp
w6C//5XKyBn956H291CXCSHfVqMVoDt/stWaEQQyrVrf4QPfKmBxppikfrU+3fIklw7aCjQLk40f
r23CqQxm6cJTDIQWeiwI9njO6S+8N1mGfyAO2yGH09VtblZcQOV6c9MC6ZKu28qDAcO7fb8oQb05
Hg/2ZFhQveljX67aYZyHVljN5ZwIP5DR9MjwLjrPUq3+Xto3AV1xfbRAxqFcrQm4HNfAm+bJis9m
sgk+zPrJucReT6YrA9lNBZw8v8P7B4C+S8qcEd2MMpBAiDRexij26DCkshVBUe59Sq5Dlb4pwdh9
aO1Keo7m1j/ZF78JyRaTp99pWi/SzFV1xJNv5kYVQ/Kyu+9LlKlwmtLZ3W6MDf/zNcZXeMjnmoOn
hfhL8VoiuR/IiYgCQ2fnTJwsr84hWXX1z9faGeHWPLJF/pNeGqlU3sciAhGCJWXFrNT7J4FMd8N3
2tRBJ5iibvowSIBiLX1g8XRb9rud6B2XGMhnJH7HD/2lbhNY7qxc5Z62vxlb1UknybASPdJHiX1Q
yeZaST15B/9+ewz7uUq7UhdWSRGL2QOTZx+heHFZ1ccr76AhT3VhEBH3R9SufS1IVDKFhv0qGcJ9
/KouU41peAOlYptpPe8k3Spi/ynQTWGdO6s8kh41u5U1LDINwrHBriVCO+hv5gJVc1JG7fyrxgn6
vDWaoYwOT+yadN0nxswqbTT2DgN+19vxhRCOZpc4YPP8d1IKxlSCSuN+H95UzsYcGznXxLCZjaPb
odcJju5aWqGfOCWRqj8c7vpONK/LIvgBp2VTlbM1aiVbeOhTXEzCu4xa5GJezos/pFi85SivFqBD
lVhSHiurdzP6iPUhuVl92oD8Xni77E5pwkOtYsjtag3mUr3bh61EmrLDoraYSHashWNtQxT95F2o
M8VQRLXDoenchKx1i/9kJu6G74rt0u8nnpLi+olRLBQsCAXTX0NaCq7QmoUriJ2UlEHfj/GdKfPD
IqOu++6m8VHNs24tFEY/MeV+dUL1tInox0ZV5VeQD28e52tKzNiGBI0HwWspZjCwUO3TxM5MzKQa
Pud2PI254louT4MCAluRsQk4jsCvHMUq85CtxBGXSGOB/CVABJ3LTSsG10c3qmCX1HQSENWFeXcA
D1n0DiVCPq2vwkDNMLOslpovc7OgiuxMuTcuEicIJcNcB2eYroSBxXK1eIpLbBAbSr5XNTU3mAKW
fprq1OQAzNIp8ZqWNPATfCac5DKYt6ea1y50jGtLmMb3BfDJPUF50WA+DD+KaW5WXkgI3KMMYiW1
b/0MMHFDmr5c/phl9DEDngIpnvS+26UGbY2jSN/vMJa6YhtjeNtWlkteZ+eLicvwq9STDrslAIQg
BnOjZFdTUg+epoC3AsByzsTd9TWrzdMh62cFMEct7AMpKTLH1KWCho0dg1iQnuprhHpl6KgyPrAl
3MVCvEINIV0XCVP74t1YuipXj4OfzgnifpG9mHhPmf1d7AcMTKBoFso6OtlVRaPBpx84QIjp2iVu
SI7d34bqe8/NecOwCoUQZFG6TPM3u0C5lf/P1UeCmBDq/KjB4Nlf7TSwxVtyvqD0QFt44WHyL+Xh
eSpB1GfwSnbyQWflvkWsnvg4ilfC71ljTQd52Ns9Us3mri9rNXI/ZiZnWHGpkLSlBqTdxbk+aJRp
SJil00d7YBw4gdJl7JPD/pd6aBLczTrMTRwmTes/oLtqc81F1584WJfABv/aWmhJrfBRgWFmQ0Le
lIg4+VFQRO/3s5d+65LGFKXVKZiQbhXJPu/MvBIVz2fIHfmPmGMk5aULdI+pqOHZUkOTxpHZ8S5S
fMJvY4zO6Gu/dMYV2LrFf0oS9qVmL/AYR9UEzGR1PLCA1E9IZqz0g1a5X4JcMKURlhPdu5J/ACVC
VovbJ6ncySS56y02/tMU9Kt6RuP1oSr2GxlBtqsmSWpPFApemibb+RnEXeZ9MpFCiPgnmp0MJIoO
EhajN1OIsdrRC3cCe06IERa+/Lr3M6TAvjsMM3V4mHAEYonhn5UvKNFRjkw5zFQMKbPFqLnKKRB2
AbmVmhBkzK18kmf7epe5EbEaLZBUJ2rEopV7K+BS4TfOrK9I5bmad/OdVTrQyD+9MG8Ah5VYszvf
LXOLa2CBirN7p31AtKOTVo7Tu3UiPIEZ4FFf1eyJaEP2E5wJcgJ5UoLv+bDQHxjlV3cDTzESUjgu
hs4RA9tJfbEQ0PNQQv6dB4WTVYDHWfWTfBl9ALRGxVn5xapWugTWwH0vVGq5izyuSsfCjm3+TQ6U
+ulg+N3QuVO9o3n4cCHcGCGb0awD0aUSwVQT4pLXnCk+QuEvHLD6LDxR9Y7TDG3+LRMHOhbSVENl
wz2+ioHMg2Aze5he8V08bF0wMhl6NjID3LRBuXGV+5xtu4cNVF98HMwjLHjhy8mVO4GEwKia2Z1F
Zjo3h8U9eCNP3s4cLQubTIWWe9hMLjigMd15Dqb6KV0JcbT4aFdDoBYMyadmqzgjUnQlShA5nqqk
vIfnWwxPWnhakshYizOxTYogPgZC8HCdABdRGpUXk4o605Ms3Ik5avotTrBP86JP/PfEjo4TuoYO
8FfPUjd0qD+2Uod02/0TEmX4g/8pvWpOpt2cPf64X8qyPNyQ/KlYsIWx7wA70JAlb/OoAhNlHO8N
nyq+azauTtjusuMI7bQfYpgq7FpX6WBhRiboTP7Z90p0jrpdVuLyOJlxI/vgb2A0gon8VN6khUjH
NQVrmWY1XokfS+h+1jWkZlLDiiIrZTpTTgMh/OtE4Q4D7Z/L8PM+gCkkTkN2x9Mji4fTzx+AqSjd
SJlmKdScijQdqNDgwtiXU9OwOUnTZmKAzpS8B647o8nn/eTJnQopvhCPWBHdwJ0NsEYE1t8t/cWA
E6T3jO21zqO3ARhSaN2RdeQw9Kuhl/bT0KkEgEIdyNrsSDZGJCi7NoOSwcR3b0+QfiGHZHNa/JKn
qswFPJ3LDYi91jp+87JYwFUjfDKu0SnQhZNuxn/Ux2t7J3xlSh+9qqBRiLVhkwTpi1ZzHkrP6tS3
VMV85wIgzbazwZAUD84rfmQvzzlx7NEuOglTv3WtEAEYq91nWug/2/CjDmkiJ26eWJHSzpdh/1XH
6f20VigGbkQl+W+80c/eMMP+oHzsCAVN34j33QQzm/OBq5X+uf08HOTDXmYnwD58RTnywNpkNhb/
iqlzImqQ4qvWqmIWywHRNLbrR5LnsaMZqsHBcmb9mfJWJIUqfZ0BYa+7drEDrx/gPqeX7JmVMgcj
ZNpRdZMrhhJleJKoQssKN/qVxpmokFZiwjEojkbLUPZ0hwMvvEwoj555yNOrcFoouua/1woisDlE
UEjBJMJZfFDJTdX3LyI6lA0RU1i+mIOaqYqZEKpRod0RFlpAHizaZiZcM9Vm1hWOPoT+RSZfM8tI
/DO6ZbmbGxhCVJ6WG716ygVmFQ/KH1GzHrKlNUqkwcZI+mjS5tvs6BbjxWzUfKWD5Y8c8ati/LLY
hMDMWIrjYzJ8OpfvBSV/V5Oxqn/yVVSwfkYJkIEdpfxfNgCs5GFgOeVed9BnHohkUtvjm4j+fHxk
pM/HWurkCcRNJHspda5FD1cle9YobMxLaSwq7FseqcYbQoPkni6ER8tMXI5iEUqUZcSNQwBSYBVx
XTa57CX1iUJfKn5Rf/6IbVh7chLNH3JZwCjZjlDoQ79aE5bvU1pSQ8Tn3qjD/FjULxo4/2QtBCFQ
+qVbNBz48I1vNsTIGEo/pm16aToO35VsE2W/uB9mO4s9pw+SsNQDJS5djNbOeQnaItGhYffmdR5L
KQlXNCEjsrrQA8bhZ6YSNeM4abXNFzK6vBSGzkWW/ZBSnAS515lffiXhOoO8Gats4diCwUwjecEF
uYX8hwXuuL5stDGOAf1Iy30cnl/+DZRugxJ33Zzovs40TNR9SyP6RnWj9sWXcofCkKFwCD75Miyq
WI5owV3TfK5TmU/TlarIeGcm14o1wlg7x2roRihLuyXqY5GTkWSlq8mYH05aQxQqqEY2NAkReg33
rdy0LCIbShVCBbjSNtsnW8PK4NWSi2ohK82EKKo0Hp8GWhR+MBuqMTs73cUUB1Tm60+k1w/7wKKk
1oY+11+6hS9AXD2JTWVRIKSoMCffm7b3DBAmbR6iAGoFZqEHuxOG+q2rE/nBGbsE52jrYM1IIQFK
wEDqumTYdIZwDI5GziacaVQf0EIaxfc6q/IQQgFJW2fmu1XEfu+3905AeufLenVGGct1aUC90hHu
w+iOZ6ipTtcmoov+Fsacktzi5+N9mXKyyIKe9kYO+QQ4fvomUpiwW/n4+5TfTCnQbGP4LlWjrAW0
3oJpnPfTwSvreJjhC9ci/Ys86l4rgTOBsMSR9HtY7V+fJbq0/mtIVG5VuU7qqO4jEMCCvI1KK5w4
GrzutpBsWjp4E/6/92hlD0uioqvJeBK8z3qmv3rPtdDazljDFkzTzlsGhiLwfydovyXDrSwp2DhG
MICHcFrTcRbjzMubWkAH6J5CnTyZCevZVt9E20Jg9pXB3U23Vz/RJC6arQsXc/IMD16gX7dk03lw
EfVzLPLppr4o2DNfbNCK1+SfaaxB20NVQ+1EVESAvShVfd/bNM+3dpgzNd9ItSTftYFicRu2fLex
OLZ3gTBtELfhZCdoG4n+M/9SKqvreWh7pw3APh7YZuUE9zGt9c9itikVCiqy7FziVuPd4cKeGCBC
ULqrLkFGw7t4J5D/DK6GM13IiV1byncIPvs/Gq9OLbBLinSq847JbmH3QN/wja1YDxX0f40XKka0
nUGmQuJYd4GqUUfuMTi7TRbOD6Qr0wZ4LttArE2yZlkgG8bGPQYud63tr8+DRL4y998JAIVk6nFA
cYWmrUFDth3aqoCqf26x/De4VT7h9dR2usAm1jyExtqLw+veVdKmv5h26n930+rpelviKfTvU+wq
Lqnoyfp9x/jl0Ds1oPcf/QxiH+eZqTopYl2jY1WHo60iDGeGtzIhXupN5KRGomCe4laN8RNPF4YZ
ykCkQAG5ojZwRjgVaz5rCIxOxM9jsMvz0dDem1f/CvcRBNMq+q5OMM0Mfla3yr13Q5DJaRdqcPEr
NjNd9r9MAqt2CWcqIuSREPggA9OQ76r9hJViMYhU7TDmWcb3l5UmNrWqMvvfzOMwmPHDH9GT9CUy
aaYE432V/G+C6U3lSrwJN/2l/zB8OPWOSNKJqcm3u2Iby1ygkqk5hkHWv/cO6xrMvd8u1X7olHUP
va/vT5HQVJsLq5IxhMjkA861MFpmLf7a3xYKRhAQOzaqz2u6toiESaL5gOm3jPNLaiuzm8yz/1DL
hRUefFrXnH/Cq4+g+vNzUVTzCcOxHOJAB4yBe8J/pGniTLa01q19Smv8cA6KiZdu0pxtvgHR3aRJ
eXLyT+UWRNp/y/NPPoWyhvBxo5bbevXCnPJoegmpHifOQg4BGdHK2DHqnUXwhq6AK6ue+iTXGK9W
9/nYRPuEZs4B5ntM0G0v0BWNgk8+vRjug/ueM1yT8f30pYMEFJ8ji+9WK8iyddPYM7LyGZV17GHl
IEZxowaRyWMPXkczPFAzaR6d9tiqaXOCgFb56eb+8AC+JiuAUI8EE7ObOgBt7SRei3418XaYj3rN
9z383dQI3X6Z3n0sO8xJ4VY5GnETMnyHLh7T9X5Z5oD2wnL7QCdyIOB3Lmn9nLeZC7K5pSo1xFCw
NnpoFq9bQh0VPXwWeMQQqHrA79JfTnJQNZ8qTMvPWYN/LlSPTzU3K0Lx0O3CQ1GB8q8YBdrd+b01
iv6INVaLAIBpGz0MNt2Bfxd1IgecKH11Fta3sAxSCUX4G1bt1eNg5BTiuSHhUYSZTBIBMBreunJn
NOfeTUYD/SJL35GfZuf4Dece2S+wdQsCBGQAIaxaTvcrhsWYfrBPV51Alobt/j7X8a1UWctzjUOe
4SnYrqeWgIceiM/Rft0BjFtpXTS+K41hCPUN+SsoeUK5sxWN0WUFTv4vFT16ncUeP7HOONqdu330
BxFNzUyFLM55a6/dU0FkNh9RtEdete9+z5Bspnd6JrHgGaFBfH2cM3mk4sfnnIho4xQdOo+qilcj
K/m0KqPlJxsYrsthdxwczgK5/K4H//MYIij1H0/do7Kvv56ReSzje1BUietsLagFOkdkkTnX+0VR
uEWAxRR2AoefCMvCN3JUCXNErakEuyHhabqwcYsVPBHohGXTmBKrJ8d2QzeRzSmrFBeG1SmzFWN9
LPTY2tYZy+GznLtp5pdNTO4ETi9E9y0/dyLmGPU7D/hqKd7JzOEQKgLUA924Oh2lEBEbiJtrQ/sd
phzkoiSB2tvrjREZTy7Ba7ztN/Mmed9EJldvQP+ki4+OOuqF5/nmy/EIbKA/LhkhNzG8fhR5rxpz
EUVJM4vUCpkvcSSLN1Qfo1LiTr5lqI6v9u6ZkcnzoVKxDFbwnNw+P7ODsO7xpbFX6czueaYJkmHa
OW0hY9UQFDdW8ZDgCZqHRFufSPE5CpH4J4JZ3p7qZsaNpS7lxPpXiSbPSJ0cwtkxexfH7qABV17N
eL52VuEw0QkT/nqNW1OD+0FSE8b9lhYmALquHJWIfyjhPtg8YHzdGY/jzdFS6dmDsqLm4E0nFOaY
ZE1iJ+ocdrY28/FB0wvKQFQpqnwsCmnmTO5tPA/6EenXBi9ofygbpqFvA39M8FFHzWFGhp/0Vx9r
ZvK48vWJICOUpnKt0FrVCp9NyCZ4xX6hh1ssEjqFed84Mv/2rN4d4Dz8PaCIK5EeH8Fyc8wkCA5e
P0xg9lNGg+qwOBJiZBsvtQXAG/u8zEqhWzX2L7izhElm/plN4dK4n/HXSVAL2XohGaCFwwpuwvjv
NXSq4WHgK5eMX0ut/qekQteWB9NJpnqxK8mqxtyzmLHrnBoNctq32hv1sg9EKM/rHuCH97r+CJuT
rsMuBhqv8jkNca3DNnW3znujWyTbqDrBQ8/TVGau4VJXwq7EylAuf/1zce02u2fCe3kBPZw/on4G
GUaOHcYmUOM6qGOKodrI6xczRYPLyyzYImkCVyshQ2P5DZM/n0tMCYk38drJunnASrpwI3lhqzQ2
PTGQbsfZf8S5WfSQ0/kE8xBTFCFv16BNrQu9plIYiONdG4IrJRW+B5KIoCAy2xD8PHYLDhsWi1MR
oOLdQI6vyflBi2tlZMPqa3Oa2yZpaYRkyucqfSLSrRLV6V4HRF3hMnTwDUH6+slq63pvg1A4h4vm
mxAsaZG+wVyVk9nWHU8HsFeS2WnLBYjwnzbY3zwtI8QAms6h9l44O5f/g6eSwXMrBQSJlYJjkJYd
uH0i4VePXzt2r8avzP9YQ9pMMIbxyao/5y536a4yySZWl8FSzTASL8u8mhTdHDij00jzAPPapRBe
22LC7thLqCYxfY7gefxbYTMJlI8jdeGMlG8qWFL6HUZImuU9Bk1Klj3nfMZk40QoZ0C3KFnRnpVR
5SyYaskC+glSjXjy+qhHqFEay6OIkKHi7NcemJ22KXL0i8oxpSZM83Qzy7e1JtqyR0mwiXxCBSYj
apR0j2cb7fOIDT6lcJaS4KVvF6/EOoq3dNyitIscU/NryinRI7Mp4y3v4PWAaKap1Viz5ECntsUq
+R1wKrcNa79kSNKRsCVSUeWJqx7kRQPthq0fA/RRXkt5Gi8S1H/BdlS1g12Mi0MDesvFjHnn04T/
9EyovtMFuTsqLnN1T1GbE2y7bYQGwc+nZeMUmfgSTl7aDzpA0uitZPDjnh9TbW91/0O4ayghyQow
NKZCkKH4qHch3FtTVMR2pZxmzqfr4l2R4VW2DJtNRpl8CS9uTQH7qQ+MTcIMuPeA8sVV57q6C417
iDLPdM6HI0sAllEwO5FqVgHedWNZWKNIL+lKQTaUFuxoQ0ZiS0pePPQO1rY/ZM6uhLJq5GKkh2rt
HCGCw0nHj2uEJr96LmVqVGgNVDyPix8n4w25N3EZSnuyxX2lfODcSvyqFGje08ZnR2i5MuScdWrC
okcePK8mQd74MI9fflb/+2GgjswFBOGmbrrer1rjIy4M+Wgq5O2u5Jl4bGp+Lddess/FrFuPFdWR
0gqNwrGjXuZLpjYg0QrIHu6PtLONRByjVhSuzqKGDX1vE9IisywYxNrTn8gZsOKTWNwjgfwb/424
a8WdIFnp+E582U0JUHsMwHT06E07zcIj5Dlj7gMSjI1/eqBh2KxUgVZJWkeJ2aMUBYvPbT5ALw/X
KnzFCkbWYKK3OCwHGlptF49FdHG07n7KXZ9FxtiF8CDzEPNINgXELwpJTeFobIolFCvrJDBqblHB
s85pXQF2A21EQFJEi9jfB5OyPD2WKfMPUTXaPY6//kWpyxDdCtMoHOIUwGYkJ/nuGD4+n1FeRtvP
1qNnD9YSzPVPB8BpHiUOtvv5xMkhNqazQosT31SANO2h9XEtC6mdNQC30/4jBsIEkw6eJxA+st3u
OlImm1G+RSe1GOKGzP1bfgrqolInxcaeg8C6evb4UhroHPffHffL6aUm0Zm82kaTuK5x2dPWBYBI
8oqByETm2CtWp4AVaL3CUpgK3HeL72oKT5IpLiymokM71Ep92JCEOiCywHv2Skgnv6Fb7X0vmkEa
z6578sBLO2nGguXt+0bb7HXI2EX7AJgk6XhhCTrg1pMnoHSmEw3NGrLHCXjt8PozCUvmRnDuma9H
djIv0ujeGUFoohvrmF8+M5DVdoBgmrDrWGSZz33SGQfdjOd6yOP1mqFKSKQFhx2148thO/gEDOOn
BfaYX9pFC5TZaoxpybB1A1HO+uQHoQVIea9cmFH47DqySh2SAJ4Ot3K8zZEK/Hqugue3H8CcMoY/
E9bCLhW8+dgBVurtKE/CGqmYJldcCNmR/U2Nqx+xWrnsNpSExWN6l4ewwRYtrQR3LRFrnywDy5Vl
A/Es3DmE9GhiJnVyDrXc3QMyV4F+zsHTYJAz6rNxBeZOV91Q6sPGKRUf6itlIocXmCGpi56cKQ/0
k1lwL3ns5Co9FK4244r26CiuOQvAwx/tVLWT0FTeT6C2cnK9v603138jECfjkdA1TfAbiYXv873e
yRNAgw1P6dVddCR9++wXLRDZyn9SsVuRIO/9EcBis9er/bpoDRXxsLhgm7GlBOD7XSGGitN15g9F
Wqrh9hcbLHFSCUAIMM5wEVTqw6zpesoigjnNXgpjeZaF6ZVu1vuKPLVcuompA/VmyNY6ZouWMoT9
KEW0nQ9LFQu6iMo4UnbYUgI1hYJi4KIJbLnM41ILkqlA9f/R8KIScMy4xYdEEcTyW4414dJ8YxeY
fnJU83yJd+VnwsuuLMxFdZojTq0dI/hg997J3H7KLK4HhUf87VGv3tF930RvX/bWA3WRIlyIQpUz
rhQ3pH/xkHoCLzhuA6qcg9BX43nyYfFeo+KMnKaqvLtZNPSdv5ABPjduZIlXp0PgdrPcj7P8PPIE
+H0kpBBJQVVssJ6fR4mBn/5Q1KjcCPPwNQiiWULyZms4+aWSwczfKRPtCKP5Iqy/OImeTn9GQc5r
8RVe/8tbTI4Mxjx+YagQo6tS/a8EO+h83EsCNbJSLcKQyskY9RohMgo4JlCzJHWfeUJz0dHXcULp
2XJNcfwak8pMHMI+jsV635OiInJp25drQXZWPoDyJrmkQ8/1DanSctNEorffH4trq45AQoD6EPHc
Ar7H7EmRjFIFquKCD8QhG4SwDRnK/A6cvBe+Ay36Wcd7KLMQtPYZ6NfeS0yF0eXHM2Now7KsTD2x
XTowRl1XSKLZ7VTYoCQGI1bLUTV0wrhq82aEQB52WLIR7X2gf3Zvfd5IkH4GWAYttC4/s2WmyJeP
sbLYqWg4CcTlyFhid3K76YRMOrBf/CQZhmAbn5rk/m4BXHuWNQVD7im+HkzFiM5sUCbPoOw82qJ+
+wviBPFnoXfo8ZvxFWHV/yLtumw3maqkKEq6E3nfuX/LMcbAaK16bmZZAMAClVHMHQxBgZ5hsYKm
vbI5S0YslTzmlBEaOzI2sroukijCeLW25Q5Pz72NOvrUpDKv5vtTwh5pNkrzaprbw+2Wt0Pe5vpT
9R7ubRjgaKimUup+v2r6w8sGKPdHG0S5fSPnzQIoH9SEflpWFsVxO3/vsiGEdeGcKb45I2Pi0HU+
piwM5YbiJ4htk3lOCH36l0z3kbIR+JmpYNhXMbcQeImPtRkCQ927TvrvB8qv+PweqWr+rCW28g4s
53k24NExGTM+yvweWgTi3k7rUAqn2+C1GNxqj2uHD8xEQTI0g5ERbfdglwYBP7373mMjUYS7JBzb
NikDIwr0j54dNSjOKOFYU2jsPyvT4DV57iQgwP35F8Z63c03Ox33KfuEyu9hcJerDw4/+ER2WGCX
gvpxsjXCz9G4PvFDESRNrOLkuMXh2FxWyZTAOOs6WFo0OU97HMRVpmFO1broYugMI20/t13xKPbm
VlEOePhle5I3bWS9V7pQWHf9tYRYNhvRTmrPvqi6Y0bBfYyvCqYles1WIcU/zb8jyzXO1uqYRkYK
wS7cMq60u8DMawKXtycEaviblAITHO5OFYW60iXRj9GBaV1M6jpAPxhW4SDJGuNWzxz8y+QcreRS
9r00N21EZD/5f4ESUGPCg6xDfzmaBRA5RMifMihfeKZv22wGOHxtX8Xq6eMMlfE/6hnvfJZhcJ6t
73GFcHUqHn/ImHQFw53J3d5LBW1HoS/ppURCJK1bQV2m1fP5E46rFVz9HqFAJLPQhbKgivlt7yVe
ouQCiutvoY8x6GDUdOzDuSefh8jokhO8Ag9RB4O5Dxc5ZGrFEvFD94axbW9Llw2p9eqxPM6udqzF
O3U/Yb1iuRayESKQ20+rDfrDnWm1nc+c4laQRkH7YN8Lo/AzyD65EJ+QnCxxcIja3Fku+hLQm+qS
TxyQC6I+Co6h0lkQ6a3pRkIUI5QXKhIjPROBKBHb13Za8tSEYpLfdaCuEClxMEvPwX73Bx9GH3CN
/Ljgt65P3PY1lmUaFuE5EUsDu/ds7NZAVH+1CtUrRUD6S1LT+wgqKFxDvSqelpIGluMfnOoNjsC+
JlLkIhDJkMEO0RI5i+5noK1YUsPpOe/29xxMzqR1SDPXq+VOdqHRBZ9uas6bEJvlAVu9BkTQ2H1h
3CU7GBjjSlI5lQzNBpVnN7O/lnFDGfmaW4JIkByvk1vR9Gum3zTyjJ535d4kiL2myLsWH5LUfpMd
Y7GUkl2MIe+U/dMBG6GORbHs+SD6AVkp2wvUTfxLZ1ir+a8ZnlVqX/26GinQNzc8OcLrCVdHWLaL
SOrNJ8y76r4DrZojWN4WDRlWtW8ZAic1ko0m85OkvhPa/7qFcVCbNvQMihtq8+Jz7DYiqwpppab7
pGrsfiXHh/TLO9tbQfLMqZQPQkvhjtmg7HEMc91zmHVvPJhyRTIaIhDwCMLejTBoEMWsLRGVa+vo
qC3A7T4rFhC/pwdjjKwgn8v1pkHXDSzIjYg8TwvHDWvCUHGeS2F+eecV19CSXD8WxVc2a4b2rUYX
Yq7loGKuIg1fWqnBVD2mMjaSMcrrEUyBxAhw9xhz3O99vFCeWcSxsfIBaaDZTv4tE9qnTH7NHT6o
tWJLTpFIIu4e83t+ls25lqN3KCBm1osdXN45yZ/yj/KhMJFewdLfBkVlgQI8BmYBZkkU8Blg2Aq7
Ur2zVc/0GLwvC1G9X7Z8UdvqECDCDuQqeX7zmicvw/rNdwqnrN7sj1YTDOsn5trFCleLkcbJQ7TE
14Ggesyw6bed7ckW96QaVfeyW8DwOUm0OiYiWiF423qwWADaELpwYFe9SZhTAvzmRVObooCgXo2I
7sG9xy3X2TfnnOkicP+TwDFx8sEogbb6mrqjP22T0zv0+ZiuNDIkzNEvpq1zoyNjmr3FcBnib10b
F106u1eQbkVZT4k9E0DWeVlVYz8GmOZ9L8tFEdmj6DmRt/tOAIZovmg8RyShbH6jr1q0a5Tyt8fw
kX2MMVRv0c16Pi/D+ogrFX9MtNN/2QneEI+QgR2fTGrQUPNXXUhhdfarfC2NT/5G+JZNBXXZ+U8G
EZ1fc1fsN9urxaMxFFs2SnRCEUj9MQ6wrc4nOzqPGGCfOb7DsE7SaR29PK82MWVwv2R1MT/89p7Y
9TPlX6gfMn0tUw8G0BhM0pCZxMR/jbNtpRkHaX5HgvlITSyeOqHDvwq1eJm5NXfMReSEdJ/khQjR
bTKpKOgF7o3DJaRriUj70f70LNEvd4s4ooWvDtXm6+8qwFRQOQFaG0CD9fW1byZfkjtAafp7YEFP
L87vXkmpcGsm0vnXBo7DF6TirjcLmskwNQQ/SVBB/g+gCkJH6o6rq23ldmMbhyrn04OePp5/RG15
zYozNol3yq9Q3zioSi6UpW0Whn62+gbBjk/yVycZWheKVvHdiwvVCffGiTwtjtCKYKK0EQKAUICP
FC3Rd5f+HYfcVz1LBJN3T39dYUYFc86FJNpzhxQMSahdyI+cVxXto+G0dSgB4bO0vYufUERGzROc
1CiVTSSnKVmjo27ac5LI8+jfhWd3nNkAZKLifmNe1WdFu+j+tJjSMXDrwQZ3h0jYeNPi4fzc+qcy
c13Z10bpMDK6UD6dW6nNu94AkXf0AOm7ndtYO4T7Hm9odQVYba+q9+9iJw9LGjyplyb28kLM5q//
JswhRPoLGb5YaUw6DbpOm153PLzZWflHqjQIVNYguP/ASl/l33EnIB/wOIcfGp9nSjFD1gWb00bJ
79n6JZJXtiFESi4qW3hF6kJmvg40B2Q/hTeaX8MAzHkwYhO7UH4i8ZahvrA7Lpj1OcAMsL1k3VJx
JrNiPdpeN26iudOYrCnlcGFEsxwgIqkrWV7cFswSVo0YfBG7HxjAl4Mp5YXcNUbOrH1awjX8Nfzy
yJs3lA9HubsybxR8wzW5XG2b/F3pB2zHI4Anklkjh9rrAZSubYuAEDd3Om+IZ0YtaHHiXpVbsUkT
uSDN2ItBootHBwaVHmO/Fc5xtyG6GRaOZjmGCwpdz1p9331UujBHd1V6+l6VLNDIFH1JJq4wA2J6
wXJPuSBmbTok6nh0vBM8J7i+LJfgq90bMzPboVQ7QV+Nt+4LV1Iuc8vdIREgnTuudeyW1ox3xbz1
UKAYcO32fmypu6hoQGsHX7+iegXxpUoLg4H9U9ELyyNCqZIjoDqDsd0Zb7VZV0PIlPMXGNYf2BYh
4H/yVbehhq6CIgb3UT9gEAR3S6bbKxhEDKdT0Hx/RicgEj9cmu7JQSnSUdDndq2IyUWmZsJxnij8
ft5kJx/r4GGs+jyLu+8ke9ddmcKYh6NOj0Ts+2nWgvpWCDbVWgBd5RJj2OmuIHPHpHJgCKkweFQE
lx1aa2/XjOjGaGRADtqYgx+SRSW5KcJ9AHytS5yq90oJcb3MBEIYD/l024n+lKdy4kf2LyeT6UDJ
lFknxFuHpQxp8LOOcrmIAcjQTnFr+z1HrtpUmcLhK2/rPgPR2ACFwf3D3eoOwCb5z6SiuLSz5ahs
cWJ3FPoGV8mnmlgx9/Sdn446LCaZRall6z2jQ+askEzGO/GUavckKUYxXsvK5X+ceLJM0qOGWEcV
Q5VY2Xj57oF0fCGJtGBxoZKzKNneBHnSxH5va69n9t2w7Hee22PYMu7vCpKNltFPqxqExl0WR/0O
b5bGUYEsUhoGRhSZDKK2A8i3KDet815GJCYScCzG9i28lENwLl/9H2bv+/MHRnESPkOOk+6F2mP0
9uLkN7fEB4X4lGUBv1Gu+OTz337aHl5b6D5QvVg++FmbYMaqZBeSNr//enpWOmhWi7wPn2a8dvVI
1lIw9BZ2Qsg2lVCyEHEz7QR5+xr/Vkxur5Y/CglM0xrsvdwmzT4WJXu4gQ+Vj7JJPEDYz0ni8wZx
wDEjIav41vhohBfOxpLdq5NP4qxBOx0oG7mZgNQneB7W9WK47Sy9Hg4uRm1Y8zhx9VPXQWU8faxi
ziomM+/aAaoQwmQfUMssRMUFj3WNa7QcpKQqLf+p3lFW9WUkurYUXdt7991M5bP9pvczSPe/MLO0
GfQPTgCGrBu2HbxYtPU2BAt2trJhl+HmskMCUWvn2F/UY/c9rAy0s9lB3Dz5R7OAL48TGiAx8ul0
aWXq42hWywGm5IKViJWsP1+cQUYZkT8UKuUNvvcpHpYOr3usDPYBicgf/EF0rJLSNR47CDVAuENx
PZfMwB7TVs55RG+bKI5vPyfH3hKHIgDkxsbcGeSX/Y/1TEeHmv1sEbcVM9xmcYMWRMe8YNYI3cix
fGzTTT+KTOn6IP1bwjkMowEMcdCz+13JkDsZltKnaehvAHT+IT8+Cm3NPySVAg0YNnsvgnKk2qEo
3JTwnJzTZp+aJOt+nTuJhKm5AaOEU9o+Efng2einG0/TL3aQ5O7o2bVEqG4TFfwp5bGGQkHW6QQH
kuXmxvU75+b5tp48oR/4nni3VmWKtF80YT20zGVFjSRuPNUnyZ+4zDTVYeyOn/JjQZRRuW3TVz3R
anlgXVIMD+xNxBGID4iYDGVsOb5+HGLQ4cdLW7eGwtkigXqQpor/jK/bmLBocOnjlgs76LE9+Lys
CQmfnEuy7LJzQAr7jF48Se5krMrA5meZFmiL/0A/APV4KPmj6Y/Q8V4Oa36RqrgdkmC3dMTxP8UZ
2VZiCpAWmeNCfvOYZibSiaLweXfvGrR9uszHjFTfxgbPKasbjx1zFWp3+UYRM61TqK09nXvzd2Dq
2HugU0gCtuBhf+ZoudZqqS6T5+J6aDDZsrKpHlinTp49fkybqruVBgedxDXrjEtYOn2gGkGeku14
Yq5LsMPdn4DzuWMkPPXme8OaKwQ/I3f7BHiX/K/YnFQ8dE345gX+9do2CkEaz5P33x7StMCCvcv0
Fs5vJ3IWTJdKErmRugSbIY0mhF1zfWaIuDqDIfFB2Bzov+j0R9WT3R4IG5bqzhLZyy6YLtOBrJ7s
HPPxlWTzCJVOhPD4qesKF98yjXxbG3J7Awhc3F9879Xl9skKyJ7/nK9ru7i7rzvq2YdeTsrPmHtr
10ISAGlgItcdCYUg/IrWzjACfgiKFNh2xD5biVPv9bH8P+BgXiZdgcIDWpOIm5dLFskKYN3ptKmY
KtvfR+ZsAlTY8hcoRkVXd9BBbhbrUNrsyaSgWRR7MUMdJJIvvjKygHMhebRzH5EiLNtyct4U8tc7
W5F/wYa+Sv/EBjoVA4+LfKOdAOGSfzrtg9rSaVIgYfX4/+SUtfr8nHm+9Duh5F9Z+aDOJZaGF4J+
90ltpa8lkSaa/KUtQ/RXWNejkwSrtLX5vKDUzqXQwO7IH1pVnwI4No6kStz+U2JEFH2ohibvY3rj
0hGZos537Mw69Ggmdctol258eJy7o9Dir98dmzqBXYeBaGANi/VD8qrsOQqeHGdAherrEUGe+vp1
l7Epvy09XFZ/KA2f/4C5DsIOXjIckS1qJRMWROnUWghIYyC6SkVhzCVwtTWV2Fp3cm7UbUCZi2e8
479B1qaSp6Asih9SS5FXsxEfq/Eza4E3kLPDk1QOowUNPchkdgg2LVv08F+vCTisUTMuHfqCrtoi
2/lh3R5AQ8WAWMY9AaZepy2ol0c8vnPWmR03kv3diOM/TNV10dqn78WckWU4qHlopotP6ikmSTMR
MPzvCcbpfgDffic9tuRUTPoqTQfst7Hki0WsPtdGPzlWImy21TDTCJ1rAeytNxZRvGNMIM9sRvvl
aibmIWRc8rY4ncleI6cPwMKmchGqZQSIXsXe7ywt4E29iKHQ4nIS1ot4EMbVlgJBxZfCJxyiVMBM
6qRMH7nOPhlxyDLZgDLDXzTfOoufxlARlpcqMM9rCYdJN98chwS2jAAhBRbeSPLJ2UJZBFhzjvgk
NPX/lY+vDTFYdPaskcuG1AFrPrlZkhpQbCZT0cMXYD19nkIsiN8W7qruHcvbcWQXiCGZlDLiBtfH
TyUEtgm8w0PA3u7rdU2+lUZ/H/3R2ktaNnu/1979HiF/nhy6hdlmjAREihy6CtK/zVNBNGR9R502
4elOk4usxZC0Ljzd+d+rFlClulAXRDCDDv3Zzc31KrXkmBwdN6TyJb0HGZ+rBic1U4M+9yYjXp8m
ybO/P6C7QTcxN/YSgmT69JLH4TGaFZasMXQuECnZgDjF6H5g3ykYc+S23syQcuiVIunfuZy/ncAA
jRibKFzljcXeBC2paygw2zPpnosTmY5H+GuKYCTP9/9ZCags5KFoEG/+jLOqYCqY0E6ged4LUQ+J
bKVShQalKUfjQDfvW2iiWTxnoOuRi7CPnkHtJwSvrYxjf8uDx9O/hrK1YpXClKTdUdiGfJxYgN7S
aQVDsZzHLreie1JpqW5CjudimCxEVK6VYvyypoRPpVo/SZHts2js7bSS3FbMisDYlDrmXbC+vDd6
nN/c8CJLAoXu4/Ev09Mvv+vU5JoHCiOTD2tMzRHGIcQl1ISs/FGCe9UZqHzF5mgAKc5qbqFh76y7
FJSPMfJKWft9cPC0a3PpJwmfxlFFC88u/IC3KE8J1W//gu0QyAngf5od/MUvs9yXdyqprrS4Le3T
qXW+y6NInroXGd3kNKlHbCCvu5YSRxlNvjCWpluNZm3cyer8V9cEbrBmM7rPG2AFcmE4drn1bUKk
EkUkWbxVmyFTMH+QW5gQT1viMoNvcgAMOHga9oIIWvOAxIvZycruhzc4/E+VfIiDcr2e4o9uAcFU
4ijQYdcKUVHQpOLkHiTFf3grahEDshz15iwuKam8AtD0Kurbs+lmbuaPu6oiiMO14XdU4xAH2bgR
0jTxHAjR51nfAyi8GVEngmnKukKV5oFmo/WCZEcVX35QdM64zD9HkF2bSbISgncZewW6v/VD3zYd
vKxjgf0v2EOqYQJ/d2+cGfdA188Rg8H+ubxLXKvwMndo1R9NDnpz0g5B0mBGwGSwjmY6b8Q6BE0P
+YEvK23gPp65BiMhOjSTa0lxfeeYeBFYhZRzpn0KmlIdqHWf+seRXoAKx1C1NdtxK969Gohg5gJY
WzGeqFr2/cgJg7YUAm3L9F1WAE5uwzKHaoHmWcPNBH1mtm4fYPIQDEoaxaZ37515PsGYegEop1kt
wQ95kRd5pYFTRXH8gXze5KSp9GeAWvMUMcv67eU1DjgeaFkdfy6qc6+7W94bi7U6MZJQ07sqgIfg
sEP3BW0laSQE44I35gMlTRDU0IYy12YblhCjihNewmfxFd6sCSIMPZCvaPRARszxk7MA25CoLe+a
a7raTUEw3/pgH6x5yaJECjTgdb0QOe7QHZnBStMsYJgWiqkKszSfNhAT8nXt+4yXi+i4zE2P5rBv
51L1vyLFiYu6q9O8Q9uEQHtn86K77n1CSpig57pkv31D8VljeyN2WdIfV5STxoiLykQc6lA0o3Ep
ttrHUppsGTa4y/Ha2VrySn0m7227DpYKSYbY+MRmF0f1zG+/WJcqrK4Y2UvcaPh5B6SOX0Rr3Rnm
MJbZYPBB8uoZDlbNc8aeIGX6LaVYYpAbmdn1QsedoPYhMrDAMzqaynj/pAnPmQTA1mlc7uqHb+y5
/FNVtVokKKSlTGptHcAdAPJqm/BtrEn6F7g+mS8zx19VCp/O5WXbvC16wsCJlcZesNNMlFLhCXJV
GCj4MS+M/ijq4rW9e8HYuUVYkUO6cZaOw1orFazGJ2kR/WZIAhazDsTKTg+ybBIm+LQ5nXP4wpG6
AvO8HVZtK9haFCX5tSNDiRKgB1OmYvdGchfrzFywA+SDm7PMSkX0Lu4SDToY6Bxu5hVZJ7HTSCsf
J6WU0Pd4OSpGg0RD3yXOVFz3IC6CDiMntkbzSoHhIAN5iQKoTw771v6xlejk9GKkVWVPAi0E+E6c
VZIwtXQXVwytOeM7Hz9SYZHZ2TH7uO4138tOJzfGmjpY14JeAJosX/+LexBuNDM7xlGsG9Dy3osX
NyJSYRJmcwLXh6d41xicfcGGnUoZ83oCYsO8x/4fKSLWlTFMh8Y7SecYZ5mRIPsnleTU4woCDc0K
qT/PUrxPejgAPOMPV24ASPToOWxd5CE+qduFO5HV9Sr0sojeHyR4hfO/T7G1evbay8mksy9g4sMM
MCppGoWLY/bo2i0dwuQp3nvzSRqdz0BVs8vgfnbCSvR3ltBNtDcA+vSyWuxC2x/wr5T4CSQ+wu09
pEHlDh7M8CWVlwMkp4/cWpP6qdoQaMbFbbMJNyy+BA8QlBy9AAUNYK8a6DTNH6BUJINJNvwFaAqC
nMMulArKKmLaqe/Gb7gxpivBFC5/UUl0SAUDcF+fhcz17uMUkUi9eSdk5EJlcD7MeOVPZACwbwve
SDF46YkScNVXpv2TwLLuM9Jy/wkixF+Th6VISsniR6ODJshDydafBdBwE53XgpVAgco2TmT8Z1/L
mFy4V7QFPzcTE4M/R9lJOl9x+d4jPiJ8AMNNOW2oYrTYytcprKiLhHqCgYSRDP/vECsPcfREhHCK
naeaFDN0Q+tH2WJ8IWMrhxM6GdTcOL8ukyUcj85zr/YgmRMSa6eSQcHLFN/WVP+qVlSH3U7BUFfD
Fl5IFk+wauBoAS9kmhrFFaAhkRGD4oDcqNNI2TjqEMr6+D+PLLXZ7BVNVk/qTm1xIDXLY8SxVTLx
ZMFPNHB+wV5dHp4spMUmWDYuz+mGcKB4fpdZFjFYb9VysJxM6ecDVZ6q81keVtLzeVbKvA6DlFou
GY310fIbMJzqA7BWjTPE7kIDvJUz8j0kB7MUuhHZKZq507c3cpju6fBQBCzF8RVcqr8S6xDbiOlu
rUTHYlTyyNchV7b77JsQmLgvu3a5VfRygdeGsgub5dXamXAJesaIjoltTjrojtAEhFjGB8ufQbUV
HcxXsjF86oemZxw3OxQWk1EtmM3A+KF28/8g6b1GQ+OfMlnREw/Jrx+WFr+Lhq4OwbOHJUESaJ3Y
I+vRI2+B1NumEpYepkJ3JcCZcdH382a+wd3hRcNWKnsgX2DLzBrmLRB2sPz6PZvPfa8CXduoCb4k
QlyJCZsHDQqsm/SkedDEWbGjjWMg5Ahkt4iKhRN2NC8xJeDEQyjzvV92kQdBq5iszoFyPobymLYw
wjDJzJvvRTW5Vhf0xvJDXb+vLJT9xxlSH5AmBe5axovaBvXfmM3E0xIzb7WF+m/ysc4vlaJaSYtd
vt4Pxn8YEw59jFwNEFS256nblggRi5w0JvmRz3Q/NqVoGuts4VUxxk9PbTiO2g2PTE6XSx152iPY
6lVOqPdgrkMMMV3oiHvYgJjv7QngU++OEjZ/kQsuy97dEuyvj8rAaIcg3A+oXHB3S64OXXcX4RCI
uBMTw0OkXRH+9Abi+Op/LKZPt4i8YImggP8AxSqZxS7OcLJexzCEFwcaFEahgf/bDVtsdL10MuNa
u9UN8bPtbhS1aYLh5Xu04fkzw/z3taPXgU+NRLq0sclPLHlr+OWR2vHMSDJOGFghg3x09Bd3t9x2
SiixIfvrmVBLPWeReV/BJ/TTj+jWSYNI/AxSuClNRdgVdMlZxqDIAuSZCmVo86sDRuWvTFZc2GHo
e7LtqpQdvXWZBRqFdptImLrT1ZTNCzpfAeOhmXKhJZN8s7MMv/nKZdKicYINM1mTh/rUvwXtUOnz
aVi+a1e/JnwYNLZhF7n0GA7hmF4NkmHN4IBC4vZsMb5VUo94AsDO/KrpStjK4KBSp2s+MpTAkIwO
pCAnOLpG48GYtNiVq0tZ+/CAuOA4cbx7S9uPSgo482nUj7ck4Edk4YoaZF9EPiuwk275yRVQLZml
vZOZuUxT3ilyU/pXQRC8KUcTcHuHaScOm5PZwV62JnhovFUHyqiyZuhci9lj36ljBkMS8RcLmjYF
WBY137tZs/Zd5veTkr13dV+WBMlZTxs12EieoAUFpvmvEVrGiGxSB8sEL7X5BP+raMp/+c9e5vGY
y4kV9oFXl8Bnfn/AOxA4dp4wB2xHhbGvi9xW1iyS9cUwzf/SYn1gN/vh0pp4ZPQigpDmgYJf02gZ
W/ucSADMvzaDgS0RApwLvUIZY1bjLnjhcaTu16lMLl8Bp1YhBSYWAX20+64YIlbg4wlsGAgaJRWD
0ig7o91AqKai6Awh5V0ZddWncbJqLuY1dTB/QPPOSFtX9TjE3OMH+PeRlnd/s4s/7XBp2yZOvYkT
SVOeAV2vbmiuszYL9Gxaay1ZjSrmzFCPb4go4RJvXg9LChstfg+qe+9Lnh8K7Wdukx7CogB3WDNM
gkRSjaL+ynZMnAU5MupzQZSXV6/shPIvFOTmg9cpsrTTnaVLEXojesO+kDDCCTT2vdO1tKN1UXPH
NxaHbkUldgG/Vqovm/uKzRFBmThSPahQonJlDS8p7Vkps5Il/qdsUb7aqefmiejmCk6eRcw9X0h6
OeuURqPU/gjLO9DV8IXn4BnYhVIavhQhVZxwby2NZ32TtErrZSghlppOER7kz7k79HvcMGrX7WT0
ZnblgGgYZLWbRK9Y44Fts9d605+ef2ToGaxn/fq87PwaV6FmCzJR9Cvj4JJ6oqExoE1+14HqgvaK
Ebu4lC4TxVDyOSpvzNeKGwiNKOvos91hOP0ex0YOlo1UBAJl68iLCZBOMQxOYtLmUuvoNqBmP6uI
rKJtqp9dNdEiylNh1GtQEpzR3LqVCOL8GphOwdJbaG/NpKuEWDTBNaoiLOv8skqETcWBnqXAcIpa
6zVZ4q7dzN7GKDdOpDMYB8f2boBA212dqHaqg3IrEdWGAXOGzRAM3HQI48mOh0x2AJBZnvMTJWi2
eL00cY1lVrMy+ulgqP6UGosyG8GSbeq5v0tTPxqcneqqRRMexE+7MXPuvut6b4VcbS7RR7nsfSO3
/2gvOwljfzJEoLhAsp4pYaXKC9eqgSsRZDgCKD9kAVw+S29HYs3U0weX8ktke4Cre+dbjxPEARN/
YFRHq/EEr3nsSFSL6OxUe+6Byf7JeU5c7ZFJ7+j0lroqcM8CARg5jrj5RZ+LKu31wJOpvakKON+4
s/SxScRXYKtGbvEkgB8bQzKAjABKoMPmwIKKrdcApgHK5xGIAPl/rNB21HotYJdOCARzJeHmoN6z
mS4SKwiPLV/73+WRde10tHaWRPRyRnl/6XG23voqP3dAn7k7Oq/PfALMMb502YSpY4AaYpV/ufw2
9FbMWCswkPF0QIO2XBu3cRGKS7QUQ8ARy5x/hueZLu4XbMj6OIhEDua+UoMoiGAyOCbak2Af2B4b
GpvlFwC3qIKn/2OUmplP+xJF+amGUgRzdfFKT9bvkiYczikLlFllSg+2j+LLdqqj2R4gaFKBDlR0
7sn3HgtpEXsID0su4phpN5rJ/w88jOrxMNGvJKKEMD3VfvLMKYswQhhn8tojisBHExbQpw7qoQ7z
l8eP9Gxgl/F/ymx37JmYuAofCNFApFUL9YT1/DQhKhesVSDyO5iL75GfQa45AiL4LDtkAKB479HT
gXzy0plK2lYYR0eQcISkj5BqiRy0svDKha0H5ZYR7ecOhpncXxtWHabxkPa/ye1XEhG5ijRJtRWP
7+AvkTsOj09BBqihTudVT1rrCgxIWSdDPZCT8AuwXXFFIq1wXJcL6rnUqneaHGfl/J2lzr2MxKt5
Klv3jZfQUM1AwX+JiRlfPUDe/pd4BqCt44oeUTU/g8tz7MfeYedMTNGi5RXaPENq3ZszI2QLQ2VK
WTPSrkRvZG7ZPTLBdqUiKh76Z6Ku+MNCv5VuCZ25jmXJ9/VXXDlLkyBTEmS11i6Naow6x0PbkJRs
RfWZU+Vkvisl1sOnc5zqHC8MUPHMaXe9Z9bxwffylI3i1K7MldQJtNejdi9pTdvuHXCQ1FmL8GJO
vTogwYElRP660MGlLHNvgS4nKQbZqat/zQ7AgwXjbT2ZhU3tcwExIWQ3k7RiTutsAOElWKGuxdZv
xDSRMssniRRWN+jkIYpzav15KaWD24tJ+2nTKCMR5NPbfPivfl8boan6yO0l4Oind4pqy5EBpOF/
MyzC34/zjpFil5JG9GNhKjmu8lrd1M7YVBIhB/y09WaOPFVBID8pE7tyKFAqYqvX0LvXg5SG67CB
KklFYC+PF7K8BwZ6S9g1GMmFX05BKNXYX6hKPwwS8RnS+/OtiZSOEKUp3vSAhfTtschd5SOywirE
aKqzT+W/kYPb1K9m7M8zn/341jUKzz026unNSyp1lVLKUsauq58lGih933KhTLSn4WU/EGLWcLBZ
TDl4CxXpVfwxfIpUqqGBOCuAQl+WD7dUYIxU2BlFT6pzifihLIxQ8uYvsOcfZTs27qHvsX+Uznq/
IOWmPGtRhoZcW6wyITxTOGCFfnzI6ib+F+Pxwb9xnYLHi68LmC6PhwVDm0PBTjoI9nyAGM+czPMB
rW3uSkz6XaL934+tAqpctvLa2ZVJDNy7xEJ5ERvm0rtMg+yKfZUKbW5WYqVqkw5meUkR3ZRag5K+
UjYo4WTlPGRzJxFejwflBttdEWGdYpj2Y5f3S8abUlKSPsT+YVcoMA5O9mljCEFBYLVhTfo/9wy2
8R4Zj09OYMnYkas6m9VK7JrpyNOfO3BsErMUlwkpb1QzCAJpHCzMh4rzQvnqlIKzyy73jMrXJPA8
FGDre5jxnHKGIPSr3VzSm+wKBVWfhLR5p6/eTU1SRFac5emSKGitOv6+7j5EjaidqHS9BAAVPisp
vmtpFPALByPPy+K/NNAd/oPf+to81AzakzsQ2ri3LJDHhKoI5yRQdMwgDZASOVixd7gJ9jIslSQt
eGxVvIO9xWTwFm94OSzdfVdavTvFOI8T3uJ3miUfUZW37lvReJkIQYqXIGOFWanb9SVzgSlhTM7G
Q+cipKA2ROj2qYfcK3wKNCZR9H933LC6r5p4+Dl1hmgOdXGyAgCoQypIIYosvhYX+a/Gy7ZaSfZX
qS9lEz2R4IdVxLnu8zVPHK94Afzq8zuX/qho1L+AWfr+71mNETD99ZtjgMycRkoS2Ze4CZEib+G3
isIp51am+qlZVX5Z5dJQmgg2mhoofO7h4WxlLaXJAVDtN4Cba+cnP7n6RxESzk8e8+vxd9LDTR7x
q3pOdROPMvz9DaS3q4YaSDcsSn3977At27IZc6Chc8JqgLIA3e4QU652exAH2yLL+RnSk18Ek6nx
1O50Kv3aT52X7g38golGRUtP+YuGLM6LLflSo2gwf8JjCwbzDEIzuAUtvFp/w6D3M4P9riwc8JL1
tg3IJAbrfevjJ2kqbNtD7B5HGcQDu4QOGvjZ3WN2NJ8BD5Q0S1YXZsbWfphh5gOJlqS1pJIjsOaE
i9FLHpUpd9QBvj3E5Kbi3NGZCt4meMBqqGNqYsBGrGhK5y0ynCO7XAw9JaYCsytR6FF70116u7bF
+C+pxGw37Kq79GA8FCWi2lrqeXlXwZ1RqTraRM/0bfPPqxDs9Vp66JMx56GPwUWiPcLGNN8Aj+aV
kFM3YUYjNCoWCYxTV6wvaQ2oTN2oSXgF3Zs3YQb7V2oAQdalha/K9XHqvtto39mLf5nlLoNKPjko
G6rf7jvm5BXG0gc+CIur0CxA42NZbTE002D7I4Lu2F9Qej9/NebTckMeGBG8NFuMGVTThIQFK+8W
mGObGplihBd/kuz1AtdDnGJGVRK5BlR0bLWtYKw1SmCxr+Gu6Xj7a8ElGbdHa/BnqfyCTFNJ5gm9
Wim2Cp6IHh+drqCA8PF9eXo95uX9rDE9BZRx4Q/BZH7SxFvoNnzKkiKvb//pPRHG1GYfB/dzkCEE
1QGWubtly2Z+DxukUgaF0md5XhQuDX77A+PLRVxRNW4aJ89WBbWPu0xVuvE/bR4smFzMrnxpS+IJ
RgRGio4QCAwNVICrrnUT2lBEpq9FbwWAkxN/IFCplGKccO/LEed1JKyuLXGbb+S+zYgciTMtIhxF
SFEZebamZa/svKknoudvqPJgbo+a4hPVX5L1RQdXv/fFavkVd2RsVsuOTw8biTawVlK+f8JrqOUU
9pr92uv6xD/iWnuNey4XFZDy91gPrgptavOvNbnzoFoAem9TcWX50qb547CTK9r94cCwjehn9THl
vZJ7C/5CNgHVFZoF9SMBIHIlXkEuM68VK1N6QuSfPfTIeuKcbUZQNJA0TKYMjRGQCAvCc1IAKkvg
iXosOaD/NoGf4zD8myvj1A5IgK2yWOO7e+cQCnHTXxU+01bRx8uB8aS/NaDcSivTzxFK/gRdxO/O
YehU6RB/7XDRSuAkkhZ2m+nw6HFDdJAVCrVJV0hs8t3j0zhTRktTRqdq3h0aNiKkiH+LPsk7VfVm
oe0XETfZYk2jQavAhpt25cCqZjQghgngtS+gpKvV3zJgX60Yeq3V5d4cZuFB1s68ajhZceo1Ix3E
/OPPokwjLVDI13O2G8tAQuBsMF81G3o6pAkLdGUKGiNhJH9ZuRn592LqzsEguChllXTvbUpXiSlN
I9+W4c6hdzSJbcZNGlGBT7YzTouWcYYsFaWhFJ0/eMorEiOssGmik/miNGDM9TK6o5cR0CE3SfOH
wlNlA4Bv9BUbOuvksiDPI2h0QiaZnc8gryAUZK0V4I/WmPwHCfzPTKpxH5au6ZYmx/tICVhxq8ac
TKvbZxeByTb6+Y7qgBrrA56XV6knRgPeEDbRLvfUT5iF1sn1xnn9/fAsA/cc9Ere2gcI6P3zQpur
DYl6t9LBST4NcmMqMF+DCdtcurG9II62d+OfE2GXl1tXbDZemTaGmoKv8YZtQIEQAuTsIR6UNaKH
scAiRzRs1AJUts+1LWmZS1RWLuH+EDKEToB+9QmsvRLDeDojAUW4dZ7uLZJWBDvQx5olZlAmfg0j
ppfQGLFmkBtdEzQ4Lcmp3IJV3BNAYa4efji51bp8xJ2m/nKLeuS035wEFYqP/U/oZRhrD9Zx2SnL
vfYBogTltytgo2GQWTd+alXpKjEjX5lObl+ASosgZerxlYToldLvOoYreSLblYh04xaT3szG+VAG
fmzf4V1fcgSavydCRDpAgxQJnZcsS5Z4qpXw4bx6Md4mMVLSO/41hrPk9WAcHz6YrfNVfR8Wv0lA
wM2lzOW5RmVtE50CpcZDugAVil7qy785PmYZVz6z7claGJtE/hmylwVFhJr6G07WixJE2eICG39h
rLbEEkNF/yPVxUPohweaGKnUnr4fla2RB0hSgjk7YZHFjmB6uA9AzOrloAVdOWWCTsZGXE97cZAB
f5IkO0SEcYXNGfQKr+FUPXuURDLw6l2136cmrkKjQsLj8hkiIl6IsdJbY0lEplcb92wej9/Kdmf8
W94HY2TdZ37Qqqkt3RqiEj0FN+lkybVLUhptzaJbtxTrJ05lTH6dfRbkhASCWvZa6by150mMOCKn
3bFeznhD6lxdHkHzB+JtRMaz/uFq89B4OIHjk1ABqonUMo9xyWL/HXzgTxon8QftKYs4Utr/AwLf
G9zJ/U5ksYA/K/4H5pUTXFUQHs/s7m7yxk+0WYvwXSh/7HAwy9NaKUqZ/oticn5CYHRNdR0KeJSu
/F2tMou7aXKVbkyitjcrGVSeX3RHBmRY4rcw4GiTCKlH8+0yAvdH282HklrGTFqo4+zBK76UxiRi
JQQD51Vbb4XGRklkdsuHWgiELNyUIv4PSQSZMDvHqd91Ua7TL45GWVXFZvtmRniQnh3OL9Awv4FJ
ROUo4NZYB0XwDBPdRPm0GW2KTUj1wtGU2mtECUbQpOdf90eCBtC0wBnfMRB/PgEb5E19CyEnzcZd
8gsvGj09xKcavvxBwMuXs4qdW8h8VD/jAwvtbwtzk/Tur+U2iwrNMjhLXnuPUumumSEAn8KizXu7
0hK4DzAnCFOSVzPSornS0T8yUfg119WXfr+e1CdwYYJXPKmYBCO7HMsELvfe1B/c4SmyLWBnIWoQ
uAZBTTvjw6z5Em4Ke7AF4aZMDQtpQOhbRut1HTXFSu1/ciDqT9ptx/kFUhSNDbsYpDGMeWGDxU+h
zSYIGGDrFlLs7xLnBWmdCKyWOP+H8wEAL/qKhrO2zMXDeTS7jhQUU+jTlM6Wub3YYIvH6PI+OrGb
d/XdQd/LRLOkM94Sqbs8ToK6eEhy8HBtsQPEjPFyedZRWMoakSqi0kVDl+yrrdZVW2oboQIt0+oG
PVwL8+51M66yOkMfxySJOJToYC4cuE2Fx5fDf3tcnIRMSrt7wVTsAB+1aYK/OzEWZMcSiO82jumN
IHJF1KuMnLq7CMsh27sppAjwk7aHnO6vxlwRzf2QQV1vmn8in68Pe7Esuv7NHoKTITla+t/thJPD
oGVExYFAZM7DTC+ufjVbv4520skxIGDd/B+u3OgAH8p2Iyjnc4awjeie+sIOvw9PbXaWk+aFz8J8
ZRaw9Wq1qo9m79cMOwN0amgNHyDPWsIgL4V72n5o1e/mtYGGgNdFM4H0VjPKj4SjrQhnhzJfhEmE
Ez+vqbPxygpR5ppHxcHWCpUEsMlHeydJF1RhbJc7zy9rnMsvcLlJXs1xbbXxTNcoAaK3VkIMKq6b
YYPcsWoO1QsNiKE7JW61rdiA2SGEQPxZw56i5rUjXjtSnBSawZCGbYJ5HbF3HoCljru27SWXRcLD
2MayxCTrj6yo7I9q9UulQcogaf5nfE0KO9LnsTMYNtk6SQ8iWn8vPQGlqF0teyTZC5yuhLKhnXlI
156YDiiMmuZ/aq8Pz+7dYWvBFFgpevSolIuBiXe5BewnisWfDPAQVPh2UPAgnKvJRbSZ6fzubmhG
zUH70q4kJM4Tcp4z1syQ+9sLC1uAd+bi4fVa34bw8pkahscWP1zWelFpNr7Hxc12Xf4pgQA1Od/a
PECkZYi2Y8UkzsTXgYd0dBNzFGSsP4Y+NjI+tqwzpIATooJdEYK5ptfuUSO863upkYI25nWTRcOx
1oOaVUZfoxaiLIVK1gl0dvl052gBfY2H19wlHwGGIcphEYHOcEUO9wAEf7vCQkcMBSyBHAFHjJln
eTyN21bH7VI+I0hfKbos7Kn0aJfpJZSj8HKju8uVyf2nL0nL1klqSGLYh0vF8qaJ0sOq3wq4yIoH
ZTQd9Lawmb1aIe4iFVIT4MTvXTW7+poJ1r0CHXJ1nVDJMLsezqtILR8rJF4L0nUD1RHlfGkcflrd
DqKqWYKSKMCVNaEBYrmipSKtpM0wloaB/et5OUtYa4vVCdOqAp4S8/R5RuavAw2IfdcmXZcvXxox
mzhKwrUJIMNsDZKuIZP4qUZp7Bwc9yf5PjfPFXTgHj5M0ISs3fwKYcdOeFuNb1amr4EfTYT8gqCq
qF61Bp4r54hzx1gIz4/KuKgqZLbWWl7pigH8F7OqpCVoP9g0tlUATjDBMdxiqZFsApSrCJP3F2KR
VDo4H34gTAbK0V5p4+Bu8C5sjbcS0QZy7EOlInWeACieYo1LCE+fkpJ1dUFjgqnkFs7v7TE2P4Mp
pPedaE7Uju/2U7XfL3YpTOSkYzx0BA3sM5vKeUIZP6Ss9JGgrIgZ04PCHoyocpYHSFiLGMu0/2db
zQVKGGdIqgOS283yVYBS8r7nzEwgoO/1ozcyqiiWrQT8iSXAWjYeFIO0EiN7tFHWOhCP9Ynr6j8A
c30riK2eARSAFgRlRMJyCucGkbYeYO2LHp2i5FEn6WNCT1Ok9tPP2NAdPpc+t++Mmfip2+74bhh5
7DaPfh7Crj3MMEWZ2o+jRgqgBUfUxZr05z+Xgg4s3m2ycBAsW1M9hpu0RQ3zuqM+VZfkfiTmkVJ/
6tKOqqKBobBgqcjqFAhpSxjYSXk3iGTwFapzyY17r0JQrIgvDw5U2qNXS7enSKVTenfn8Xs9hVcN
luUBKRffV+HcXEpCtmtNzvl1O6f47v0/qNsU+M2ROgHSecbhFsuxYn5QR/BVMcDV564hQOnu7hgP
oGij/sIo2MS9rsNhWm3DRXZnPtiiLsW0faSMWb9lTmMPs9LO0HfIUhPa2gIuSZwU6i1MuUxlgoEK
oolCwgQUJjASJheb15MsB+0LgDWednujhVmtENTWwXj0WFqkE69fXeKbkIza9nwiTCWVWLuVVW2Q
JnbSYBuv6uuPdVl5pGTKCrgewlAkLElz2aHeI1o7Fg6uCgysfF9G+xwk+fJbab4KdeUW/j+60Lf4
6eySbUwRTQeClxdtR1+RCW1a6FleIoo07qfu9Ds0cShZyAcJm7t2FNaMAC/yE/SiFHfpiNuBnmLt
7nAF6dhR+YWh8WJKRX4vltmQCSTRZX2F9wepMb7Nu76h/mgyEfx33tTRJl4K/ewRQLUoQhUkiFJH
toJByH5VRyV4PUswT2ICtCAx4GBI+sJLyFAkcx2VZutNGOVGDHwdRcgNu+cWKJ5U660UDzGQoFnk
DWtmBwvECZklJQi6BFXZLEWO7XcnN4LGKYpj20kXLOAA/Y81Giu9IJKkTn1qzV5d0mEKP42uQJk3
ITTdqQaZECg0GIsBZ+/MGd6Wsro8zfwpk1Ynr+P0WxKzfVu+eTy77zZq8Od0O3JbBhl3ntfJSWP+
Ev27jr66DxwECW2vXPJ4Zx6ixSX0fhyevlvrUziY775rkP34/hv4P7v1774UEDR/KcGcH4+tXq1K
BJz86oiFkV9tE1EQOuAuN7cApnkZ+olw14FHFO7W6uqxFyL0g6k7wy2/p+Na+ubrteBiFX74eziz
6pSk8/AKgpCRQV/yQ6NoF6HYPnsqQsB69dIAMdTRRtbEoItgoXK35eGhKGcAhTwFIfdyGorh8Kas
M5JnaNKBt+3o1L8A8ipnU5DkFmd4fZPVZZPEbJU0ZYTtGG80TUJgJeCPPrV6RAXDs+AFtLthDT67
IVlxff8yojG93XDNr9Cn3pgf+MjptzpPbsk9TrlzCZTJxQpxnLa3gxbnXExT4BX/1f7myIHGB0Vx
2DcHlhq8KGCSNLBry22KrDAIbXKfeaksaa509VHbOoffflANEym68PEgHtPXJeW6IFTzHsYrV7hn
ugtyzXxXx0/IA+5ArxkdsrzaMkh5SCombrCdDQ1zAyZf/2X7AKvrcAV8um6hbkb1X8WLdkBqSo/w
F971O7DAoaur7PwwRb4XY+8O9gAMPNi+EH9ubcKxJtNWYb7EtsCdsJ/HUjH6ZxZzF5emV1rtbrHN
TSiPtTfqytSFQ0LWcEL/94fguIoFW06o2peMCNyP93TKlEPj730w4zZvDZpQvQrSi9QYMPLghAlX
v7kl8RLJJ1EMMdI3aCWoYeyrh9WhqFOR9OTkD++njeeB8673ahkYjBTfYMoEQIDRZm4dpGYcDNNW
iOJEqfwzoNr7nc8yuKjObcP+iiPfntHrq6nslI4G0Z4H/6Zg+aHVaXA6e78wx8npoqYqeRTpKGWu
6vbQctf4JtDQVxgbhe3x0yeivo3kDgjOtb2r3t3bYK9DHoTodAwVDRXd9W9mufjFMTCa6u4gLWZ9
6G0bm0wIRs8GycrEar7AMHyI6PPoyBjVKB3bjMjzW1J6T1I4brqLZAQDBqUBdQ0hKqDtI/GLiWnR
LhWr/RzanVy33s1MR/6/7ZJI3YjIA+AvJ9UhV4DuTQtn5gx9xEAmUgRTjTYuetuV0v1GoB17JQGm
941w/JTAZJxDLjYwBzMz2ySyjENwHEgAq57AV79vXhacG+LZuxqfzLionjYXVNLySyIod1Lrw0xL
9QjgNHtCLgKeKVqmn9mS/7UlaZRprD0FGiTAdV0trAN4hraDCHzLnU+hNoVk0AdifdlM0ZLmdaHf
UcOugZLof9I6i8ts1kRTdDiiM6iYWE+pVazOhPAwLk+4ZfPjlM3VaRi4yRaeUTzxNZeMf5YnfpOR
rf+tW/fpWkLnkPwlqNkrDof9IXlFzbodnQf4R57OOwKAVnN/3B3reGgCxuHH4Xh24w8+fvGSPT71
5W9mm00h7lMaJCCbAe9KK7zRx3bdAVU3Sc6U7t15j3kdpk938wZlEXxJRdJogt5yb9B+am+gGeCc
+ATLK7baUTyve4eaX2W/6eDIhhFMHr9IP/pRRj9tdgrxsO5ENMeo6duSmIoKj6jXUknsp29mfozu
O3zU3QIWhbhrqpXwgv1yCke0fvzBDEeBnWMhJUu46btY7S6+bcWWRj9bYwrRiBbC8kpB1b3UHcfq
WQlcskpZGuD9L3BeDBPrQDED7G2HV6VMpoGEQ2A7idLlmo6aeiAkBW/b3nr542n/w4EEW/fBFadS
6t6aFbn6fmB5chT21lAx9bKFO5PnVS6vLgtmzcu98mSp+Pue2Klfu4s76UKAXF6ert8tmtlWJ/Gi
rVZWU0+trOK6IGoRydwjM7MahJv6pH+MM/CTfsm+fq7MKwEZ/b7iusmFFYUW/A7BblwlxKdjkRKy
K8XK3e/RGlTkvKlrCU4hMMLJIOA46jxx77wNndi1ENxQdxG5PBA+DWPpMKi4xSoG+AX8GQdmebrd
A4V8Lmsr5A+sz6QBtTciSWXpceWNMStLW3WcUwu1lGIj8hTcyI11SpS40Qx08MJokb1Vv11nBe5i
HsA0Gj+m6/N2rkeFfYopDpB31WvUASDs0K2I6SnG2dl5yNz2x7Bck5c0G0aUyTrSsHoOICwn1oeS
tYd3vMEZjrBTtYF+BtLgLPDMD5euG5ANgiqjO4drav/lL9kvwcrVk13vddsQuUUOuVNNf9w6bt8v
LEAGpX/GqrYTbNzNafWHmTkYema+Xh5gYfQT4UIkAEdi0dGkxg8k3cQDuiXBPAAsQiVcABCddg75
eUxjRNdM0eI1Rn5RyEdY2RHxlIhgibKLuvMBygGO6Y2W7usosAycITZtZVPsamJkzkDRaZXs6WRv
C9GWD1VJe2WlKGdqRsUB6o0QhW3oF47YWQndJl63zWxXaRv0KWuPqQQixmSdUrborVM0U7WukEWn
5XbfHAPJlsFUP4GZwaEt7QekOQEBdRcuFL6NfgWZq5dsNjBCE+26ySdmrnt8wool87b92/ziOVi+
Cvu/jh3G0NUkrndYwUNwjGyuYN8xw9iYDYy/+XbnRDqbpL5yYlxSANiTial8Hok7+KlZTr89t6dk
jY2hpNcQUcCr9eaqaKSkDYqkb8M32mDLyHUsAAmyNdwlCWrexEkmhv5zFhF0svHZJu56+evkwfMA
UuX4B9ptcaopZnVC9Flx4fXGDR9D1gPN91TpGLEc/lmuVwuCZBikefM2in+dnkbUFqLmATVr0hvB
4Zjjf1sVLWFpd7qARbjiR3I3ZKTxOKqwKz8cODY5sgfpS1ZrCOUpShr/EpbZstZGnpaX7iCGNWq9
RRU+KeDHy1Net8U0Z7FN1ZnMtkUnn1y6KdNLNZadrn8fXHITRHp2MHbvW69YrbPAbbhLHlC1I3tc
gDMZdwxn46FSCjcf/Pelqhdi/71TDX/oyu34V6vJ0yGaUymk9ac0wnnmol6d9AEJDpwbHM3LA2ld
VYkaqIaOWNFJgGcAuyhDYlfBgKaL4gL/6eqe3JweWFYPvBx86CIqjY2h5KNzbMoyZBRfFn5ifEqx
y0ahD4Erm7zyGrAV4TCq3sEbYFmy7XLkCVVmu1N+NoL7EF6h8M3XNEOLOM9FrcmJZe/hArJkzK8B
42AugqV9aGfWgMnMe7Sfhww1NPs4DNmSJuOOTMMIhi89BTuZ8Q0W5Mv3HqmRRK0sF3rPamACY9KJ
pL9c5ZUAfqDpuHZGr0j2lgf8lmaA31hYKtmPRbLpe0PQAQCyPvHH/GkAseUzmY0DTsMdc0EN2WIH
wj3KL91Q6i5fr6U759ZZDZK7YSgweQ1VWPwQyFDzIij2CTP+qgUHEqe1l2U7sFVhdKgN3FKJv7T0
SUvW6K3w0BX24n8om+IJwl5mQy6Zei4OPL62iybH8e+WOM1OYXULhTM3Gzm0oJcjPzfizGUg6Gy4
+zfVwzUhjahRZuXtVazWtC3ukrnpXj136AvFbftSxi/gmQRHQna3YaFIsbmIA9fi+k+JyDof0tv6
UlfdpAc/IMeGNQfykQIK2SApwHJ8oQyQwXEaNbWJbiGcf5GQYjY8s1XYm7Z8OUpoduP01DUzWlT3
TpA+ldsJn1iq8YHQRJxENoaq6hG0/St6OnBdv7fLqyq9/T6JKtJmyW9ML/ZqWT2Q52jebCLP4SZL
ZxR8nwSRnUTwUfAMY7V/RbilBozzLwYZgHkSVtnMbK1cvvL3+hc4RZHffIUPJhJtRtvYUiCSaqIC
Rg9NvMYahI6TN2Ze0qI7Yi1/p2w/X6yw0dm5hC2IvQX2HxUZ2kUWQsmMAJTRTCzhh+BelQtVJ3+C
9NqFGU2nJrhOcYzZwhi1v7HxbYaNtPZXPO3/VW/vrOJKw3+gpOMFwiYRG/kkwqa2psdZ7U1wUl+7
QJwgsD10mG1kAjAgPqKkPc+bxbRAtHR+ATduWRNs7JA5ZDR2yFivW24TIoD3HxVkt5eBrd05aquF
ZI+5+PHhBjmijZ6up7V5PWIatdi0xv46qQ3mzA8tq6jXQnJDj3pfW7ocvh9pPZQYypp1ZOGfInBk
ByhQYDKYNRKLtU5O242Ak7a4OHfHSQnX5XSVNMZLgfswShD0HWGKF/fFlpYq4F15LNaUJZYxUAfr
Xw+VDJaVEBjjONnnEhMzlIivyg+E3l69j91B0kcJwZG9HPX8YKxpe8Z3w0lfoTyszkJv1kKzUPqy
2ySf795EJ6mk6UP1EfNFPHHIv06GN0qapHoMy37AIkPXuOMERGJ/TIGURpu9h1GeEIC0rPZcwser
JbRI9aDOl0sfIyEDb3PUZciZ8eiIDN3InRFHP/sV54R8zhKtSTJms3E8gLKbz2ygSKdobXjq++HZ
ThfBSXneZoLVp/RztsN3g2KNclFO17yXwMPF2VhU1vKUS7t+VjewlLUAALK5QyPm3A0QAer0pH1u
d/9CpW2p8+6V4xc5F6X/t0++EnPxUW7BSwuhpjGbT67JjtP4WxBPwE9HVxaNMyCI/pXVa9p9i/jh
uaVcyGVZs/fd+1bkQJvMd07M0ynTXUu6b0PXmRZ1CzVQ8Vg5KfWgQubBvIKOiynumrvGP94pRP2f
Zy/9L8zov7spTn1uJtelXU8XhSly9oVIpBcy4TNseKenhQ/+dGfqodsdqPXXwcpnFO0vnkHWFHVx
tpRT3FHHShDi5GslkrUqnrdd7bNUDTKb3HK0CkBTqz3QAcggX+ML0pwdDg9bD4BZwBAeQeQhNZ4p
HbyP0yjAe/9+jXHQRmCWeIJit8KUDtpfzFZd+a7PUqXsxmcegcqIM9rvjMOFXR6dqwJFrI0LEEtp
vbUeAkFYysIWqK332OSZB8Zah/5Oh1GEFcQA0uOwi0JUdigFo9QDqwPd+yxutwVySrRIPFAF8YDC
CDvFvm2FvQBOC3kEZ4/vOh4Ow5woKC68r3azfblKk5H5M2xCtcFdp+XsXPKUQrcMi4ni8VKQByBi
3vYghi4jRzK9cetHV7qHVXw3oVDFHnfbY3tNw8lJCFBXSmcoJoXK/DX8+FvKncsWcDnEJuTzvVqQ
ZOWM842r6vdMGjkzZCyLXbipgzTlNJYl3LdSMbSuRfmGoUmhrG/hlRcCgvF/6xpmIJqpXb7wEGLH
QJYsGNf3ylKIzRjitWmma4X589XrKql37pADcwN0RD2/L3GpmBQLzdDTpfIDk86wMKtlmtp0OdeE
lycqTcOhhd7BF3c1i+TlAs1n9rPosB7Q0e8oCVc+8Zix6IuF6vAuyfKiInvzhUmbEtVYatFHj3Po
1a1ImTBKrs/ryiYWbPPSvM+IoWYWY/MzzWWeAuxXcjV+pRRV7zWZT5wBBLMnCBw5wc2fUe2PGswO
YTDFQ6bjLVkwEnPk0d9XAEMhtbyFLLoK+SVaFGiHLBOD5BIHxBmD3Mlr3a+aWn17EtNfnqhwRyPw
JiBtkZBDoiFSzsPn3tkpAMapBIpS+OISXLEwH7d/YyPiEyZ05dTfKA0L0moEoi8ILUhUJJkeTric
dV4FxHJm5iHu8EouGk8Iz12NdfZm0kO8WGWB5kqq3y5nYUqP8ELlXzQtT7NXcxqDsWeJj3ZRyJr9
UgMHaInl8iB9AF3sdBfM6VQfbB9MGn0hZslrwqVuLFkn70mMaQf1oS/qDMJKvplhZr5D+fExOYWj
bvvTiLxQy5oIG3W00DVpZ649X4+71jblU484FOxvyPKQmWO6ux0dHMFjGUH4Ud+8Cdhe3ybDqgbS
2bVwsr9yLbliPxRBrdqHGqYvZl57Spwmtc2GqzroFkxEY+VZvRcFFLgYNaTOJNxxjNMrNIC9VkcY
k/1I5ikloSosbX/3ljMDxwYaVcChALMlqb54kiVpxlsJCCYmU4+LoxqPlah32/xSK9hr95ZwojBW
auc7vz/y8z7KRbhcUkyhqxy3GUX2fzXOJhJwZOJColm5bsjd2qR49RO2TBXK38SKYjOaCfk/8Jkr
ejOLcGU5igjmQOTdHoVnrV8AFaDCwm6nVZ4xzIm5EpKgFzEv8xYZrCoybAIODYnMLEmVpakzdLqn
7B4vkX4al4rodspm+egpfq4+t2OQ8myfdEjDBw8Xr1zyZ8xSPmgyGixSBRkeyEHBI9BGyZ8iKnUP
DB0SeJYLXcqreLUwu3l3kQHhZBg/hgvEvCbg44JmVd4VWfFL6iIE2M2k1lsBk4m5J+sY6fn9fz6M
p2l+WbtDm545fBsNLrVfh/ngitFbwRkFgqbG4lKoFR6GiUBMmExPIIl2vp2iXqeRqpltuQ8Kkvrc
XVHp/c+6AABoZ65QzlTiy27xw+QFESE45fMcl7KRn+Vsx1GbwmKJQtw0cGZyuOjzdwH7I4fd1IpM
eC7h0q96nlV73As4pWKqAAnLmcyrDY/hfiXIhxxcZtMIjfwbCL19ADUYkcMyMQW2+eEAiT4XRixk
Qf3I8maRua5YHl4YlCU1JmYf28HWXwfre7A1KLnEhnEQqaJ0dCo3wh6BsqcHqnliLo0y+oXpYbVp
mFYtngCip2qNJtV8/a2xeB0bg1P0J61MBks3u4IpXQN6WcsNperI7mt+9/AvnHyrxeySU9Gz8nU6
7mVTh79zDAoR6aOzbgQuWrvWr99bNdWQphHHY8aciDtgg9w9QmwTYwBqJAJBkmeB1EOE11RsFW1H
9L7uoKIjWZbbVGjB3d3IN/rJeHobzPf6WPHEJAmIWaRrPAKBW4Ry7fjsASy8Pf67bwrI5+f+T+hl
YjWLRVn2lFKA2jbGZtZXMfw+Hnbrqk7oqwWM+ILJ5GdlBDFe7A0z1drj45PafPulV9E3H6AX3wxH
Ht/9WCVX2/wVYIkLIdQbcgNV4laScMcPKgNjOvo4WYj03JBY0NUT08PQvNYsTipcg9ts5C0hrrz6
M9IzyLk+7DaTMFuFpC7kacd1UFOH3/zrPefE74ZxW2CJdQ2BOrVJZJzEi5Q2dLbTfEtGyLEyxpF6
hWXKBXa9pPawfVven0doGoWHyRsaIYNrR36sSEOmTkV/4M0Yx3l7Q3B4JZ+cxDbKRcXRNqmpIVIi
AvI2JHlTz9/ih492d6SL8rNjaqgVuaDq3Bhg6PjRgJSreDmohB1e4Js9DFinsgiwx5GTkOSG6kYB
F4+oyo1dZeAHwVc70jj4qVTZId9Y5TV7IEAcLdHTnKHEc2byOI6QtGyaqWme6Tarra3m0cwBkA22
ztDGoRQ1j6ZyROJQPTHzKxbiYagCGVf4M4uUERdceBDz1BN2QquQGUoX6YHpUAt2nMfpH0v4o6f6
9jkTNp6c+unKelPUX5hASXZ8HL8tTsXa9bchfS5oZGuvY1qlzFvFRU3OsXqi3/6yYPq72urxnwWe
RjrWfI2s0NyMGfTMzov+EADV+GdByO6qe6ib6lyfCMCIdfS88vEjxZO17LRW6uPzpEACDBrh/qN2
Mdl32QFyraw5j6rHq2o1Mi3zDmTPuFJzPEBdevVGYaADVLzYACdrtZCHYZm95yWA0W3/ab0dZuqb
IjUjhFMUWSdNjTjtU/F3N6GMyMmu3qi6yofQ4vFiPstcXtcc0JOb9NsOkwkY/2axB9bCH1LlzegH
AqdMOqBV7AIkq3QuzpzuK2wOZS/0rVsC4DH6p0stD5Qp3txEqHTyyx3jEHyP2n5GF7oreNT7fHgy
da++h/Fn36B6mTfoK+Oxo3pABgtP9hJMmzWjrXTq8Isxphku9d4fSuNEsVlxZtf0P6J0xg607yG+
fyQ7gbgdkIIEznsgctK58eU5MuY+yaHgwPVRQGM+aDlOpopPuuwWp/LkXBoww7fA4vT8Vsi/Z0NU
gQzwBTmEWexJr/CxnQqhil9hFK+LZrp/UP5YueT2+TLAHZ1CQevbnnRDOcx+6QKmhHGCo9dHrm/6
dt7FRFjmgrDln2lROmZNXNKjyCq1H7uJuam+CRs2uQ4BCBNGVfNnFPz0GoegE3eOvwGeCk2/9vVM
c50C/iZ8hOijkyI68E2ayAfDL2i6HhOHHigcWgz2rZJZxlA02/I2EeF/NkaMIBw604bg36Nxepav
Kep5EvQ/UMfXms+r44NKjy3zvulIypeN89U4xNhvggRnJ1HDYrIu1PgMOQPQtFYUQ6+A1JARWKO/
ax6BBw1+IVGt9899IDkbSBEk+8WtpoZJwuiAliizbH0Ayz8vYvEu8LhlNTBlf3urZv2VRhFJkOOq
rNLtM1x3FPjJMZyhM28Ro7HNeacY6dmW4qCkHS5Uob38cAWSuFRRhIvB2WpmuUVTt4w6sWN4Wx7Y
I/lLqNPFgZpeib9hlQvZnsqqIuczoR345GH2BP6MWgQD4e/FKqoWCwwfKWq58Nq6/0rpZUuuQFS3
5FZaoozZ96THslPBlBUBghCHjw7ewX46ts6IhQv8zspMMC66FxunENfpHiGcrtHG4CwcibEo0NBb
jKh/qJPQLWG3j8Tl2H4n7hiFH0aeYFMyunf12406s35Mrpgu28oUhmiNuw4/ZF5d3H7R8ipxQd8b
+DVoouaQZ5HS/fGFCYuSDzH6j+QQIe6KyX7Ixpb/+/AVKJ4eNLGoooW9Cg0inDiSYEuUt4KwfIDm
yqAJuNDU+2kgB3adhkgekRAODMHpEuuGdNzIo/pwPqw48FkRNHH2s4/N1D+w+WkAJimKdA4gZ/lF
IS/6ClwBfeg4AQaBHZHYtIzisJ6lT57iUJHOO1ORdog5ouiMZzop0R1YuJTRA0ECTpV6SuzI1N47
cOWkhKd0fDH7pfMjxQJBL/XCRJIczYDvsZb2apjBlpPqmcmx4T/on1YrGd2/qtaiigSWZ9+sXog+
WDdw2u9e78pfQzllBvB56x+wK7tYvbN5xUlusMLZb9ouiGgoAsD6xWGcpx0p5YOti4WEDvMIsVtO
HH1DdVjVTkiqrCcx3MJkTjergE+BfEVyHKDNsfEiMymugHQFlTGC7jfFzpyED4Zl2cCybHgBlg5c
rJ/ZTvwgWb925YaYUeJBo56NSLkNYoVXPNIO2t/lNChIJKsAygecdlzb5V5BGvnUuPv6t/RE9k7e
63VzwbCFMHwZsWb/IhhpFUueY1WOgsehhjIlglN7NSe79lXKLq2Kha7/+4+d2s5lqoPZ0Em6LnYr
9uThB6FdbS2sAvuDD6qaBVIwDNcnLiI3BrS8wTF1bQOS6GZC0+BcEj06lzO/sTFFmJKKXeL0zEiI
sQ/GBX4uCFUVUVz1UUgKNdnngEWRJZEq+3kGMbyTy7t4Uu0UmpIoDIPxPbrV8/R7PHboaiRiXtyp
Ke906Erui0Qz0s3K/Rgwjt7vvNnhFYcmXDp5vhLUrb14yJQuNc4gpiCF6TO3+qIfOtZ8L/9oCz+I
se3vdsC0usRVk+Ga82IKP8QAbx2jxbITBA09p78sF6EON6xmPW13+5mjXoAkvSCUEcPvBdGwys5o
jXr3cCEHfOMinhiBkCQqfZlJEuAbve6yj7ZEbfz4PdDrvlCz2i0BqBhmLkUGte/U5E+C/5kVdwvg
JUVuMmq9rsYx5DW1uHLmLwKWD5PB7EEzYhNiGACNeHynyMuJbz1BpQL1B7DjXKWoc7yJETLmWu2V
NO9QEszjrL9NH1r6+yBErfOgkHHCbEYPpjgYQ2lyEVEjekQWFJUvAnFmFuMoTM2Gdet0wPW0fcA8
FaC6zf7gVmlbogLV2PwwiSbE/39kq1btech4h0on8/Tx/yufAHYzMF5ZW7FDyXH1Xg5gNQkBEmJA
ae1WuMQtRbKArkDSXh6ucH+Vd/Js9bkll6dJB63Cz/s+bvsnXHjtSLq0LTau6eHRxYM0f7XqyjMU
swNscj0KtE9RaDRlCNYcay92Cby/+5Uvpwi4KTKun53iz64z0kAqTQ264ShS2aq48u7G2wVNItyB
wJKQY6NrKT948049iR1xmR0hwUV2+mqJzmijOHmrKx+s3sjwLPmmXQQcFp8G+8IIfRRxKj9J9slq
A1UHKJcVP+QbSyAQSEWLCDBesz2FHRn5yzjkpA5rLoiz0N03aGpOMOohBVBSsJ4nHjdFgmn8cXNU
MlGbRud9aomYV0I/03DESe1eXNae+ojYgHvMvnB026IFN4dkWc2xO0DnfMbra7fx6Hf+vXmVWEYz
DNbg/DaWx0+Z/qiFeB1mFqk8iuhiNIPAMRGEeC9dgJkfuEGt1y716kGklSeyVkkUstLqylcjxUUd
slCXMVtAxn7NA/bv6CAzmLCacY6d/0T9yKB9gzBvEta0XbEndJ7peGvFGssz8ZEeMC9OwMrxTK1f
22RHMItGe0KkkMw8Ewlc/mgXa5THYznWWviMwiE1yWo3A7kbNJiv90VW8HfYsAF2I8Jtb5DkqAwW
F2dL5GVt480F6R8k7x4+ONEz0t3IKqGzs3xPUkKGt2XpsFoS6y9Wzo4plsdNLVnlbdcVhfpWENfR
OvlqxwS3QMpwV403k4Uo2NwXAYsXCGAM0mdtJGcQjzYAb9FMQhvZTwNh4fmyZPKCh4a3BrGyLdJi
SnXd1doDBej1Ckv4UmxJ2YapNETc2W5qonyX3Qc0ee8EiB2rlwuClH2/aARv9N5LQyk0y6TPvaJJ
4+G0q3UV87H6soqfBC06JN87md5sTZNdGGzmgsH48zEeAABU5N59tAp11mdqv9HWQ4DW8Wr+iVv1
k9mDoFkf8p2sWk2BSiq3r49cHbCfcx+Ot7FLZlG2IKy0dAAHIJmp42eZ0a12zmGfDzYebEwgxg2i
F9ZGfI5D3v4086VR/eUsmkaUv4waj5A6SlwfEKxiy4NXzIcEcB1n0Voa7IOvOiXBzgAlkLZjsKC1
eNtklhN2SH1bDXB06Y6+oqAhm9wLhcUMWPhkQSIq+q6/PWO97bDychmCcMOoZZpDZrTOeL4/xmoZ
/pTVHeEdv7OY/YTv4uaPo3NdDU7lEq72g8PIZJM5bHiQ2yThiCmJlAS6/V6KPsk/q+z0fPj9YviF
35uhQdi8mSzNkTpJe4Ob4fzn3sy5h9kYEaGH+lzQNpnDrRCz3BCxVBt5GLdV1SX88vE1rFXz1Ssf
gU7N5Y62+yMtR0ACqdc1lSd+MIO8c5TwMDDiBxFx3brZqFCL5Kwltt+sYPQ4dqUf5i0bDyAedYtw
BQu47PeguzFYqcii2Obtcg9eBehHfRqcvSbiicEkdVmC3lWQTZwlUFVY9po4sUsdfd/TOBMwGNMh
4wuodk1WC5V9S7yoaQfx7tQmaWYfUqcxZlHCPp+js1kZ20hvAUPLnp+CEjpYqbrzXFB3SuCTd8so
jZfRUKGF8lfbYsiYTDFHMzoHYDWEeWJ7696BMjTlmOzXo5qEQlSQ/1a7dyVW2AqWr1ovGfCwTyeR
F4rln8uesYsTp7WkYwNLUz1z2vMsBvTMr75AOAvVrcwM1Al6ty0vYcCi9EHc3kgHEFmZhBf+A5L2
obPcw/cTvIMg/cbwgOVRDI+eXt8enKmCmZWPyDLAlR9YjZE1HM4itYEfCbS9A3xxuQl/pWliTJNO
HDd74ARUZbUXuS3RnE9/HfDWiXyL2/UyBIQNV+04U+OfXS93U2VFq7sqxSYHbAj+lPc3mIFkKPhS
aikVL6XkxlfmtWy9OsSy65XUBNd93ilnw/TMbrvM9YSMWnHow/hXKKqH/kMmeFA6pxeK+lL0DkKD
QDT5xJxxIoKAwa/nhNjM6TYVbUMjKBYH0Hi9gNZWrQYWF60NPfNwip9WI0UAeAkHAcGOeXyCGV6L
vZoGrNmoi9GFWepuFYxCcgTmsPBjtCq1JfrsYlfd0anZtNycUNNoHk9Z0ckecy0JHHXA7jogs/b0
+dY7cz0UUYFJHSQffUJ+PGshLumDdKxmPFHRjNtMRiYS0VpPl6jfQkROdRh+UKeCpMZTpcwYBmHq
pSMuE++MdOhb38HfjfwznNDlkxKc5VO2s8a3Dzyl5w8MkkhGzPj29nLkRynpr1hMCeFCwQCHfrSu
L2jlhcwbocDsn3OqBx9okKQqRwmdleuTkBLkXYPLOusGIEzR7KbEkVoP4wxLBUV/P8d0iznHwMmD
BnL7zTLQ1Ukq3lkTOcOZo+v0NUcDm6C5chTagxNQOBrst7wcUjl/VVkGLfwYnB+akJz7008ckR/s
dSY6rhc9ASh4sMBSMwVW8KYJ0kWDy6VKU4mVr89E4pjzUy/fO8gz/8ThrfQVz6PUQHadFeE94MRD
SpFBtx1hb26eOR7YYP03dC2Z7rt+5MeM2U+2L8zlOqTt6KEM6Jwig1chHxchdz2PwphyOo/djzvY
Sa9FiFhEjx87jUbDBWp99mAwMAnoK/teIFr1RaGKRT2ajokudove99r5/9b1AyBKJrQGnV7/h5hC
NiXW0ew5R4FIw779KAyhL46GHdW7BnF2XjNO174snILltB2hSEsL0ceKX5dGCql30JFXY+twQf6a
/qcWJwVnLU0BZTeNgiVl6yzBnpYIwqdimrZWMmDjKUP+DLFOTTPjJmrqOXUf8qhxLrLD8apSmnIH
qrpOFgbnZwu1QVAQIiSa5fN88ykcKJsrB5xyxtGgx1MjKMtv9O74+SmKq73i63c/1SmruQj1sO/q
NUNO6BktvWflmaiamiGqA+ZOWf3Bzmadh0LeTjKgrDimiMz5PGFdVsIw74fq1JQfxr95vfXC+Qf4
nfhwmJV54ISlzv+PRY7KRkRGeqU2o9M/Kgocqf0xjlyfYhkZP/Cp9by37UbvtfAWDpxki7FahKXk
0x2y1AYevUn1y+kHiUIDT9c8M8dVjy+3CXePNma0QVIVubbVeRO8fXUoronT4J4117nuglrx6qz3
FgRn4Fdif7oASYJvI4zz5D0+E50U2nj4uENFM8eaislUW83mpKfiVNix0+336c6coVyUxSrupDTY
BGjBaC5W7O23XSAzkeP6rfq/cVLmDR2StStUeeP0NrmrS89RlofizzIkX32hzDyCLxeR6VxPkq2B
SZj2KLrfyJZLHvJEewwhIONfQMa1btSZBhgbrQJ/DDJMeHhd0WXUhAMJJiyagDmRzcarlOe6gQyA
u9zrmZ/LjUr/Mvtnse/MtJrndUVbN2MGqZCZQZPll+q9GIs4bC2aou/zMLgfVC7uEl8FKTpZ2V+w
04LprPgof5mtvWR51MlEbQyQEvgrshgTN0Kp62pbxT/goeB71kHcDyhZn6jVHRu/3umtjWvtbeHJ
RzfB6MbBrjf0Cj9OyAm252pHpS7IZwDNAf8BQ6kPHxQbCn7GS3xamrfnMTLvgRAvK/L5b9RYVsqe
W3OxmxNQpkc5XEhyGfCCPrUsqVdyGNBxX9poQ3Gcua+COQKyEn7KOo5Fw01eEtPDqGqh/33XWtNB
L9Asian7YcGvH6LG6oSyhdZA21adA5OzrxPnVfxZ2JLwX+rcvZ1BGlmJY8/s3B6nDqBfovWAzRaB
pxgubHO1ZPgm3pvRqssYVNcnG6YkvhFdPTBcqgM92O4h0EB3JtnFjDKSb6PuP+/0ijhPOkLe5jgu
glqBfDkrm4MC1Moowva6Bj5ZVloFdHDfR+AA5V7NLBb1Ap9sHv2JN00YScJ1rvMOBUkvv2FDSdnS
qSdUiJmY+1hNrugy7RmuVIC5yLz6LgBItmpmw/TmFECntQ1RaKfx0gk/5UIBVkJq38/t6keCvJHu
oG8TR/TIaav36VnHYgun1mT/ls0lO5JywIlTK1y8VgZNYPIypaPq65IIb/1Lgv+uCMaDymKxgz18
IiF52bGW7I7TfyjacDqa26VeWOIOE+rynXtGT2jSPOB+0yDXdvsqbDECP9AapyOaUNZCpWhP/KMc
iDp11smTVbXf32HEKAC+nHy6EulKigX+8OMUy+3BmoQ/dypmeIZZStwdlN8eIw70Pioi/V+Owpsj
CIMQCkjsB3SlxcpsviaXU3BQ/fp7U/lpc2bj0JW75dF0lZJC+9TfoiR/lfcm9TQMki+5aKfgNakU
xf1ondI9Dfdnfdc1hXWr2D1KxkraJlQebSISDbAQtfsCPj4HS8bQR+pizpSkm+xKwVYzUJgUn26y
nLLBQxVigQBDsR4jLU7kEuKvsRmafK35LTn35sYe8v1uCdXTgXLeCTp64+och2bHeESo7EDrE+5T
7n6ArAm7O2GLxOeYdwrS1ljUiFS75tAsbK9goHknwwLcHIjPkjo2OdZc2kIGiPKYFl/XgFUXZPff
rhA3TodcY4sRkiYWOvQi+YBlK1iYX3kj13CECauMq5UG+pZ80YwCtIaFXdsb0r1tNEE5QfFfh2c/
QqaB0l1/VW4ErGbNHmL3479FGfsB4oFQizLRZ16en1MWkV0NALg6yvvzLqH1oNFyl8wDXvqq7U4G
RMfHMzr5XEVsWx784yQjSzZl+Zz7z0Vx3u6XPYuE6sZqGujotXdCccBTkA9hvt3s2kn8vEAVEa12
7on/iOfvVitlErGLt1uqeQ/RWYDpIRL84xJKgK4CnMInQTrjfCWW2n3uSjW1Qj5peKKdDMP50MXV
Kp//qimQWXCyXQRKGvwv12lnhsks+riRJpBKRw5KsjMkf2wuqFG/KwqMf0imR8mi3dJJUb/WC6cT
DV/qnAtTPMMsngb4zLRImGIbQ6bH5B9q+hUbiD+r/uy+1eg3MLbsQzhD9Ec07+5xQZi0Ru0x8hqM
4tNyG7KPq3rX0k/R8XDJ/0VKaK/37HQcEr7illjgkGf4tlFZQ34F2fmfU8HaMqGTfa0G7kEonjtD
oJBPAGpWYmixX2Uz36ox5XWpG4N5c0xq9pyaIhzPvohbkjcGKApv1pslvGazQpEu0mhYBvWrQBYr
t5k1iCLpsc20z1uviXBpIQqgLE6mI2FuqyFXR5GMr0r5+tQZuEkZjMlpsBwcuMCDSw6MsRs1hh8Z
G+g6UErHO9Wf74vu+/uFHTA6RJlwkZlMbkBV6gV1cnjhiIizsVBS7ALLJKumzvyx09/oUqRKtPT5
56zfr67w7/oPG4I9seU/j3F9oFWdBa78oYzFh4Tg5RsYWOu1Z/QavUyi678T/6LzkXoL4LSuZTtM
B45EeAAnASSC2mKX8sFHsloZofrq7z07inTr4QSEzf6MiVkCSk0Eq01e60jWZHsOct6/Jv9berdJ
CyoajnDz9VWiBFzoxKa8ihv/Fi4lJkV3sZiAcofNLhkJU7rhMONhdNhIAM3547eQpZ32aZuq1im4
CyYwq6ilLXVOvV397uW7syvQr/YilI6FC2Muh6Z1eGNMXTmP/cdpbFwN2E9iEa2IrAkJqD+Jnc9e
0TvaIXLB+GOO0RdgjErVtfKan0GGlMV4smETBrDCzWiJZS07eLeLHajrTKT0bClFPWzvHaDX6h+/
JHqjQSKmPTZVNpj9aE+axZeOT/yt/Z1PT2o3lN8GE+LNX2WF4Wuhbm966A5ZqJwfvl87bhjnzp57
V8nsRKXAKMjhZ+I/FZD3qAy4i+41Cl1y52Nd1QWWBA0FQWFpaDm+p+PPem299zbzOGBaT1QMjvVP
Kt/1zapLSTeptkTUaToHlvrsUqCLbjks/Kggik9XQ7/0mTBLvdHZSa6oJsUV7Fn76+eJ6jjLkCU2
0k7jlyeiEcL/akgF7nsxXhmUibf4ssUyWfPClyEkb46kFlp7No8oc1cWECnbpPYoYtxveIThEOft
st2tpNBP9RWqJvj7d1aoJN9uv7Wh8o/7mn48srUOujUf/3c65/ptpnHyreAH4f9se1+xv8Z/QjEi
JT/pZoD4mrokeShT3nLpaomp9UU1kNYyXyXoK1s1m04Dx0JlogmKKNzVIaSYtZVDczjHuHR46PLe
3RRrFwvDN5CeM+ZWn5AaOfDN8PAB6GrF6qdQh7EigS5T5rm3sUPdxN/po7sDF6nz7s61ozREnoHL
M6UArcuNt7sjoRhN+TOjZ6F2Zr+FglgJXFKoy57MpEz3C0e1xliPabgYlXbDs3cnA2TkzAHCbC25
RzapR1nP9YR88GFuNCmFPCY+UQosyTDmiUEBtGkdsU0rUCS/SqPFi+g72bwqy10d2mUMHkQbDomz
LQDB7f41PaGE7zT2hLMHn2b3VIoEMrGYavgY1UAINvVjkqv3JYnArAKqD/TQGfQaC5kT2TMD+ZHO
9Dt9xGxHSmokxJhHZ8Vn++4mItAsrxI/oG7GfQZNQj9zaBGhWaOsCn+UROJgiu+BwCfB3E9Lkny5
MOyaqhsI6DPYO9lTnwQjY6I2q7t0ZwZiP7kaitcEjL2TCSCs3Dof+210yD/JtPNnBDxvHIpO2TJd
aGYgRL8ya4RA52srEGzunJliDb9k3JaCpyymLvEwypy2WHybFTcvkYCQJcP8YI9SsH5clGG5bkGn
ZSAsBIIV4qqSgmVpztZpMjud2rfRHsDCmOErbVHCgFfBEq5R6mu5uuU4slbSSWErJESZRI6Fggzh
Z64WnqVEg/4zeU1Tjx3pm5kJNvD9sl2PmpFizeCb9pSSfytk/NkYFZiAx7PkjVRSahdvF9KRjSSB
DdutYbMjWOZTlBbpZWPy+Y46nScYCqrm/c/3wiKN3Jm6bhhPqMNOD0Yn3+lZ9MzCYFSfS8nsazHe
2vVyGbSC/5fnxYMLDcXs3QqPuwFx/1qmlO8VzvEV8gsikkNXcRnLz4jtzwe2i72ZjCk+pGed7XcA
447mwwo6wdaUm3w7DPSx03p2qe7bIh6lgA4/msoGvj2bVLDLH0+GSkX2j6CJ/We+wWaV3Kjh1oh8
nIfcjUA3vvmdQPJHOzqR9bw932V76HnDnl13tEgUMHUdmgq+ZbfF/r66WJxKOGBtDIdxUruFw2ch
LOOYudtqHGRU1eOZjC12E88NGzbtzU5cbCItUIFkTqZ4bmpYcN8fMKav8nXbVkj79+W8M+2AuA15
3SlxjcRTDhbUGZKmhOh+40ElUor9H1D6bPTRPqleKCU/o/gkYsOsWYswD/CafmpOEIK+n4LkdLzy
BbkM+iPgSW0hILV7F28E2FW0M/ojLJ8BN8WlF5VmOAp8+MrSaKFCF10UmHsw/mK7ISyw/V+aKhDU
UL5OK2pG2p3YbU2ckbytso90/i5LllLOM6kYi1BcwXU5ydET23p/Vos/9/1U559ZwZUnQPeD8LTX
wZ1PYlbthswjaw+HynPixKC6e42+eAR9psvZm8TDZLHyx5q9JM4yisbUMX4wXVaQfxRhSmO+fclL
Ylx6EUcIg4wHBokMMgoqz/8M/M6E5gzg0oNBSEvIbqaqoYbCn+ikav0DHJNlJuyUEB0sryoKhOrY
woTxKbDZ8L+1qEvhU41DXmJtUP2rfbjA5c3Cnp17R5aEukAruc4p/o0usm7HRsYL+m95NHo8IJuf
76KMprzGbVgmjGQDEhw4CHcL38myskEqdKbv7/HH88jZr4zy7VpI0eJ0skZoS0EzoKEbiZzg7eUo
aPL8sDXxOnNjmKiu/w6Vu1RnVPPa1urZvTYqWsxktm8Z02mlgH1pDvQIpS9uE8lXNQ9oNnpaBqDC
l5rMN0g0RCMwy0/LihA99D+QgRybiiuVH5sVesXCzx6c3EkomDDmYbAQheV1ipp+g7k51ZHkNnKC
XgpjMSRR7LZkFgzdZQb8Nq2QT6nSXlwDGdBzPh+6Sv1ehckb5nP8Dagru/rswTHObPrWgnyJuHlS
TWa1on3iY09xr1+2Rxy00bbf698AE3cqlsvfOVje+8VFfDVgX0tyvVj6syHsalgvI1NRo4UYDK6q
5oL21kBWy9dc0on+LwNiBhqXpocKgko9pXVPGgyVWm1ZIK0GMfxH0B9nXUgBY62EMblTcr/SFIMk
QP5VooMVK/qzOa7RzQ8UFPzQw9W4yUcAURB177tvnwkc6v88SyT6Og1n1ZcYts2fq1Ph2ZJPT03f
clQa5DYw9F70eEPqZMRpqrRRtFApm8aPVpLXKO3d/To2TVhvVLPZzi2SPratXpRKhMieZA7H8VSO
igERl6B9tPGTx/F7UIH0ZzgtMAyuegpE+BJXrcij1Y+zKjZwTMKilTFaepG+qMhjkAcKM3J6cXOC
P7jcZs5BIf4DwC7gOomP2ZxW7LizhDFatg8js/+/7D+IXhbyY9fhYCU2yEpCznGgzl1SdVew7UcP
nJ5ORVF+zkvt/JcelTrO7yl+72KHC55O/Kec5dZFLDruGcgcywBktmjlHh0vLC0g33BjatKN/o5w
u3mYtxHiv7D1DMklc4ibKrDxE4/GcVyEKdnV6JMnpZeS5yuh6MduXNDpMaqR31PD9Q0HIknrMIpf
IEl86aFepSZ6HGaOc7dUrL9mgHsHT7I0cwW3+yUHkWQ/u1jJ0sxVd1LEEzUwKBs7ZYhIW8rl9gLV
CRBAyd+x4shFlXse/cRk77sJ8/e3QjZoeobkhZNJTU4shQQPi4PnnCxkayWIc4m0HndJNjSAcB7S
2anFIZGT3NuczHWmGCfhSYN3wFgdfdMDi4DSQqdXdEDdbX6WPIUnSox0QSw+XIH/fK9uOMd0CK9E
zZiZ0OoF50erKU4RERuNAMhPJJSI10YxdXmhdIYUHPXe3+LLWrwr3xGmf0KyDeCT9ySCI9xY49Z7
wb68mV5igJqx6DsQwRKpYNN6H+0wW79M4oViKdkJjJ4MgXAqK0EZTMsPDP8r7C/q4p/cEBb18QE2
jMVSaFtQaUZG/iRq00Tg/TGq+h/AdxTehkLZpEdVUNzEXT49mq6/VALd+7Gw+n4Cc8spwu0tlM9M
nIZ1cCeMcZSUIiA3H0F2DML0SJIFV3ZwZWBi0LEmJTCWLrrrFfq1s1SpIQErk8QWBRuTNoBKVPo+
lcabv/JBoEAcZOkKfE0flMHxmBjmaDnbJsc5JrfpqZW30D/osnZn+nHi+siUPAp/I3rGna8Qiriv
63BQzqr/WnDwu3hSrGiqoQhL6ZEugPaY4cv8UTXq0KNIgnONUDjUVlPGM8OeI4bhKgDUyE63ZU3S
rfTlRzLfL2pvVBh6ZkK0jLppNaSiGf6c6Hf4V7BgzWiGCcXjhT/7k4E+dfu3Sz22dVAeJKDdKkM+
xovOjOXvyqlvYwWqJxqM32HXNG3H6jqobS6ULb14f8iRmNf9l58wqJtMGzAtG1ULWuwopmzwC5iI
KF3EVTGDbMXAlL3NRl1vTfPeOLvC+at1gu39bAoUYu5T19dDVGHNjIJmi6y7bEmvfh2L7K/nStCE
weTjUAUD0ivMhYOf2sVm+1ZHuBnWDjKsZI56NgGBcOnTSW3b2C2glgnGbhF1DfRtJ34gpXFNWQIE
OJcrWNRSDIsGZGoxPyjOmkHD+1BB2qXfNW+tD7enC4u34v+cUcniByFjm2VEgJtVAy6WLVMxZdAD
6oWcAJAKS9SZhANQs7iDkWYMI9J6cyFz7WkSbAru2l2i/JadUpWCxME1ynug8vK7Qlfgc5OHOQ5X
NHHFO0TZkYH4a8oZjOfvVd98vbuYxv2fMuy9M3DGxf2AfWCWdKgCbkk1deV5YnyYvPJabCqho3xJ
BxREeXc3Vscs9YZNexiN12BQVNNBULtx6XEjm+yjxSdyN4cAs7Mu7jePG/PSLYa4uuGelwj8l1g0
qtxy8UcBW6JWdiCqU/Vd1loJRaNWn1mqvUUjGJabtFisstgY274iByaYhBvrCdO05zye50yN4fK8
W8Dxp4f/7c0zap4GiZ+yFXGOH/zQada7NWEzKkvNUIFTeUYDqEWAeRObOBRW8bwHguO5EVyTf7DN
BuIkfVsRsO287wLsCg+Foq5r4rgBCSxdCOL2igDduDpZcdHXRL6gddDeeBhD/X+S6j3m1gZ4U0x3
PyW9INYuzKc3vvYh5QxN3GvEjtGq1zj8G59If3az8XaUvp5deuP2IZVXmWKlMYA0KkDeB7GcCk/7
9JxKzQSNBgzIaH8FvVIl4G+eJDSelczOYRnojvyPD2G198We3JOQHlfGE0Xj+4xeus1oGWOn02W2
JH7SNahciMNSedl2Vy3pfdUSIIG2O+rtSf1fz9gcGSWjh8F5fgFeQcwaK2XUQMUhyooEX2wwNVZs
2x7yERhoRCyBntOu8G+pUg+FZNdjfubhyS4rUARmgItKv5C46SMyW5Bal+wFLzoTFc6TWaC8iqv1
zVnMoJLdqlRCo8N1hgWzbwae1+ieHZjIngTwmbVFnc/V3j617dFdZu93UFDY929KTfhJ5n5BrRjO
fKOAfep9m/2TxwISq6gq2iT6QIALzLNyeiXiBE5HLS6omweIIdwjDzlJZqWw2LaJR3g92TzDL0fj
5jOY3Nz3k2ocHfTX6a6eupqcU1sb55vqMEnFUPgXWc36gwpZ9bv3tgtVo/Yk3EO80zdsqb9wLnIQ
js+TA7EHmDwAyu6a/VoTjBdnqnH7sYp/sr+l5UAUC1oq/ssTmQp+gSO6V0KLwLr3MSPenmdqqOKJ
BsKdeI3a3DuVDqZ7j8SFTCSuIU4u5fjR44NlBW9kcebWm7r+h0O2Y+YAfKkL3H3txB3iKWsNoRq7
7OS9F50qyMX8FyjaNNh+xHlaZLldGhSq1Z0mIaY1GEeqpf6II7HgQPJUqrS9h0RvACuOS4B5k/h6
1APHhd+T0zqPG4adOdCPlmXoOPGr90alvxi29y1sUVrWm5LXgCErkBfHHe+hB4fh7r3DObMkMLmw
3jJ/e/Czj1GujLmIC3OHBugQ4e3GFydB1MvwlRzOOKrJT6snVKOCQpqv5/mvZzmC6mAPM4mx73Qd
aby1VHAL0BhVYKWzUpHvnNFg6OaNv4j8TxnsdXxpXjtiYuCHDxQVEYQQtl31FazfqAYC3grO6P4L
SXJUqwETzsLrI7B+HfGN6EkrAH8wYBrUPqYf7VFbhVQdzoe4O4X5I68ERO7+L5pCtWsmPXbDCxSp
51JgiYMqHoFSbcTiOITanDt/1+Lup7JT2AAoD/v5aspdG0fgdgv1N8HqynBuG52OAFmPdILOfkdO
YosSF+z4CwjvJxxNn1fztzdX0WrqZbZV63IqqX09n4hTr/azpd8MD+po3ZeAF730YyamyJgoP6fR
hkgE2owTBjDxnjgF1tyswRuzGih1P+zYCP45cr+4bfSC04sI1HLn8pJz8ixBNwMFo/0JViaUhu5V
HwjQws/Bn7kMHqyneJ680rDvldK6NHWBSg0cJltiriBTU1QiQqiKQnZzjjiL1X+nI86EIAtMGQbR
cr253cQvflfRG2uZs0ILHp8UHf8B4VRDDgjK9wmxEUXuapjV5xftyvCsVmgleFO436weBZ3Xkp2Q
pNeiNZmHWuHPT8YG9rCWIwUiweSBjk8aeE3VPBAX6d3LOTBBQEPbYh17aMAHSG7MBuLt0vfQedJ6
8HIcHuAcMLoxNyYLm+hmvcQ4q91bscFEqMVzEkXKVZLJr8vtOa+jOba27q7AbMMWAg4d7TIUBlBi
E81bYlkmgE3dxnhQvI02FoAmMdq3a5uGiPW+v7PoEKm5gdwJldkxGOMoMaleuJ0SnqyhDTeRGwaN
T2KroUXOB1+4eEiFxpt4luQ5tIpO+FJ4Emg30EN63a1L2Oz6cOzn9omqRYbR8BCYQ1rNqhe/ETNn
zYAnGOY00aLc3KTpSGqh5vgZPEi4IRwsH4/sXoQm0P+mivKa9hfRqOMmHghcU0cZVjmbY9hxqwMy
hQ/EWg2s8+oIpF/XHuCB05+UrThoymeWbfJuivFrAONhgehY8O5qcNAVze/JLMjY5kiG4JKYDvCO
99MzNgYv5h1CBNWJZi3qwm20fxeloiUId8eIDj2oZLyeyeNP5At+cEA394pxSDe66qJaQSkTmWg7
i4kkkn/5mVzP5UM1OM9eLeC0wmfqZr+RTnz31d+NaoObtQVc6Bb5wR102FT1tMrNUkP6SwrX8E9o
0abEStgZtTiALw+N1epwUQRBYq1eq6UeTplEVJTVu5jA5DzLBtEYd8ArrQC/5LspItdX48ksUEyR
CQ/IF+KL+PtGrLjK+4ILu6+vqJPzuHqSP1RP7Cf3kMM7gxNc2w17J965MkeYDDt8I68pS3ihj3YU
mwUzEPvU0Hnwq+vry4xJuYThdhNVWlwqUn42Ckq7ECXH3679BktZuBppYY2MkfQHRtlss7zyppqA
/vO8ch4tw17KL3DI4lZhQY+pr17LgykW2sgTQGYmtWid2PUHicfutOiy2DgyoNpicN3DSujjnCV5
lpJpMrBQhovL/koT2HqREVjuCdVk72p+wG+Zn30T+CyEZR5Kp8S7q1+aJU4XlpAwBhaVXJUlrqVD
B8DJnxFjcped0uOXg5G2NYO1YfrL+V5l3zG/7Pp8qaafNMoq6rfK+NUMlKJ3EtLlV26vuAALKVNJ
ZH4fVHYmPMYlpLfJCs/0v5CVWZSBpLhUfuhcNbLMdlEReIDSFjb5Pbif0UV7J7x9vxFt1OI9HqRT
PIyllYnAbrlYq/MwP8+O52wCJzrDyBlvaCcbfSf+zZBy7yH+hy27AX7ww2+UrrfvteXGyeCatf7j
jyEsOmfricRIci1bkU0vZgibgSJ3vLiSxgyf/cPAyc8UnAozzBpHlGA+7jRl2Eo6WKLky51RQWhB
CmNAZaQ/VPpnPcXk1pNVS8NnW6QXf6uy2HmF6bDjHtiTvPFKB8NUBf0Ln3L0DYJfjw+aDKkhz5cn
p2fl5kI6UHQBBxge0poRrsLuecFVHlN7TZF5stQ8t3uWguoIxwR5RK29aInLmGjN+r7VmK7N8ayp
kHziA9ExML2qRaKp/m3V3hAMAVs9b0fWY7o7vTyug9aroB9YbuN/Juea+larLiTJcRP+Bf47RnbO
8HYSEGFAqkxRnkKrKOvXQDzjo22dagnvk3dRDTOBAtskg/pj1VCJHtuJGrVmavAPcnXo4ztQ14dj
d0+rVShE19Z/85wfuU9gEQST+JTMXvCm0JU0tJSXBW9ApDVKh7Vfk1nSIjTnrAMgjqrHdRn84bTj
8eMlRwZWQoibCZcJN4GqVveZDOhRvqIvXXuiiE2Lhu9GvcXW3341HLYJtWxuMf5qKCCdzTLb+jpn
6Rh7K0pFYKRckne0/M9Xawv0t+PAM4muIs6vfHirBQSS1eVBo8KjKYn4aKGa8azlAyq0fFs+h6MX
JPgVjdiDHsHjTsU6VueMedchCtifovmxS1vdQyxcot/iX6bOT7fcu7XgcYl6sBkFm94mu0Zxl+SI
zE7aHJ5jpLFofJSe6J29+zceuW9dsf5XXupPSfTnF5AqMAjfET7oyhxTzbQ5HmmnfdIsqZeJJhuK
0QfDAz/aA8mikotMH+PoR2nAGknZdPNfZNOmzU4QL9TEnmjMlmwaZHE56fC7G5LS5t7xmJ7ZJ5XB
RNqxn3qH/umbdUiJ92ABrFDTgf2QEEja/Rx+SZqF+BD/Lyfm2OhK+aTBzwq7x1oEbTlDHPReFVlj
LAioWBlITKmDVu7K8WVZ/9edQOXqnWpDs3FRjY8rnfWg6fmRxnj8XOQFe07sDH3EQSAdTnToobmE
KNK6JUYyUTswfB7LS0rnMi5OQcIbj46WqVVth1i6ZROoU2rLY4tOYULF9I1tykHnl3OV6V7P4xpY
mDS2D3V4Dj615GIny3C1/O7pwrdYIP0E+QHCLafJsojpROTEGawXSxtawXlneRg9i3E8j69uXPxN
4Ud5wPQ8DqFmw3Y8JywWBjCYYwxVqpR+soYyjMZFM4nhQpJQDuA+QQ21wjvprJZKKLuD/K0H40mt
rWYHXqzjc0gSUfATJtM9D1nwhySCIDE8C3++OacEnCmZPGayfS6K7EiFypc7ODoM3PtLWHu+H5cN
S75aIRmrTyxhnF9mKdwB93A+I2HsTCIbZBq8v8xG4fRMyiI6At4i+fKSj2DuCFMkLjsVwoJxVROy
TP19XkB/zYFDmHtf/TIqJYXiv1ht7Y7xuvxp9ryfi2ibdrmLuhIroO97NI32YgGiyobDaA2zAjjc
wlceJeU4cEaiuDdgUq2X+teM4wac0yJtx3pSjKrw6IEthfjE7Me4elryZL0Ze5K+Ypmp8OYEjWCh
mtD6ctOYW0ZuNDbY/yPoJflWAXbfkZ5DZu3w1v7D8zQsvzZZJ2aS8QkCsm6XuSKgFVFS7/83gMhx
hKwTdKWv2GrrQMdH1bDaNfUvK26Le7XqQaNB1mQg/6bqVQOeL3PyenioQKCnUqltBOFl2onqKVCW
PWki5nq54gI/DpUj4WQO+cgBDzBk2gq0RTRX6ur1iIDQBcaryQ4JAVqaUn5hQSDLFQk80e5axDfM
X0cZCesca2FjPoNuTI7/h3Agijw32QspBWzDNuyfWND55i3uG2F3333EP2W2OTTCsH7r+WLwwHU2
sVO0eKPWeyJCDwU3kPl+ygjCPi9rchEMtkkjg4PHnrnJTpaLhbiHvqrOP2OWKBWZ5+4Xv4WO47qZ
exgCm2IRSpk2gUKyrWMEush53+wdUtwlVAxUJKYttOj/XqByMCrkm+gUAawUZ6SyssbXa/4An318
mGgk0PlsfJ2vWQ81Q4e3J5W++t/vRD+I+mbYTXfxG5dZuP3PWh0jSm8fU+5e7CfnvNUXYVw0Vbn2
kXCyQDUTKW/bKot2FrMtd1qi2n/KBucj4RlA1j8eVsapC/uWh/iAjlJREw8szeaCc27BEjmcXaiR
VIv3k+VmO9pDZ/EIr+vyGigSTfW/rSZsunaCylO8nIV4jXydTMeYRvkDfAGWhky9ejOe+7QTfuSo
3SDcFJKZfDU67mxBIxN8ZG5l4pi2ck3Gg+eV3YQH+3hB/ks7NEVlRD5w7EdDqr4//ThCw3IveORH
ttNI4+/nP+E6iGXmChC4EJorBSydzaEc8AlBLuhrtGInqzH3KH51/TKhSNppqSUEHia8ESpxgIDM
8wEHnmkEEgM70YogpqGQL0simyWhDtficuUXgDb191b56iKSmfcSvyB8voYfxekLbGDcbhvrxGjw
vT/pNu0QRkJl+iF2oGpJTeOJxAxhdn4CzCZICEpt8KaAm5s7YBdPJp/Mx8noZH1iMTDhi/seRvg6
BxLYGctx9ombwkyTTowTgqzto59k6pC2BRgrOr53bZdUf//PgjOS6Qj30oGCe/aTZRWe6lwJb6U9
vOr/Tt8w4MqemEc/rQNjDbAOKcLi4FI95Lgnk0Ko19lPNyDeZP9U5CKviOuo9NUx+JluDRtJWocX
6KnuEVP5XBRp10tGxzF4w2b6KNocb49iWSVhoyMQOYnI9eBm2XCM8sTLzSzuH4N84SfAFDtFGS10
4IFT5OULaLvYgwJQwK79c4xGSVZUbaDEI6cAruxWYo+qVqJX+p815zq77CTIJfw0SzGcOxARDuyY
/A/q8c1Spd9CcCcBL5/DhD/Hz1Dfk1Kn/z9y/dSbAC0Oc9Mmx5ujARUfyzmhN5cRnclJjlkHsHjz
jPUR5iZlapvVuR/lMZF2JxmQxWYxdkDkLqx9UTlIGGVtygPYwmrmqx39YOWTpRpZqDMQGWzt4c1i
oTuVLKsJFE5U2Sns7HtqirYq+bEA9T5hmFmFxWisYHt3p8Oem6J/yPPlcXaOzFecv7n63RZUw59Q
FyreB3dmHZ1eYyKg5iRt/XqCLJ8U4oU7NWZ/WNoCwk8CEK+SFj2CLzS5S4EILvn4VUP8MBegPwrB
0N814JPwKE01RhpfQvos9R2/tHpMS/BH6s5gCII0gLv3wC7xWI3BuFrFTWwNBa82L/e3qTNiIjLb
SsyXHt14tQMZDI5eYCY1HemsK1aUCiALQELICkGYmsHi1rm9NBo30nIfpj6Z41jJ9WwaNOsepyeo
UcKVnDzeTkh3/bQgX2AdMTaDW/JKmfclfPLpZyZ5qaLXIlyk+eUISmW2sIYMsffgV4sxLNkrNVpg
6SDcnpO3Ie5C5JVCGZxgCnkxWY+1GwGGcx4H6BCT2k4CPdTYPnn+B+dvoOdRGJhwPgiHZcZDvV3G
PPBjN6RZ/6HZU2utx26AmXvJ+eJWWkONHN+XD9cUSBYjJ2qz0h9oxo+WGQzj3sWGtsL0ZTg6qJQ2
xM9zBRHHCIzoERiTHhfvyLFqFogps8+EEPvFzA/lLIfD2OUcEU5e/Z8n7Ce9Yz7aedrioj9feFaK
YhXmVPzU4P6rLXtreQXGSTBQAVTUzEWx0v4LdyWF5F8WydAGILr3Ixa4WZn6KPrt4KUsYSsE5nov
jQbHgQtUgiU0Zw8lj7dVtazKdh8IfHuEn38MxtLcEG1K728nY2POnJcn/RB7K8PWWqi0zDPrtjvK
BiAGB56Q46OJnqik6aJ7BBcDuU06ruyBEkazElUdUBgY0bpYCLMHZ7MxlD3zLT+/7LBPN+lXr/r8
8/TD4t3kgRY5uAMqtT819EdE9/Hj/jNRugpHpmoM8Zl/X85Mk428V4hBa1xb4GmIOH2XCoS0rhnU
mvw/JbdFUFf2Vn1MLYPQS8Jsh0a/GMMfa9ZsjNNcKaF6dm+4ofMmwvny9t1Ay9dRmJlffEHMgOFX
ms/jxKu6bWEtVz4nmJHasKz3GIMFu4HRFj+tFYxBePAcjD7Gm0Q7ukDABmrC7OJobnJBWciJtZnu
qwBWPYAL3YommzdN5rNmXYuYv3edR8VpLOBfBaQPrBcgLN3RFdki/cQT3u2XRFH5HzNSZSiqUmNt
7Loibhz1OHC4K0cNp2hcAuFlqma3uERn6SC35TeZcUXlNubNWNA0y67Izi1/Ka9wfMPhfZDdGnNl
yG0ZsheukKibHKPoT9D8NmExhNlTcoiUNbJqFt1tMWG+CrEwCFjre1i9aeQpN1n9rGGwocKHYGP4
G2CKooGOdjff0zAoygHtMspqv8Zpg5fGaO4qKYfp543UZ+1Z18B9XWHdYbUSR1nlUF/T2EFCgdfd
TMZEQAwfym1/Jo1TiLtguyxFc0ZIaLVDMXOSLK6JVkfakP8chVVB8cOWMNqO2djd7QuG9O/fqMDH
8rrAm939LQ20N6o5DKbtcfsd06zfFnd6MHBRflVciABiE+27Y1VVv7SePaxNjJhgSnDR/r+4YjVU
4wO/ylNBU7p2ufIjmbLow43z/J2bwVPsAF24heIzQ120VAstJCnGCsihacGpOcrCs7O1wGyq0jAX
u5fotG3GKgOov/ayK5PGxuEirV0wg4oTIYLv1IzcZTjtovXegOW07QX+7e7RKhelP0RSFhi7czdF
ybGjEoPQ540xoth1LairVvFlEjztXYLUk0y3yDxEE0vNn5zXuni3JI/EFd7v10TLxborq0IbjJqd
N1xscYaddc4jq/ZNMyxoCRZt/D1UAJzDrx52mwxEIJKckU2vcwII0PkStyp7C16SWZ1bbgYHN5BG
dhB15yfLn9B0DV2kYPAdftwjdiaTA5MHlE6Cpg03t7t7YVcK/+JSDGHZ1LpnYBzKTxOJIDrkoIXH
FwW+0RnDTxbew55Vk4+olTGeWcMuFoqxGUxfmr5aoSX5APDKadOlhZjMi/I7QIXRU5vkG8oeaAUI
gtCRMA5pguvjQSFmDzB00iOUxQro661ZzS9KhGi1k+Apg1iArqjkCqYn8j2Ewf/RS2ZsZI9Xd4/P
iNDNFb1Sm683QG08Lg1f1n/OTTAG8KIE/6aN4Hnk75vv1tOzo9/jV4xALtJPhiUcF7nKOJWcSZtY
U3X9HSmdBsj/+GmDcg9YiocEdwmXudRqztAxe2SkgjMDatM5LeXdsHBnSihgcgS3pKCQZwfot68p
cDECCbTyozFXs9SYJjrsTfxwLE8GAnJu4cT27hr9ASE4ypfVfdwz7CL2Z153ZVeJ+NAbk0TlhJbZ
SDJhrdI4F2fAj+CPTwcVPSVDcGaehatJfvkA4uEmJ6kdQbf/J+KGWILUByDPThhFUdg++M+W3eR5
n6jCzZj3KjydAIHAUl9cgGqfBRax6r/BQszOaHIRtlg9PQV7ENgcCETuTI0e2WRUBW87kWSGWenG
xuR05GY8mFcXIb3827e4L23S+VAKVbSf1qZur4ZYkPiV3l20p0yKnYuHK8qH5FpIXL5TVfzmSjed
yu/SmjE9nbp/E9mO2j5vwi9vByc2ln+Qc9tNcFl3GCakaBQTQiQfM23g71k3tRveUTjYphhfSyZ/
CKL7q/2CHw6rk7Ibr6FdxVSkQc7RJO/7md1nYQSQrzrM/SGictTkkIEfV2nYq/alems8HVrRsicD
rZ6oLvrnsISGotUb8lLidfaTYovDVPD3Qe7umm4fom9oOvb+AHnnVgMS7QmnDreECokcl2UMYqsw
Tc0DP3S3rz4enRZmMFIyd+w3P8h9hSZ5cVoRrIEfemlvnxc/2+CqOSuGd83CY5TmiUxfHr2+zCNa
bwWW/nbTqth+5r7YfwXejW6isGEliyFQBIQWfyOsHJqGi+DSimCWQvUcrErj8D+TPmA2wt2KBH/G
jys3l9uPIxw3ozYhCM9jBtoj3ZVi6aP0K3GTcSiu7tEWXHaZgwW9Bb+53rrmDDRFZvc8ARz2zcvT
Lme6jIJ6QA0c4NUqVuU8A8kkqrRoShjyXaUPOXKIqO6RlJQ4Zvpu35/f2+s6jzIImbCX6f2SojWv
l2IEHEGXJHIL+2Qp7zY7Ax3ENyC6AGGkKWLUw7Qx43O6JQR9etLJFcocObkIFdyYwb3BpVI+zXjt
tVT4uQ8q7YU6XeEjMzlqFTI7j6yLOtvQ4MoOzHat9SwkBXgaVJxcRLTxFu4hZ407Qj/JTnhbaDPn
GSDUT7o5ZGb+NH9jtVKFAHpG7k9TO+QwVT/D8yiCEX2rOOh+tteNhPi1DeFPfN1IXiYITYBMlrPf
1SGcrc7Q0aJPMYCOrgfWPer82NlysaSfVb/KES5JPovCzKadhdlSmygPNq7Jpy7yEWuM4E72Zu84
KLvB2j+6US3jEKNQAn5DiRDMpWFTerqn9GFBkAy4EkC9WcRlL8TLPMKUZaIDyWmsNrCdBp21LYP6
0CNCUn7/vnwBD/emDc43a0nOtsBUAUWnXDzPWnYlZxo6gO3zVLJa1rYsMhUtbUF+5gMm78U94bCD
mAupiU6YaYnul6SHgpIR9YWYojofZwJ4c0vFqG5N2znC0PTmR5HYCraIkK37X6VWmuOClt7xYucg
CWdrS6A5LlPCE+EYZO6l9yCfYhyYwz45O5Ypme51AKzD8jp7knsiGoWi+4XWsBLuSszbxtOxZUmX
RFg0xUs2DjgQddVdt2Zhswl/HmXRgw5g3BpSgxr+oP7Aa8O6uCd5ENCFbz54f53WHkTd/tCyER/W
TtiYT01i85BkTFyawxsd7dqaG6/JBzK6nts3lJd/EtDSKOF9XbB2XAAoCp2g8kt1dxL7osrjbWdM
KJhTfXjekpjdojO6GqIstchjfMsvzOWvsnOlSXFdfqO0b8zOR5G3L1LoUoRmhLVbTlcX74WFNjg6
DzqDYwX4B5bzsgpCV6+pdzq85dqrUNR0Qw+dQjRGAP4Tm/iohzjuifYM0iuwD0r3zkVGHT94olgI
ZwjkOlSa1dIFeAy7PvzVecJbswfQlcIIoYC3u1nOKQmD3Jy9DbmqN1PLaV5ROFZo87Agcm3mefsq
ftdCtY4jYHlaymqS6tyaUXx2sunHsf0hgHwXS8jT29RE47wwMteqzwvjFH+8tqFdtja2TJqP01cA
c383dsxafDww3MNH3ft3WEe7LS2TLM3cp460bmpAPRM/JIzfVbNV35jW0SRiSOj3LwN6uNJgKRF0
lwBUU7HBLxo2jiWxtEOM4KWaNqUSeyLlUwV5s9uWipNLrCgUIBQhq6jNwz3GjIlyRjJ6aHvCiV+Q
9qggNnE3/MEjIBCNKCuKQLTTpFyA9lWNQzKXDrks/EdwaEcjPdziT6X7o22s+EBj9Hzl3pNVeHs8
tNX7bIazAQHOdtYTuQS2dFPwRk5PUwsJ7z3XedhGuhDG/VlWwHeXgZaZC138OiHLcr0FW+x0W1Pq
S6fga0eIDlXcrLzXI+v7EoFuDcZR9SlXocqsxf7IjKL5DV7LRM6ZDe9ufz9H7jqhvtbz+AeSwy8T
nMPoTWitRtNNSbcqlzfAEYfwk8Et8Ru3XgvvC7OTY0y9J3ZIDLFG+5fuszt66M0ts6JRWQ49XK/H
vAly60iSYEQfIbzEP7OL9/Ej8L9yM16gxY3+dZ29ghVluteZFToHObpay232fKJtIaN9Nv3HWm0g
jTibQY/xQqyksylGExwZQdxe6eB+mYtYRDHVdTZ9QElJ0uCmRiwE4JdIkP4uwt45L+JiXueBFd2h
O0Myw9jv9EKxgBdyM/B69MK5T7FpGveI6CZZ6PMu/WW1FwrWGhD7p6BS+g5t1icThost4rJwUuPv
4iCP1PYrSJ/0xoduLIqrj7NYwY1XD0DKjPpDoorvV6PHiTTHDJPfv/yquZzqBGhcIrhpzOsJt3/i
TdkV7YKJkn2SZUivlWaPu0u4F04ntRWIhSvutUnid+gRZY0m+/o1DqOuPuBUoWL00gngfLsxLWfx
OVLkImHQyReIs/zrN1JkJVzqHo663xRgaRa+nJ1RSpxFnxdHi8zclE5Y5WMRl685mfMkiY28MKn5
g7oTHTIXc6Z5QG0ZFYaK+ZjjIdF3ObmlCafSMu33tPg+8Am29WG0D94KzVV2Z2V7MzOAAPlTMQL9
vUeVRMWViFyWThfzvNS1uGQVAP0BAc21b5w9HF2yyBxlImBv/FinJFiHvey1EMA/VHVYVi2hBv2F
VHu3VeEfwO8RLyTGbTum34TfQfN/AMPt+UPoOoIPsRk1Ueztw0apL09/fnBs9cEQTG6X/rO3WOvW
FjCpX4J0TCgtxgiDaJxV1msPRhplOa+aOekxCIxgOgMKbUwoMriOYwBSYahnZgp25s98R/gEFbmq
qhm68ft4STYC8Oc8bGQFqAdNbl2hGEYAi2A9ji8gLq9lGZnY+MeR9ILDe0c0RUTSIvIGu83cf3cF
8FpZG+Z8Tet7tesu0TiADYMEn6lcX9N+ku1PmBMUjpoX2pQAfhalFEoJfYHb+ZDcHW2dpEh63ZxQ
QFCkdEKGM5erCAec+RmZHei4bb8Z1w9ooi+wn8JiCj9e0wgINxR8IFxeRctB7eN1PPinJ2IQi6ib
0gPj167OthbWFyED4PNfyGYPv7iudgCR0teHjvWDdx6FRQBkCKWjhm2FL14KANlHeyf+XLeJT6qu
ifQ3BRHwJQbgkQ7qYCLDRsqEgty8EVvgRXexJ0WwEr9qY8LK/Kww5s2IEhlWqLjSZDeHxtBaZdQv
SWFbcFUoc/pNhuavXNBdVBarNNqHGM+jQgJcnTYX7t8YDDNrO5ilta6ksSMSgPBEUP6dApZmr4hl
JlzxBZDseuEa7QwcdEBLOyJvAPXqMKtwqvwzb8h04n7+O1FwQ8hwrKVOeYhTyTNL7j8cYA5f36+W
Sc0GgvLOPlGgmmUGT9YrSupfKbJcCyOH8gmb2kp1JPBbLQKLJEDyGHaRn/cjTCw+27ua9EApNHgF
woGGPbausO1Vxx6N7RiGhaxWlHRosPO3t7ykyy71BVPmlzOpFuJBsFonS75QqJBOBOXNlY70+QPq
xsocJeW4ASxQbzpdCfhoBmhigCeSO/jV5e7NNZ+3p3EP8POcAFrcmTjv2DfGeZ9znQ5Svhv2ajM1
G8+u+9oeT2q0cu8gYyv1Lb7GtYPm253A02q8cSCcubZsLg7YkuETn0MEekeN2hJ6eYHS+ugaCp+n
03aRTCOKoSBuAupvA0Rd2N0h6Sm0Q0arLpcb8FRoh+BCioGviYKj+a5q2yL1KWQyCayDXVudD3pv
2MQGAilNhjbAwfql45GW9qUhVX1MGx+j1nN0zhRhA9w4vZzJyr0GejJDqO8sBAqZ9AxNRCMLSu3O
q9t/FfQQPK0wnrzEzsT7MywqSDF7nZ3OaTXmkAWavgAOIH0utR9y2uwgkD/09HpFh/IfpzVkFPqI
ET1rVJbyYmTyXg2Ws7xnhXi8i/RzEX0m1li/a6vfeb8RHkJNSLf1sA15A1MQ3wdyVkNayxgGdrqT
LU4AK3cjYVMajS4y83+BTH33ftICNwS4wqg/oVrO9LVO3M3jqkMtKcMHIJDlHkiFBVOUWaHI5RS2
r0K+YHa3gwXhQR51U7hhCMrpXZMfeSbVAhrmr66DlaIB/YqrgNlwXMWIkkBYfK0EIV7f/GbpjhBJ
p153w63lzHP+KcV4rmdoQJUrUAutknyWyAtLtTh4mX5W/gzYNhAj5O1EJLc7wSMlm1CWqfVzN3Wj
w2jUHiNJCSUvoRgxEc8FOLCcUt3kTsGS/eudDSzHxY2xbMdVGpkzu+eyXdxJT/ZGnexT4brrEEa9
1CGYwoG7hqLHGAfFfb8MHaAd92kWEUZFi1ia340DGn/13uFt4NnvtBlyH+OCqSlxqRPT7u4jHD5O
4mKiLXb4f/j9IR9GOGi3b2UE4zF1rBEBtoexVS0QZG/qKT2wgFlZhTWEeejJoSzVBqmhqA24+WBw
JxUpFT7amVVyl/yT6PPb5JZ05ttbDKrjMP+b1ZEKXuroF22GJtMa+kY4rKeVwfVOraECM6LHyWwG
JUoi4kBpuDVx1Xw5jSzOYskQdzwsL2/e4IEXOTp3kj/AXuRAkQTciUoBiEPtImLBpEZVWnp0yG1w
U/N3JfrDdCE6DAYAWK+hUlUB/xJF58jq1YA0yKTma6botXb3VjBcAxDpZbjeWxISllZ9Cwiz6uws
7x5G7FUmYRaMEr4tAoVLOsWweKDsevNwLxHejPGY87jeHsj00bnbztAnxBVlUYHHyUNcci64ZA0U
eG8EUQAOqRy0mbbxMZYw5IpcwbiyAV3fnSiWAYTiTiqXxjkgK7sexj2MabMQDtgDHoxy9mja4Rkn
1fgGmivrrXw955ZiqL96Mc5LMx7Bnj0rhpDINj0G0a35LXSdqY8b7sY18JaF4K79kykvXXVA3i+9
SXBEKkWoNMG6aB7GV+obKTt+PBT6UANJTFYuD4tvpIXrpQLuIKEfnniZ054dPi/IACsNuDm6s+4o
KkVSVLqtpDmIIt+fne9p6tCmpkqEyTTx7tPdGsYmjUVliKuxw5kU9g2DTVkHYve8tiFpIBJ27zY7
BoSdAupE+9jYNUeB/0oyUEyqa7IlLJA28DwmeUb96KRMqwxYG/mzQxiikswSigijy8A8gpxRlR1r
Z9lkQC3/oNP90sWIERMc7skRtnYPMo/Ili6H2XxjGlcZ4MsF4WtQ8qErBS451/Xi4qYDiJrOzGen
+VNUuKHjCM5KGxI0f54SI91UFv7QN9g3Pb/Gqh5TEX+9E3IQwawsWCkja0UNAiiUVfuCOR17uSCi
b1X0mSmxf+T9Ik7Sldj7flwmenPdG4uBHAuUTfAt7BltSjnwdI2vP6gXkGWyfG1393qeUVtlmcK5
NtC0p57ajitunR3evQ/2iimxyCZG6crPpMSY6uzHRYcnOizhEQRr+VHDnZE5X6B0gHpY92JCOXpH
UlTe2D1zVQwklENN27pdW1+tf/B4VzmLD/nGzEJwr0xQukhOYuavxDaZ6Er7G4TEISgzqLNBD1/N
ycVlivj2XmLaLzCSKymkU9Vh16LSu29eNJh1GUO5w67hxNLS1rpmwSgJ6Ou6ffb0UUKB3K4v32pf
RM+OkZKuh6Mjknx4yFn40HiJheZhraFivXN+e42svIYxUZrJcNZjxGaBfaZB8N7RW08Xf77WgFL9
mVzoBM3RKbOH3zFa/jAsSdyKLS/qH19Ec8sESJ/BR5+SuCdHEB2Q4/W72MSVjm+2Jq1KlXr5zuzr
rvWBCry7eSgU2VhAycdT5LvB0/mfCjriQHN2KIZyk67SaMoldRAHpyQVbkqT00RJwJ1cFsK/34Sy
zuA2PelGROSle3l7YbkRQsXMd0ijW2PPBA8q1OT4tA82sCQAuul1iVHVWpWiGA66d3jMAcyZ8pag
yf41P6ypjecAXdXeCpEq3n0qz05gSKu1tdATGZNmehp/J2nFj926zZOqltNcX2NanEngHw5MfOtF
ojygk+9navv9EGCwEpmzhLFGZ8LivqNXr8i4g5HcyTWMc9LEJaEU04LM2hg3EGlH4Af4MXSU/+JS
tmtjto5qMAiXKmtVgN4BgB8VWrz9hjmxge8OA7L3y2hx1qKYRzMXbc/RzW7B10e/dGy4x6cQksRk
ddbTrEBJF0PwUgacfgQ5I6SSgzft0nyBlcULSJFlfrkwlipm0A1QyKhPJg+wRzDf1nIyY8mbEjDp
h/rXOCQe4wJgd1o+gFu2+t5EZFtF5luwRL3vlBRLSy7xZZ+oOu9ypsfssr+On93Mzg9vsbx3iuHM
qkVNxUVKOCehNjY/xlq6v5QHtahQaIGEneb6mZXP9K03MdkMKuLvaTO5gSsK8+sZgzHszXxJFbBm
FUYjrSEjUwlnJWnseX1HJusrNWRJSpfKoNIJ0GpX7Sda+gj+viucHvoqYXMfKaPUmv1ekVqfrAIL
1i0j6Q+W+hq78Uw5VOdvkUHLt/MNpr7ktIa1tKLTkoASkvr7vWKmSt8VNuBKDIOzJ6nLEr/p/EXl
ByrT+kbDXUJaNxAL9y/AhyZSDgoJ5WJPRDfiwJDWDkOIMuU2b4PfIb1sIXSb/TPDhFYmNDQqFGZM
LfRaKXinIJbNgp8uo6fzlmQlUyI6GDBMDWBzL7ydAibOKwL15JoAXTQIFh6Em9PLofkcE5VuJ6Cp
Bntx1ngpc3lX/rPAuCvZatgTNJDQdgaE2LNx8mRmwRQZPuhwWWZhr+fF2UAnQBet3GBhPQA0YmNL
rQlrjS1KetxHkKPBzNhGxcvOr4MaoO8mqtd4tJJVxPIEqpWXYLk1NfBeNOoOvM4JqLUyHW4fZZKO
qwzmyPzl3NSzmCiSEQdowSk9rObNsCZSyt8D8rO4l83SQsdOi2xuHjyI4eLVS6WvwvvBQ4Y3JlyC
OuHwOiE3PZ0gd6LiqtE1UTTQo5RxJB7cFgQ3c6SDf30lMm0SZ1j1cBr7ho04MpOYUYWqIjO5RWN/
6OsN23Z5faUszbpxCvnIboihU8YvHBdzC94zb8XAurJ3wwuSnLuHRYu7V8FQsGMXfM9Y7zfYcZOV
BZgMCsKnFobWQpyYys3EAiQ5cN3lPqIb4CjMmQBy5zzvpyA7dCLQuXX5E/3BFVo02/jwPEBuoopw
3dQPFw6QYiDHPeabCwN9xWHEV06SbN98yHijQsQl4ONxpQCuIba5slcCAjQA1Vd5LOkJoER7SiOF
5pSsk9bJstSQ4js0o/ePieW7IGNXUVWDBeUNy4ZOERghhn+5C3VHqDcCn8tUhrUk0/sudb++fE/l
KlDEs/EspjjRTCVsSUTj9dN6yvWuCVuln0hQ/O95oZvWTszDLNLahIgalj5WyGjTejNuLNlGrkWb
nEda74rcrrvToNnGTV2F2iXtbe9p0CWnN4KOQ1De1966jy0EeVu45AUVqsp3MPsrejZo+xPmMcp4
iEiKw6XoxO3jqIJjcz/1nora0Y3VaVWtm00BO0XwSkreW7obUHklVKejufaOMt6qKayzr1SO0gV3
VpTZXrbqy5TFJtCLpDcR/e8tEGbqCa73wixMWdqPoxmQoZBU5IsdRce/t5/BJeNiFUlmCabNy3Ja
hrf/w2PIw0vjcu3Q6vpFVtx5ECLqeqXtvWmOeDcj9VLRpYT2HJSXrKPABjbiA4og1OtsMz4BBAXb
pXyTPl82UHD3u5QSki9JDPPhATqy6a4OEAPRBPXafZdwM0IrbIO7P4JOpk64pC7fEPvrncoAHNIW
hb6u7WBAHU5JBfIeGd/Cfjzbya79BK9GGejWxgPrKg2iGAfKjVoM3at34FXxJd7ybgxsCXgSpQZV
Zo4PonMtJ/Xwm+39OS2tZ/TF1uuzpBSOm8REx0A8FP64Ya3029RyGp+jSm7T3asD/ThzEcp8Ugm4
R/OI/gz12yK5nw+N3GyXXQ8q6X1V1ZiQsJi/RwFtDnKlwB2wBp94kSP8Ve++oYAJkl5iNo/iqRoH
OMjo31zlnshJ4teX4wWqb30XJhDH98bmwu28+EfGCpFTsr/ST2IsOssSBXDQtemGssgKpB0XVhu9
5U5wA48RC0ew24hXgP+ZvnOJxpldyiv1/rgWWaTzdHwTy0OJeNJa7euMIuteD5Ynf3jrcvn4NThM
C1o2ryYQXO2OFpPXWOkkjWyMafsYA61ojJ7VQkwiqKgbSFyzh3YnJn7Kc8G7FvieLgafAO6hSe2p
mH+medFUAdihmx+VXqPuIaiyP+M7e/5gmo7Lnt//ew2v8iU+B5T03/XnkxUFCkdzI3PiM6Pq/7ve
K2WerWUVy4oCK5lHug0kd8jOdN+SCjRt1tOgRTgytji+QA9Dk6/2c7jyZukA0dnRkydgoHc+HO6e
bJTdVCEMEfXjfuh1pNepopmo9NnZO+v+oGjqjkj+fz377Y+ss04S/JiHwYycReZZKHp8K8Fvsgt6
t+CU2B4CdSX9KNPxOIM3cfd8ArzsiUjLm4dLCaiacmKXB23QoZ/CQHQOlzTlYJNvsjNcpbAj0yQX
bipy1i6pbSeAh86TLKruyw8HD2P4bgl2xsrs+91z6VGezD9myR3ProKMKUFF5kRmPXQVgEE+hX8o
5+QEjT4hVnf9kVoult2wBD8J8XR1LTFNxP12RXjjOtMy5wZFVHgC2GZOyZQdEwLf2/oF43tAHjkg
dmN4tIhYIwSU+QnkuiV4kni2qnnu9Im68nDurzLL+C8VWcwZ4QCxsEbQsV9boR9uxAg4vdlDSYKa
Rlciwe2KYC/kxijJ4cXH66nwTgvaNQKnNtMeeGMKCRn4DYtUhJitU4fmSjDOCJEAOrDClpK4iXsy
F8bmE9h5X5rU6wN0xadKkCxnofM+ubXcuKw6uPyEhTrPvh+dkPszYV6bMepoiuvNUXjdfwIWpFXI
pOCsLOdGYn1vpXJMJG1vpaGSTqhk7OqDTs/T9xDGqdigxi7YCV7p3PwFrbNwcMA9aQakRvCZ2Gnq
MihQuPQV1TGk6dsvf4oi0M18x0rprdZmAULYnsHN0RIUptOyMtl4l90De/bQ//ATJvtgIR0st0Hp
oTEJ01AcKn6SIQ7ioQeMCaaKQLIUkY0VmMCccMs4bM8MmI4/nHzpYZFAPB55l2Mm086G9M0mFJpx
QuNYTC2ivLYVCSvKvP/xLWxVL7sRM3EK/AgLiA9VQHq2DUOpa/Or7AemaKKklkNO3j16iCXbSGBP
EIgmKyqGBj+XBf/wvzSXItcAdiH7nZ9VayPanZ+R1IWUcmmEERczRQzFp6uSQo4GQNF/4PyOXdHp
ahGW8AgxCjBCRWl9N7vYoSlToVtagowk33LPowiUwpCAYHDEppx/tpwMVjDR1ZIfjE5lULls0y+T
d85XSVJdAviJaiAXmuMjBNx6g4Ut+4KlQYG8OO8KRDcDBUUtRvXaxbgw5k8w/D6ZzyngYihWEmp0
D7/CU/J7pMKaEg3KROZ5dgdbi3SKgKNPm6+c86twk+M35KsVXUVgqj3x5vCRVunJkngXOSBBZlBb
LwTMvqURQUIelTcPNYKyHHGrIGPq58InK34dvHKH7WkQincBolGYayFg6/foIMyGBse5iCujKTio
T0bQ8aHEr+GHyocHmj38exHGkwMepo+hE/boQdcGCFNTdizHbZFxsRTSM0C2uASWNt6lY6zKbizI
XvcgKA9A8eeSSVu298/6zzA183LoST4/2XgogxOLkK9IWkALg68TsQlbF4Tw+AewFD7jO2mbKQOF
FRyHb77qKw1XCKM08Lytiv2TQ3wwN9PVH9dMzXAaTKHA1HSwVG/vQY/udiBRlOp9TZ5w/UK/GoJ4
KEHvdvmhQe+mK0q+DzV/VGpbOvF7iIJz5PIXbGB48yZWzJezZvj5RiKXjBspA3OWqVp+kXRhCGt7
fEhAgws9YTTEV2+5IkfiBvjMWI6aBdSn+GVusoh3jiQwy/jaUZPA1svMW/zigvpUPDbcOZZPX6uB
OWj8ypvrgnXfzgYXJ30kPbuefPkLqnaF1Q+GNHLsOuL6d2cKLo262mfdnmjkTFeGCN3aIsrGu9uE
C2bpS0YR79p5fSBkfF2SuomnB+xoQW+e6OdU3ndu4/O9573smHbZ3W7UM4K0Jr7h9L6TDb8ZRzv/
i3Ho9tT/NeWClT3qeWK0+YRdeCBOZhTq78SDj9ilsiW5pNN/fHQ5SkaL3G3DKpDCdC1igCi1/fHR
MICE8yxPoiHjjnwOEkb+Qhe4nXXOfm7anyiM6/cf5FiqPgcn3RHZgYX+HQ+X+ORzWI5mLx+2F//o
/s2zXLhZ8HZ3Hy9vhhzIUCa6TIJApS6ZfdFObcZ402mF12vCUNlwMlspl+fJViBRVbWt0t9bF+ZZ
bhEMpjRIItYDJ7xGK6EpjfwDe5yCxYg2YBYXeuxI+/j5DiaVRCQ7Nc6QJe7BEp+0vUH1rBdnErtL
WVHYbyaVdJsjZhDJR838hKGhEsOhFlfp4iec1Fu4tPZ5zNkjIZtXgpzogts3ZhoqZXJNP/owrp/V
PB10bV+Fr4sUh+GcJI5d4ztTzdzlEAnc1PQiVVuTp2F2LRmCxzwylyIlvgRdr0T5fCYFpkHGrkK/
caKtEtJkoRIjWkcxQq6aGlLR2DkLx94NE31ui5o1F46yTUHvW+L5rb+zs7i5TAly2Ifd1H1AxGsd
zZ6y1SPbzGFQAMjtNz2hkB79VDr6Uv6oB2pZO9gEFfEZP0Kv5o9O13+Yx+hTEXX/6vR88BISqsjW
YYhf1rhwRkZgTmQIY/ovcTiRXCLYVP9Q8a9oZqMJPa7DG3NlkAQ1V7YKcaudfC6f2zRs1Df921vy
wONsJI3gCyvKnkjlXFD8YvJwsqZhJKzkD1PE5tp2gEt3+NMGd2qjbpyQqywH3E88YE0KCVvekkGT
nEZc5lKA0LxnWSgugLtMqJcMOp39mBOxhX0ulGWlLRrc7g/9ZRRPFc+K7sPsdna/9chPcRSTFkwp
SJYxOeqsT5N2rtz/oqriPkOjeal4TrqhIurtWX3qBPsIBALna3X+SYWOhXUoRUDlvMaPGWJy8fea
2HRFV2FJR70zUNpTA5kjJpEQwzxx6xkEgpMyM55yzB1o92wnxK74LHkUWbLo40p93EIJyTNina9A
S8kYLnZuq1mkvMGBPZA0X3Dk8KLnITtnkFQcWpvfGoBJG53BW+wg58jeXcoCYrwc68Hr2j5NpYsx
Z2qaHKbv9xRtIZamfUih1heATRsO8tbGqeEwsvu1QxzwL4gdyUOcNSSC+/z6/G56SREYo/UAdAT5
4O0YhIkfbgL8Y4FnAzv99TSzk19EYbbVzE7KZtjkr5Tm+qo2Sa2sGZ0/84O3q4+PxWVCNbI3xxXQ
++Rrx4T0KaoD5ib54jO7tMLVy1z/aeQxDNp/i7+t4zysMw6d0TMWWWiRLifzzPZx1yH9+Do833Nk
arFO4rLs/pVDqTCWXP12F0iZNTBp+P6luhXClV3MOi4DoBRafqi2Gcft9H1KTaRluAKahr1qoJ8o
my1aRD3GLY5CWtV7v4LG3dtozZUMT43xjw06r5COs0+DnZ7wZhH9nL5oLW1mVgf/O6TwruEq3AjF
pXIMgO83f5o4MyQPrDYeMFzLxvyXdNfKPV5KWc7dgAKKTi2x+WE+R+y+E5v/1eeA7sWLhe/EHhDD
r1ZTFX+y14DJcfJMvVEVaML4F3Z3INOUnXI8Rpl15aczk7h9EqH2Qkp1lpoi+lL39FMBRNbPaufy
zfdYIXNIZB0/frhrmGATz65Gk9D3Ocg0/ufmS/dEMNAyolqM2oJy7AtNTuA7UufkPE+5j9Bq0MrJ
TXUA9r+89jE/3UfMkpjpgqsFT6r8jS/maGoWzdhC0CWnjYJ8Wjm6tCWLfHzletT15JdvqvPYK8IS
2Fn3eQq4ii582bT8Hx9vfOlIYU7DbzgAKjSIspi4zQryTp7q09oREhKAEi/QDW5ezrBkqAla3awR
LYlTxlEF67yO0rAhjDX9iGykPDmdR79A/32/7i3SibbJpFEiFJLfo4KC8wCY74g0j2HHx3DoLCmD
bV/deLo00kyWK+DeXYqZkgyKEkSLAfUTOkVQIlVMNrBD6sfXublHvLGvFIsWPXGvvpQ6vi9Sz7s0
o5KhNdxQVaCPoZzILmWuafEVfx5GdaP7FSJ89ls1IxotJOfXUhzxJpZ5uAPQsUwMaKeTRGFc4iP5
e4VONe0Fx53L5w/RSdLTkSCdyjmWgbsVfqrOf9IirxZKRwczIgcFwcjvOFGeTtXpv/VUwkPGvMJ/
sq+rlRyCnHD9wTn19wvEnZxr/PuNRI1o+p1507sujMHUO0utH1ImAKTZxKWLWfACYXzpEGHXlTRZ
CWj/j7plwuG0Nay8RTn4PwZrxOXb+N714bVztC71KRKk0gOxn8FiDqzHbZ1rnx1u897yyf3TVytr
Avs/HsXPLtHx98oUFTmQf102MJyH6Ms3obsxtY7xF7xst0sSpQtqbjOQfjtUNyruZh0RJkE4Usey
SYB3T13yysZWztqsJ8MMyQeFH6yqW4tjPaulvsB392q4jcGv8rBt5PfirpuXuLABG10L36jqn7UE
6KqRAgivk2/96D68MFjK+ZKE+Dly1uo+BDMnmkk4bHudku/FXEhTaiy4180EEzSaofmlIlIxbiLs
LZL3f2S/+/+jzaKJStXM9vjO/MgVvfd6ooWof3MLSLOOLImA4OQqIsFfJ8Ufeoo3w3kf16Oyao1s
H8AnM7Vvm5aNLwe4FKNpALmDwEqbh0opGmilzlvWVhW5NGJNRDmUPkxcEx4/6tGl84DeP03wHgn9
LecwYtacF6n8pt9cO4It7TNr9RCZou8pdNAoOwm+PNTfxByT//tlWw/Ev0mv/l1rCfXdwAa4U663
27aS+anu3guBODglVjRVbKe+dR1o+l8WPk1U3uRlRvUp3SCBpo/GGpVigRIUzXuzd2FuTLDMdnwB
eGdCIgLdTxGH8mDUNGZuAHTv1l0pq9H2QYGXCbZm5x09BB1IpQjwG271LMexBnp0m82w09Z65eJD
OgsulHEfm1K0rahvBsu2G8bUMFqAkR8EtGJ4V9+4C3d20QoQMTuyyCUIZ9jUsPNTFrkk9BfbriaB
XhcMJA9m0Mmthf0+jah9FicXsRCtN3EqKf978GmSpliQl03Y7i/IG+deS1U0xleNeplLczhBYKpo
AKwAUiBATwlvhJOebbVUwa4uKwGOc8lWocoAhEiKKWjBCFt9DpBDvNPyNkZDgr5ici5hwjmE7IxS
NgZlXqZO/ZUsLzZhzk4YLz4I0iWso8IyfSxnx/w2hSE9IzBuQZge32QoKODEmApi2w0zCYnYBq+L
SLOkEHs6zKEaSo1U5aGrlfc6qxlvqODwvTZxvuN4y0rVSQqntomYnGbmiCr/ja/ZxKdF/AFwmB5n
dM0FBexVumD26qTUtwVKESRw7QeVFhvuPGyGfiTmrcgwsOaHKE4RJBW0o6WzUizeXW07rlyy+olz
9rW2U5CIjqPK03Sh7UTPthrQ3ZygjQLXVOSRfpkPpXQMsd6ms0xtvJvQCOMlI8VtI8KgE8mAyH2J
Gt3iFb2kTn/RSxu+eWEVgaO/D4rb18vsmjLvaI/TjVwjEHjjimSFSR8gBg3jAEtQPfu30y0N5oAJ
y/bSCxjASXdAr2/p03JsYDf5Nc/ZeiX1skjGc1XYn7v7jDBaZQeBCYr9PAMIPh4NuGrjfHfaGl44
yE6fJoDQ5Vv/9mr4jd7XKIg3VsKUkt5G1anWXwvGAxP5byBv3H6Irb4kLz3cBmJyRie4wjzwO2dG
z0QAWyyf8oy9ABNfqLZJrjfNb33oVtXl1k3vtD/0GPzwaoEzLX7Zm7cMx8owf+aNznnGADnqHD7L
7xIGOElkbZfNnL0uPi6311eT4AHKLovEMucIlq15sDDL+K7gwmjRW5B54SJ94KHh3CQYF1pBvuQI
ZTugEEWCOKwHpXKeGtC/r1gBoLyAHQx0mMSAPvIkfIcvATqXlCqT7Wmjz2nbdu5vEPl1uVNneD1N
nn5n9k3wcPOUcVqBJmfNm09RCKhG1FIiiutc+7E/DLxqVltbno0yLPnbOC1fP5TOzBO+XlDUxrPa
eoRACagTm7GYJM9CYvbwnV2OaegzOJHoRTlzmKg7RVDcucpyDYvxRX8qEM+sw++Wz2PnoDUMDjjj
s4sBo9gsI+kQacviCDuL/Gw2UzRZ/bA/hlGmJsUh6rUuvo199jiqV4CgDl1iSexU3JH8hQoUHYi5
+KdG5JTHOG6FLxvfkLuEInezP450UddVJyYddjKD6zHlfZopuNfDEWV+935h0oWdvdIRE8udBoK9
ZNCNIz5wNC+vpmLodEJLqjyEbSLg4JQtyXCJ0ERiuMjSKcLUL0I+NwtobGtGtpNfRmt4P9iHvNKx
0wR4HLxid8ZVDwqTJ/HMdQAL08A2EPqUW/r7Qq5dHW8sMPmQaprtbQO9w2CVN9uzQvVSmD3xMS9h
YqEUUsS4/USJ5Z10oyAextm+uAWabsZncT0X2C5KwFODLosv0fArrkZArivqEDegupJ0jCPgqj4I
FIklSWSExSbutvipOYlLmS1dRlR/9xqKzps6iB4AoHGey7udo3kQH89ALgwv1yNE4I62e7UIbBad
nIOpl31JA5X33txi3Z33qPIkkZpwmrlaZX75nPPniS6/v4kOZNamVGJAdSTbvKccg31pyPxJKc1f
d9HvSXRVy7sYQeXwT0bX1yhdH7c2uIbEWqLGSdqan+YKNzjR0/L1AOGfmusqM3j/6ssltETygq9O
pbijmyB3kXh65E7eOrUQMyPkCb3bIaTf0lLji7VFH2CZ6BBiQmv6rF0CrfviTy2C1aC9sOOZoQoC
zXgh6se8j2+FBi8RDbT2QKiRbtXme9XYZGFZQHX9cFz1i+B89A9fxFE+fkTsaQv1JpZZWipor6OE
r/pwA7XsScMsJlamnRxU+Pc7eFeWKqzavjrx93fkvMtR9KCSSxp8XLOk1lRut5UEhr0E5IGXmykR
72RV6AzvIapzP6iby3Peqtjzpn0YLdMarb+Tzd27NQZV0KTyGc3uKxYRwZXsFuMwRd+CS4Xg/fyw
rTos4gszyxFc5lOXvp5hylCX6MbOELWnxoBN+V/jnXOwVTm8GWZu6V6szmIvLar2yeWORLzruHWe
CoG/UoU1mSUqwEIgWnWMzXSc0UCgG6nI8oaYpNDYi5TCvdTgxK18lURZzAhwDLIN9+xMr3r0pyAZ
aPPMigzPQJFLRACZK6rVahK/AgVCvxervCsNyXGn0h4A7RDrMKrlJ9ENcZaz7RfWY4axgWsOPn0e
Nu6lWjfgRqGKAUBntJwdTB84hHSVVcl/qh4moYDcBXbYhLBciJuajsgeaJIGcjSM5+Y7ijD7ZPFk
Z4roxpEuPxul9nd5Psi8mR0xa5mwQh+hIUy5Ma7cRiOcISI4ydVg1HGxf7oMd6N6305dC4kAp17V
3zVy0PCJE4aL1TmQlrT6RvOc1h+Hq0gHrIFtgL7TWOMnesfqOGa5XfptLbqyCuOAUNAfOGC35Cc4
FMBsTKYh3UOW+Z3RWHjsQGEZizPqb/iVUEN1dlKJOd0jqmiOWou7BtJ8pxZGRUmHSXauU73hCU5Y
lHLHWr79167kHwGX/ZptuJHmLOeNOCkc6VY8dAIbbUjKZb1XMH2FttN9nZyHFIKjrCy5ylXjkeFz
xrLbEjs/Da/k6s+wrMJqrmvomL/BLnmkz7X5L5ujv+0AZI/L0D+UY5szn2g3x2ACU94Bnc9prKFC
qZXs3aRTlkftg7KANG0bIsZ4sVv3YA87nc6R8vvn5Be2A7v6ICshhTClxI8vI2vP2/7yWAwoZoIv
F9FClQ4DylYjNIsAoXfahY1J+Y8jgi0Lz4f3rlJ7Hytj63ZZ0ZOs3z5oeCc+vkdi47iZxpHNuuLd
/7+HG8wV7T7ikNno9bekmabzoFe1NIN/vz4pidoINhli1vDXbibizSHI0C4utdjqLQNWMcKbvYDL
3cfXYz4BKj18eztT25xwuJnn8NGFsq2c1bgTcmr2uWPs5UN/guxCrbmFq7eHzUdKsDm0qFCIUPr8
nGVF/MlrmWBH9KpmO2QFDXC1N6NkX8wp4s/102DlRUYlNsIgv1K06zbhAc+xO8aDnYyzqAOqvyu7
gKEFK9qBwCXi6QukPHiI1D8SbhXZF1wlnWD1e1J49slj27JWp5U+ELwY92lQpeuKflJM3lcRPCHB
NQ17WIxr/LApQBBqPYTTB8kJ97XE4NCNCgKB792BaSfkYK5XYmiCFLMXbVMhGh2TDkRafNlkPxLP
qycwVS65JnPX01DEDtMg/f6Ui+C9MqLq1MnokwV4w8OlM8AJ31PD8HCJ7QAVoYyX15aDF5nYgOrg
YgyQIW5K/dHCUpGajDbuXYYr99/UZFNRiItH+i6WqS7d7D2Nv9zdx2q+wShsCBmq5mA5oeMZ009V
PdNKV0oGpde+4dV3dhsJEBbDzo/xC3yemIJzlahTHEcKnpuRKgP8eqnpKMiNByzDzanfRrxMwH2d
sTrj6N3UtyfCYPFjnwLhDw2ngqSeL92InEVCLczsdmxQGcnLlX64suR5TJ12PifwvX3IWdAPzouA
/vAAyQ5sepJlbtC+TXxwaNEu5+VNXTZDtdz9wwn1YRLZSNBpjFCi7zjE1AfChR/9GmoEUFCmpnbL
mC1Lxtm2C4mmeoHkyUEJKTm9zx1I6hyO+amtw3o2oFUwFUKDtIZQOJiuJno63h7RdiDzrqBgC/3G
kPMOyeBOjWdJViPSzATMtal12nXlSeasjYDck0EF6Gq+MmZjFT6r7nYZCJFAbwPZMobQvZ84BqXD
3dgYN4fFkDwa0TR5X68tq7nCk8OwWRkb9cyYW01o8nCJwh4PJN4qKiibhbICHWpp8xdl5NU0gu/k
iqRp8/U1HPu7K/9aA5lhRxDmc38weEpyWWHDG//EW/TgUFSqGuffFk8nUBz27hfg1dxhPQA0XUDG
kaQVDAYfpL/TQEpToAPJNeYaHwn8HhmCBAYd1qDBa6skwSy6P6KBDcZ/DOKJoqQOfW8S0W5p3HNi
qqiJo+Cwzp/qBZMCkYm/avLMrlQBvd6V29ciygip3J1ml1nwq+xTXBhwTtnwdtMxTo06W+bdzsLt
FMO2uLmktQm1NzlYlb+zMiQqFQIWyOlxnElCjc2wYPIO7i2a0JJVpO6u6WGsLQdC+eHoVm0KU21B
WP0eipPhJU/Bheimzci4logQtYrxfcf2671Eb0h6PDcS9X6oHds1kMJihTHVxVcjEcmDC9qfxEvO
smrHX+w317QKbELrJN5uS0uFuhtoVDt/9sJP/aC5/JsyKS1hZIszsdI4mbjr1/iJqOtQ0fNUzq4J
nfL606e0lB9AsJFOSjLkfOCcpfJ8QOpukVcyWbHM5IPjYS93OL/UuqSGNOfRaM+V+5FawY9reSVA
n4jD5TuEGgDzbpCmy47joJNnGcU084ChcG0MJlBO9SSsXrbZmILSPBowUzv3nzxMLlttgmj6kEcF
yPGH9Jkfj2/aScG+2XkxlFv8STQN4Kr+sNnBUwGtwMq7UlwuS9jplMiP8VANvKyfcf9sR7OzV+Oq
dSpdQnbVTnPHpS+ly08ocuO7pqSyZKdPCoOGHSd9wAN2p51ch92Xiw9W1iQUuth64V0GYvwuE7x4
J+faWKhphqhJdEJk7e0B83vsoTaWviV/l0BXYPKEjxxOCJb2Vrx8Mfr5pqhPWVhetOM9fyEhqUVj
5KcFwjR4TgN+sbeMlhCSHI512sLm0mZOqJELC/kYt1VVgVP5eeLt7NP8ZI2bm4RjDf0iHDY/Nem1
1AaTeZ6Qubvk85kV3EgeHo7+eINdLpTDfgjt6AbN4oveECuTUHHQ4eI8BJQg1x2vE5DnonuW90q8
/mC0vj2lotggOWSnDBgFsQ09lQKBpXmcSBTQ6zopwLpmF/YPo84OIC1LesP+o2xos7dRZKFxsnUE
kIdMIAfMG6gv/wp1wPAdN3cKR6O0khTJ9MmafSu7eKNCEaxN67dlqFmDdTFe17lESY1/ni8aIW/G
meuEioZlVmA9z5AjWymKNz57K4nrKj1/8qIbtI9HZeUcxybpXUQkTpx+sjt/NC0dbVZloauANgkH
XsgHOE9nV5NXtd9E/LcTAPvVx2w+47xTrec1b8pnA2hvRgsTMlDJjGUwdXhP8LOvzsEnTdxph70S
uTnTCruybhW7z4oIO76h55VHJlzE3NfDmR8qNxs1F0YHgSzaLWuFMpA734thA759AzmKvlKNwpKt
vRyl6/d3UzZh7AceyRlO1UUT2t/hp+QpUwYm3Eky71EH9tlkDU7Ge1xhdYEjw7dFTWuxxFp3tdOl
82dL25Y23KUY05SEawdAE9n4PAtFJeElb0jULhNtG27aPe9dhTWP3c6aoOXkBoHPEFuXO6wQecKc
x3Kd1kTQjjOqTkQrpBZOUJge2RxBpKQrTypC48lsWVd5Fw63F5cnl83Jf1dsWGPSexPBY83NgryU
KjaQRWUHlyg7a5fhIi2wiVGYmI7J99a6619TURBXmrlwh3y9AQbq5BPLCzvSARZ89Fbt8bWg5geg
LubeOD5IW1cZPM/GjkQlsd7DRRu6tZElmpch+ipN3g+lxtQZ1Y8ZAKMv9cYiFOjBHjfhrhJVHUAr
XqSDVwc4Il/2fZRuwDtwaGHZStIQwUVcZTKeI6x6rIHO3LtdBbGJ+BKu5cQNLeSiU/H5h4+FjLfi
vg1ucpzSYVTrwmHC6X3KgKfJoIY8eo4F5WzzBNvRwQDwR7xgghkxUVj+v7moWM6EGLZFipzepGsl
zzPQmc08XzDAxavLKi2DlTQMEUabR55vrHw6sexYShA5GxmgoGxLEA8q4yxy5YNR4JZ3xTOpewRs
1/9PW1AwuE8rOmde4E2i/liONmd2RMjndMSPdOjGbqtytfZmCETt7p8oXCNlOTWiwKOINw3KkfA1
nQW8WBN5IbCgAEx54HUGopawYP0QKsleZvi1zJuQRybQOIyoLVFWqaGwcLeUvLm1ZJl1lk7LXz+o
I7tb07rHuIE1BAkw1uXmqTP4+CVnLtP1/ZT8KfNlf7Iuik5VEi5ccEZ6T/zJ5b35jTagvS6eK952
CennnANrVZaIzpvDx9fLShg2/MY/hg2ya6RlejFLpiamuX4ih/HyQ1TQd3AOs3pieNRr8up8d7hN
I7R39f3DkOvKICnL6+wPqmk2dREHjPdCCOZEVdjzdA+nRr1JTVcE/JlkLCPUBW4igIFtxVqrtMbc
FBV41lDy4OPpPJ99gSC47T3wPxGglL/20sBgulgfuW3PBsdNXO3hCNmex9BEAUIAetE8EQj4v3OJ
zXXr9DupjPyifzxW43nCdJa8fedf3KWbTtWwkRg5fzQ+B+lU5FA+9gtLt5IKm5MoG4XNDzA5TW9l
zEQ7Kz6Rvch9DJSq2fR4b7d3wtPC4kCZrO9qVBvorCsCScY6zkFWZkSUVFnlwKtPfu/q8KC+SA16
niJ/E2OcW0YbxLs5s352mzttvsmslWOuYB241I2lXhlMySEUgzmqkUVqQhsRBlOziHSAX+qewm26
pOVqM6roL/Ht0PklC1M2Jw18G9d6BAhGPprFPoh0h+Z4kMG8d2j5MQs8ZXXzU5pRgc2muYIBczd6
D7EnAE5sPtZbfSl+71Ro3uxXA6JJcL1TtTozcQI3SararKyHuVx1nKqoczzUVLn1rxzFd7IoEiYF
jDthxpaXtz5fRgPkFjaorR9jFzkgJcOAs+R0Q/onDIsbO6m80B4EH5gNZ78wjgP7mi6AjzEPg/e6
mm0UlfNZeS63OWAbfRKkc8BwCSuCAWI34b9j3RkzPLs3M+Wf8l6DDLNLUXpSsjhgV9+MYbC0ulVo
PwX3hr3vjVX14SlxnwWdjzf13u0l3SZQwgMR3XKbhHvRRhp5vhLyE/S0ek6wktBTJ1GT7birNqSs
8q+L4g4wqorsVQ/dLJ7ztcGMy8zFdyLtp/9GuLfgzDcOTfQfYsMCIPb++Y5t6LsQCc7MicnoLftO
6Aj7UhhJI9yz08RTa2qUBqjxhvgHSjc9hjtFjRWMfhiqEqYz+hkpGGSvqrK+XQWxTwfmFnwZBC9Q
CktawXSqRamP/REkMW09hUGz6VkBKV4D9Dj6i9oCt/60w1hJSJf6MRknqeMtwzb16oarXe/1mC9y
Hzqb1xvj/5WlgYeOrwtX1UN0n+TtvnkFSMtvzMJxHJ2+LgI8DShpIbZC+n/A1rvNHau3NLvZACK3
Oyhske9aie4eGLNX8d2bvtBfXmBmIKufhUYA7hICed7QeYfnMWvtb8530Hzu+p4hP/1+MPI4u0Ww
ndLFBNHX7b2lUlcsLBE+ktirFgWE6lk/hyBDIFL/XROrR9U0Fti9ilV4AQ+AvBSqRNc8c6Mp/Vxn
ZBjMKmJ6OigJrl/AOHqIkltTtjPOANCOu7tD3l78/RJ/HS4Q3WC9NfOkZAtHa+HjZ0jjvZGfZlWl
ldcLxAe8nqxNubfDwhay8eP6fghWFpxyK3xMhQJBGVnlx870+cY3hXd62eu/7ujCmxpO+BC80Xwk
G13DBuQKSU80ch17uHEtgHINCEhGHdo66qAvk6soJak/q279gVDf/+mOaFiUthhNAeFzNuihSZnq
X6yUqXk89SeMwkpLuLx3SOSx/9IxRI1Otanghu+rSp0XLFlJWU6LcX+0OWz+hxLjZF8ywx6T04Z8
6QgPmk7SeBhcGjijNDLxYMrtZHpuhzVoj8qyaVk72mxDCYi/ins0AywPhZKEGDcV2TRs2KBqL3ia
LtU7DiFseEnC3Y2tcI5RVfd3kT6hKIN2wIbMHY7wa7Md8SsBpSNa2el7Zk68j/aHj8mVAjkS3Xh6
csnrPnmx8Jcq3vdz6HL0pVf2h9U7ilK4fBP0yvDoHCBEGBFNrZ+JCCn0yh1SkV3uEpC4VUivaz2x
BGivhIndkkBDnOZ2jKPgQQYa2pyV5tLQUQJ9FwgQGkCo0tFGTzGVvqhKlyYXqmOkdifcophtUT8a
LgLe0xaXUGe6GBOGi2IO05zw2aylPQ0BhOFVULzgnKaMWsBHLDtRZ3k42IhwApWGeBQlRv/Uzpzg
3hmzuESm+C0WcT7KWdp+9P0LFbatZF+ArAGS03qf3jdUjz4M5XmUzcDxWC4yR8uUNajIZ/szW1xI
/AdO1I9zZzke0qNSvWKA6NJj4tNLVJIOkJRVVfD+6HCkW7XVq752MU1oPZl25+JfBdlzjpfNtmle
CSXMB6mXuGQakWz9jByCMMeIB3AixK2U/z9Dx6h82IYQRNDNY/6tnwkm4AgWPp42F3vHI/FuBoaR
262AGJRz0gLso05h2OX6xb9cu5o1IZMTDBwHm5WupwXHs571lT6eXGEURvrxOp3VCFvqrZze6kwb
gzrYnvaYIHRNTN83+QkJExVpAn1bdnmSykgKYCK8DUxY/iF+G7qXpjYc+nnluQBB0e94aYC9NoxO
eJAdf1kmGKQE6+Z0R4vLCBvgyt62QpOdR/NuMVCtm1GUu0WfEGGZi0PBGv0+RnqjbOAqZLCHrcJi
5NENBDI742BZ/LgqlgJwhfxfigOZNWjtQO2badBw9ZynFV7l5i0MjkyR0I8zm2Maske1//XZUc7q
nDKO3xEIPmxdR6mm6hVUqZxWt8/R7NfAxUaZ3IGsqAzfjvtZORBZK5/J9Npfv3RDPj81+1Cs5yaN
gbTGxmc8o9/Pdw0nHkxrNK+ln5zgnxvfgeH+oWjatsoC9LPylREitB0g+yX/Xh8QssuERs4WD9Nv
zXCLhjICya9IoVLsm6U9EOQ0P3Ai7qjPtTHWJPz4/NETyLjdv6h9+BJwzynnlUogrLEq7SNF1csq
cvZeuPX5CdZY+d6LmpIF+r8cu2pnHKlbkL6gxrfF+NZ1OhJXRGEy3bY+bVY2ffMUi9HY8szyNh/e
rjjeK/gUS2KXloIcVPOYtu15YMf+I3eXGFpvW8FXPBAdNztfR843syUyZa6R/lRF0cVUrVVWvhAr
AoEpagmUmTo874oHOb80KJ5ormZsaK6nkbzfi4oC5q5dR1SVZBy+eG/0WL1OhVF8+wS2/YkQ1WGo
TtFoJD1L2FUqqXgAQKCH7Xj+khAC3e+/rD4sX52tH/uHlmcDT1q2Ahu+lOSIfkArRihI2Sf3LXVx
muO3SAuPqVjc0eCPIDtEzZZBhiiWNo5C4aYjSFaJBtqBDKoIQKYheprXb4A6tgI4Xz1wZ56l1EUl
HK7BWrNEUAmjlw59F2KPBI9SlSll9vl4r0Nwbmuep9GSYtGNL0BoadstUTaRxirlxKjHHmP6EVy0
fsu4UrXoDgnYfxu9GGn9Hn5ROdmwVbCmzzFafwk+RSM4Pn1gZKe/kEw5vQoecbuLJDlEB6zsx5wO
jB9aCNN6wHhrehKhvXcg07qEZstnvc0CWIphmaib2d+6Iw0EP37UcYt8kb3XuZ6TBaI0kdG+nCYl
UYQcrw2VeUUpc6A8C8iqgcIwW6CN1WUyZ3hHXSl2Gn4WV+OiyweE3Ov7KV96adyYLnKqXCMEbhxq
2MbiJIda1M7YX635qna7W4LCl5IYsUwX0YsmU594+ElfRjXhX97XXj//+H0v5lvBMNJNsI8RT3P9
Oos5VxiLygTGzShKuDJ0cP7eYJwhi4fy/vV4VOAgnW8xAhb6RmsC98ecAWjvIKowx2uKHw11/2SD
aEAQKAe5bBXjwWn1a9EKIBuccHF50ivOe7h252SUHjKOj1I6P2anodUfOGi2q0SHIDWGIsMpjxkx
YTBdR9BD9/nxvMHivkn9Q+MVNpOgMyl/TeAY6K8DP/Wp2TOAZAC67ybjA6b9kBqMoI94AqQOn3RD
wkHNX1whQDuHSb0ic2RgJbWQpUvE8RwBfkcJaRj5sO+4vuE8RJFoG6L5xvE+eU6dH/qbZbx5blod
pL2hKObSEbyXpeLUPHrtP4AE9d4WErrx9o5wxh8BhtPAgr1QC2Fs3mjVIMPfNaSL1cyjaO9rqN2T
+p/UxHnbygkjWxpmQlHoLwcRbWLW6GmXjv0YqCRW/U87RA60o7mn2sNLlDgAnR53O3mLt46i712w
8TfHWG4LPtolHLX3TNK+oriIrSe0++A0Fddd8hZk+2MFKH0vJ/aqJMkXSwFzKmjcKuwEpOMtdqtK
Jpu5eo440elCEJDLT42wYc4eM4O9Wp6P4pYsTWGJBnyLqoVFSFagGHn6aDDadpgWsqNbR9SqlJ7X
amAKpe7AHkjvvtOp65AFCBK68R4KbzfmFpUOvc1/Iqy9w1wdRHo/o/Fxw67s5X+rv2HeGQRsOOYx
AsZoy41ll2xGbB0JoRbLxmXh/9Pwgui8FNfTG6NSeG7UINbpi8nsZ/QGT5V2NBolxiU8zYreAmzC
DTs8Jw5B+BnQh9ueMMB25VKkYiEzaL79m+BPUIdMQ512T+1gZacKfQOSjnpeA++hM9fRxQ/UWyoB
neI/qZ426mcIblHZkIUysiJ0o5KFTA4omp7X82RYvJQ9lafW6x8G32wN2bOpwD599t0a5D8WndEU
nojPEKBOkzFRe9B/m0tZomNjkT+SAtP6ZxtiNSs74e970Lr8s14oU4/JjjVnuUvcYcRSxJ5vEKmq
VseFT+QFwAgxBRWq2keCRby9RNAjWc9iOSsTV5b1GUUlP1T8Mtx0bIvR0qPtblOPTW3jUqe8ipdi
/QWewuflnHBclMexvMSNzpPV4uViDKYtyFBSRp7v4RFEQO5HaqDqK7juIJpniKOh6kSHtJtK95eH
N+zoEXovR1vhLTtQtD5f+Phj7Ghp+j0AV13rdNmXgCdI6p4FQWo88dL3QY5sBA02+9rX2tQdRxww
086b4IG3Km9UKuhC/aI2lhnPdnsVa3S+zK4OAo2PTeLMeXTdqK0Da+swbF1E8aLrK3OaRc7vlpW5
FWiEfE61tBOvBoj2vpZo6f3prPQDUJZMKQvffdmeuZcdexPSHI9LMl6oMTpTaQ1XXA4PrJ+2uMVg
1EBAlFUVn7avYIdUeiSaGjUSn26ec9Q92p4xT8WFUuW3Karq0+FDY0H6RWaY+biC5l4/hJ4+n87N
ZoM9XnL+NJj9mcG4+WwZKdL+4M65gL0cxzVbcDBe1Xbx0ruXZEoJFexgn0M5OZ+c3wOe2zQpOt5Y
dx6yyGc+mNJOdV1+7awN+U7Vm4Pv2F/KkBcaEAHUyLdWYH9MFsPkl6Gtc1qtYOJjFP/+Jst7OU7e
8Or9Huf0o8FIE4MX11TaXHCpDDAg7+fyj/S8JiWAk71ZM24x/Vzegu4pz375ItgBobjTxjTF7/MG
oVzqN5TPJwCWk/nRkDo7db3VOkhxStCHli/1fWDbzp4ARO9LzTgp5Q94w2kNg+r7VHcZpTzyOVHD
YYDzKFTOmknUsnaSGbeadIjQ+wABc5a0RHE8/D4lgTAaRq1e5Y8oIDETUAJev7pICdl+NBflFPDr
xbbhAmvBdZoe4jNJUw7VYwumVI5FW/ptFjF62EJd06UNnE+R6bHkjxMR7TX4hXQzLihpKb3dwEKi
Tdv52YpazC2vvevaeweXs4jesDlByuR9KlM/BzoTzUeSn4cck0Vg/GPSYaQBnQBgCc9fWxMP6ecx
unUxfd3N65smAgBAeq2AFIIMgGWEf52mx1UkAtFwj5OFVW0ipLHH/2Fs5LHWAMAo2dxFk0S5OlJQ
GMix61fE0Oy3vjI/bkOy0SC4/MKo+dz/aplBNS2gCWLpC2+xwqRkDv/PrMK2yBF6Rq8rCTp4afYu
7+0e/RCfD4o8O2W6BmSTYkvITwpVtNSz/dFn2vvQLjuBmfgEtjyj/3glhGaN3OgwuNzRmg7otsOa
rzcLLigEerQdgXOxNbGmrUxfDI2WMtLXZZGrkUteOvBB3kiUNVx2xhzqSAbq28nQCH1i9a1dztG/
DY/Sbmsb3EPDDpDEsPDhNBdi/sjqEiWW3miAjGcKIBCglDn3Wwr6PKc4q3lwlrS9I808ZZ05CgcS
5k1B0RlfNBG4n4v6CuuqZgBI4y41Nenbgj/lyTl0LkSSjMvkHJs77NQKctHvEODEdpwh7qkkYoTC
ImGtgkyPmOsO71J7iF6IefS+OX3HVQwSfe4ad4Awy4dZ/Fxxq1ZzD6XQzCiDzfEi87f+s+TxCXp6
Z2o+HsY+5yqlbTG63duaQFYiqCY0Ug7r3d7nSdZasw8xF8akdibadKgMSfDaBVKWlNFShgNIHfVM
p3BZmY3dwq8WSaT5J8/9z9fFFhxXkmPviXzNwNjIrqHIozWAcbEkBIuF2YsiBANIRAG7MJUDHUE6
RgGmP34iJaWEN07niX+COMihHQMEvEygUIa6fFvzVhJMAHlejoIsI1EHgMP0U29ZdQr5st3vlsuH
PHAse9qD+EjKxZITxjTVIY3w+GrMWXPRAxNMCY5d7WdOpvpUuGDPd6tQsy7opN79rrB01niudpMs
oHxREkDC6LrrHj3kZxSjgFYxZSNdhZxU1cmesdyRp1hrdeOt1kgwZ3JZAJAfI1MThrLN9Hd+9mFA
gDt63slZvNt88YQs/WdaaDaWNUvbyzjDJpUhudu70QvwbEx9MfOivKTqMFgQWrnVTnpahV7TIiMh
YtXSmOKQzeZVVw/rpe77jLC4nFXY4vCocPhwjowJxKLqpozQQbWP+YYJFdun9fzxV4JdBH5qdpy+
R9+uvov7Us5e4u0FBA2yi2/jCrhU2k7bjHc6k1n9CxgYFoNbkV6+0wniu1+0D4myispSWVInDf2L
tD7zcUJGJ827jLUUkfz8yOkw8rbet2GUv9SnNOSKrbLjLngmDnyH3yHVqXVV8BW8C5GGMF2i0l6R
A3bB1Cr0sxi57ShS6neeKXJrLSq/LRY9hV1wPmJ64r6o97xf/unIIaSRf+PRcsHxqrqQ5CXe3gvT
AmTRIOAJxB3ndzCZLp2w8R1QGTzspePy44qIibvuGsddi8JvReZf/FH4McIMtWBmNQ6BgT4VDb49
BE+TFoP9SVv8zFIiaXfauu4feBwlRuozY2bU0NgpT6i5kQ1EHnMN2IgF9Ojz6kL7lr/dqMWOySCN
neL3bRxhQZ8tknvHgIRwSFpFWmdDSREy0yKRg7lqSahOtwN6jpXe8qXthgZskK1txSYRBLcIxu1+
Zd8vh8kJ3lYhjszlOsL2OYwL0EEc2JOe55t1xPtMkZntMAcZUBB1gD7AI+NOITTCisdIEcWMCNe4
VevTCKNEuFV0V4a3DDSadg00KzR4wubFyguT26ww6z+HOq7UVISeC/WHBPgIj/osI34BAZ7EIfU4
QGxXouLovAoy3Xn2olOM6PcPBDomtzBLpfmKieQ0i7Wqc8XaPxk8+Fxlfcw5k9RyKYxY8a4UfffW
f2sQGmjOdCm1hOOxyGTkFx00qqX+qPCwau9RkaVrZ8k6vyeHAnFmg3zYNLDpzQ5/zJvY9UMhhGKD
5X8Ed6TkkSSqKWigU44zxiHwuQfPQo1fvY/f4DfOnpLo+fGTZvQ/YCBLB0PsZNULeetaQOucCLH0
quM9UC2+NUjVXjJ3GiIUNCoTQK0yXu8/A56MrRNoJr2nkuxfBrmFTWeCFmAkHPLNZsA30HOHnB0O
ogFZfXuIdxrZgntjclfLOqTTb7zJkj0C0hLk96w0QZTWpaEPqTtFoQcZtjGF4p5MvcbwbTkseqeU
BORnVi2pyngCNmhWwTjahv7TZJYx6VXAuRGInWqorbX+NUjDAksWEp2d4Cqlq1mQTtaJc3KVv265
YFFOsZqwPafRyjOVHIABUXX5Foyvr6dYleAiUmfnyH0GC6n9UF4rNoNkd1Y0o0RGAE/IoYqWFxQQ
yn6FD1m35NphL0abCvXDZAACYKTyl2mpzIsh30kmmvticpN7uSJ141NW6+IMAzTXZDdppSSK8Pz2
dUI1P8TTKc2fjejq/SpNASizzG7uxY2l5M5CsI+HKUMY/+ZMYgO+u95O4iF8wS3QEGsBaAsn0glR
esf+guDeE+zMC2JjfIqeop5tkBpx6kg73t2zUWCt+Y100mlS30yakzNXUiwgCRK5VZUlxitg6D56
M1PPdejqTMl792QetLnbqLmP89UO1mcFkM1ejydoz9lmCTVW93W+4//cFBnk4r2CQIr/fcoizIHi
crsPhrsvTmZymMPMv/d3kaW+lpX9gpwRJ1jxF7HB4Gftu36bKQA3ycvcsyrYGRKs95snyLU+bngN
YCYx1gB87aSludSrsj+zUQL3iZ07vx2xDf+4xUIlzt/KQcUy3OdjSOieUVEZVhw80DCvf+6f6/jC
QCNIxOzk9ZdzCTybYSE8cmMkhU4xGawivXcv9TX4joNYKwACeF0q1jIesmJa2gXwp/OxPzXQzrX+
TgQqc8Z6xILdJD8hX46NT4YtaocndCgbF2bXfP5cqCIcx/lLHPPPLg06jTzTSeFfBUBOKMR05lpq
E5+EiKRt6SkTG7YHYzH/Cp7biy9T9fX9aRWnD3pLACJlq3vruMRFdz0QgBvqByarimACbdwj0qPP
fN9hZgAsuDLxkFJ3oCpvqzzI0qR3qESocLM1XPlRPOhYGRoW0LVt2bRG5v78OPPSYLySL+sEwy6m
w+u3BboXV4apeQVZ6nnSveMFIt9xNL4iiPwmUhA7e2fGG3uHSNMcGxOGJJPxXuNED7P7xNKyQ4/9
a2GfI7TtyCDq8SECK5A8ejXmkc89mUkEEC1bkKcnzBnkMROAHYA3+nt3+AB4UvON8ZCbS8UMLCE0
Jc1cCZgWTJMFOURuTST8Gio3ipLWM/giaNC7wqPDNV9IIWaSP8Pf+0B3O/QxYFUORGCFr5/DZ341
0svH8dONrKKzMsGMULrY3w4EP7l+zPQTd7A6cC1/4chEpiURHGm4iEAd131zbNRv5FTc1MwO6r7Y
uchUtkibz7tjQUyuoXH6ae1rXe1TIP6WsfzvYB/pyOp9qnQdl4OOAteX4JAp/riec1IAj9FvTPVi
4DUM7cj86NPPjq5NfhcVfjo5PbXTrJeKfsM8rARasJYyPnup9uaP3lxiVQSYU8ISGt2KDN/zJUMd
TH8AyOsaWkS6hKSff4m5AqK5gZIRBSPpgrDnXeVOSeaKQ20MrVcs11lSRFZ3GBru6Igrlqa95iPv
Y6z6vVXS6pG4QH/4Ourh6UOXNPn0alJCaJ6zBavVf62FCYVwLanI4DeuCo7PMd6EEz/PFQfU8c8Y
yk4Kw9DhwqkjUtnxotW8E6tvn/TuJ0x6qCTNTzBbHv8xPFPdxIHbrYG0SFtR2gSNqHjY177YFUtK
XRelm7k5bJo89BkNdJrN4fPLSfYG2Tk0GiPc+qSkOE6nUzQpmL6Iqai0i9j0Ei3UyHCsyB+gtjHK
a5sCkrgdN+tS8Kggp8IOGUxzckK/ybBG6oWOYBi5KOq/iR0Uwn34oUYDNC3nlAnDyTi0g9Lce0iW
Qwem6i7X/d4NMkLSPikTCbgR3UKTFCDxV8mkKdf5xVq2q5iqNlqpGFGE9DMp2EqMuQfh4qDJmwyK
s6LtHrKg/9o76S1cXU+ByL5A5y0Ctatta76u4oML9YCGvQsaYQ/V7QB65diMtS3WgHO5Cyd1/VdM
quLvBHi2PGYGE4fqJk1zCboPAzGp9mE3qSoyjcmJsThzUmemYO2/YKQyavr8S7goNI2biiW7mkT1
PlaMQF6nUwrxurTfSrqPyeiiHTUO6/4x8La/cyITivGHGRu5KjzlS2Vu3cTn3nT3n39uxsC+16fo
PpWZ0qIBppNHURfMj7Ba8cyPcbyinP7s0R/MYRF3F+KrP/JKwC3F+HQzKClUtMOrCm6qFXtedVeN
VRCJffdRXBwTtqe0bvq4mekb1++5s/XgxaS9nqHqwumLin+ahbLMBURvFbODjXlt+r5xRZciu7Ww
EMcj29caYiy+uzeODkMb0e+99HFajvrXHh3uyptKj9PhPDaXOZ3wUoQfQXbw2j2Y0nYUem+u08h/
EV8l+JtN2yTQTXfMv507dQ9aL7xjHbdKsy1H1UgBg6rbHF4YQGE7swmc1jawpI5394ZkYSpehMgI
KnHhcR/bpEAdewDIDCUcOlqRtRaFC5XH0uuSuzWDvh5WdjCsk28+0d02UGwsqA1Htb0mOzd3wkCQ
pNv8l+63qAvbPiuJdUYDYPwCn4jkUkxRGRfE380XVMY9mE5gc2ScpS58J+Annzh0ERGPX9wQclIx
NFMzz6pUDAao4CPgM7Wkx2it8MP669qPjm/bC4KhC1qZA9fSTk0iSZz7rY98dyuZ676uv8VTSNoB
o/ABrXk6KT2SGHdvTE9lXWLXOiHa+/Fd9bv7AJDCj8eRd+84gMJod53WH1ZZrNU6HNhI4TkFnuik
Q2HgWsqD1EDs3eZf3xhcVYDgszc9gM3kcDzvxWPQ5hHvHUTcp3kYkxquiVB59YNRnU5Kg6GDTdEy
jM+5Ksqjh+OjKojUgHlgj1aGVMTZ9UP7LT3pgD+8rqUUVgGSSC0Efr5LKBOFom8058SqJAlww6Gp
j2tDGbeaiz12va4yfXYyhKgUAZnBeyg4XRxM+soFmoUmQ/J9m+wf+3BjCNMQ5NEynlJ8urOO1e30
p6baDz3VKN1hllkGT5FKmciZ1Z3/8oGesckF7GlnQFJGE/3Y6niJf2+tq9/MaMUWsrgDRHxXDN0+
y/lpnGZVGp316Oc8dBNq2Wf0F9HrZfkgMLJ/ljB2WmriRYXKYiVdy7ZPRb04KN/SpxosNHXlLOsr
tgiIwSnH8zJYZIRomwpQd9u65Gn85+nmQmnymnukCbX3OB4SwbQ3mUDjczVxHVjEg6QHEeghLExc
tsTasTBDcfucZGdIFhkhAwOTE3Lfj/D+RhtssFNoJiqof6bjRoClp5EWj4jk9Wiv1IEv1EKlsR0Q
AfHoAry1ROhomDWF0zA1C4Q9rTwXPr0H/KFALcZvtbu9eV/f+lLZ8Ns4ms/IGDNCKgEBHlvy1uHU
icDbms7WwyNJIasyi3x1uSu5l2Qt5gmC4rYURxLloo7bBojmfaoLUvJAL3CeVapP7+eLBk9R0yYe
cL5QItOMRbumbTWg4B9YFJTePB4Zwacbc7fJx/nJzngZZNM4ZNgc2deoxbTNjVfJ5MYH9X8zQHEZ
K/cB4DDpdcF5ZdQI2VHxzGPTFqAfvVoJYAH4mDkN1neN3+Q3AW90lLyz+GUBewLZZFQxGLyK/vDu
SV1vjFLX6jHOXZYb2G40bXEl2S4Y3x0MISMp+9yxXiEwtOx3tFDK+gc4/RyOk90fB5rtRzfkHfvj
DPTPf+8bZ6Vjc/XJepA7uGDh/Ajnv+OAigis0L00qSUpWJwaPEBu4/vA+k39dlDINXGxXz5ONcgw
pVAVxQFv37Y4IMi0OwjOd0YhGHiSDpikl8OLqPO9/fmn/hJhP3vBLDCjW9OFpDpxIAc05n6Qvvr5
+rYjmOw7gXYsNMjfB3yg0E3XwjOxQpOQf3BWtpFEcZp/uRKEXFlWZQvLNeipqv99xoGjqBdAnJla
y0kyVaenqssMluLXmuI1uozej/ZXoXQe5xQouEGpUZRhuUztW0oT5Act/G6Sql4KauVrnB4haryD
Q6HfckhsT/gFl/mOlAucUqhBQ2caAE1L8xTt72B01c5aKJ2ea7M0prYBztl2q/K8xShh9OnOK4oM
CFs61Lr3XGxMihjhjno/178flncTQB749YnwVbcFeoYHhu9xeWukD7mTkoDcevroXxjf+ZroEKE/
fBYKlj5NVkdtHX2whg3/FP2KJ68930NabUhwsdxrxAdFZJ4DRjUJBydOuv3rSKqKBlQP4P+SwkCM
Mv1FTEfXh+3vJO+tYRaroAqvjeGpKx5N3FeC/NJCGFzbo2UXjYeguRhnTQBSTmRkZVMF3BYLwmPt
jJrOIRinVlJdmdzFhLCnCKh6K11LV46b3i7ovsXOROHTJm9LlZ2TrgypYbzSxf3JIG3lD/DkyXFT
xvEp0t3qz6+0V87TOoOf7VyJQlnriASXxIvXThuek8EwsDtARILfGDe20ruDnovfvWHrWX7SHS8U
QFURANtJXicoCRoYnS9xwWlTDzlpQVyaIkPHwlqK6fPZ3jIYcg3SclSAFrTiJYBmp20JrT3rxENx
02A6u539LlmwFbzawR+53tvBuhdUjFPDfLl+XksZM8xDQ9hqax7Gk0SxsgkbyKwbfehmvPZlrXJg
Re1eexTOPuPosKJY2mXL2pa2OlLqj8PEejKAYsV8T+a3EzsNPmRLFM7cpZ/r3Kcq0ihyrz45SdiV
j/VXIjJdbPGzYyptzXHEKqPv7N9c2jSEnwkn9zQi8GK49Ec6bwBKpCN8XeccqCapXWnsAY3juHsZ
rVThwNsJQLu00D2vHjj6UzvZ/lVjDXFD4DF4Hf35GXYj5PK5n9/LK+ardEW7grijfzPP7erloIh2
HudvMNHlfGiHclMA2zHLtcbt2lTfsvsKmTHLwgPc6pvI09Z+bO3QzUHiWbv4SBCtEVuszyIAQmuK
LP+n9iVE5n1Jjk1u/9JZJ+kDIlZLDrN5bHk2FEDzwHPu9whadNdmtmeIKwArxIAtdpuDQhm3GxS0
oIe88tjSiL2c+RQZFI6hHzAd+TyAwU1x5x3q9haJ3qQSelxqHmiB+wQyqjeSJdhsuw4Z7nb2vZdY
nbbaiO0u/54WX6DmrJ3XpZVl66wVb3bmcdgnX7xslMVCwyiq4BNhoW1eoepXSdoGmBDHYDDEY/xe
fsUXfpeCt/pLhv33o0ptsXwkLnnqZ97YS+nMbc4fM++g1MeFxiz7ZkHViZMztUzDZI84lzQtqpYU
Dnyt5Ha+vG/okGnVvlwrkVQTYM82CVjkyikXuJ6olPy946jh2bssRgziz4C94TWGZ5QvzJ4R8CXU
WQl+91lwDJotD/oqil0/96q++PJ4RauT+A16qjm1GAV6lrHX+u0nghU2LOY5v01owlTDQK3RiVxq
m0SYU9u8c3I7neZrHNtnbiv6YusRbOp7owc7aEvvhkGUN1GbzQmpNpVH432WBQtPQ6FLcZVYV8pV
G7nDE6KTDj5tsBDiDfQh8oYGAO76isOcEBlnkEFHZ/9x7RrGujNeeO9D7+y1p2juaAim+zS5T8NO
GKZNPjH5yCfxPZpK2FjLbxauyiBuuNODs8V8baQUeJ1QFfVNlVf5llbHeJ3urgYdGPfg10QSycaJ
phDiIwXuG5FYpzSVnUhs7vWzLIwZb2KvjNsdJfsepOiu6VlQIp2mB5i+UVLofdw4oqaojxsmjeKb
QIW9J/MMkXdWkIjmCCWT24fcNRG+mpdRkVHE1D7zDwc0OOaiWoJO3OXMNUBt0RrldufJWMt24p0N
qWXRE/6DjUvQLsUNIJ2FVal8g0E1tGHYu7BOV8e46LQq5OH3q6goUe3Bkw/qZQoYVIH9E4Hewltg
WJpLSxGSo6m+qVS2a+ZPl6/nIpKn0KZkDChKQG5vo4nAy9lceWqbkpMPXATVxHGfXCz+TZTaBu3t
qv6ROBjOTcyFy20JGGcdXJ4qn+VZ/bM4TDPdDTADghqFaKBlJcH+W3aFopdmQQ73npgRH85Jz3op
kONbJvafLDsLhfPBTKs1B66hInz0dQ+WBuY0gvzU4MnO9x8+63vA3VeEuhUIp4HOhPONPKA6P5f4
MPicVwlePSEkmEQ2UB8Ul3JY3vZ8/mvqj5MvD4vXuwENTgroE6wLzWKlD6YsATcVwuALlN52f5gm
g4U89KnZmJ51CXFt3H2GyumozN3aJmdJuWP6svF6lyxBUuE3I5fuGCOFE+6Qg663knbTB2RCKKzy
qjjVo7Uf3sMa7NrM7/xSsZVFMGyMxKIfPLULd78oWZTRaMdSjPrjp02C7C6uUb6+XgebEjWsdmEY
huAYHi6D2Rb+f+cJqd3xOTlS2goEO5+Q2IDFwJcj4vXyKpLrSQr5+IiLzOv1ChNEzGotSaPaxHKK
PvMQUf4vnwYpzr9eEK8kvRpeXeabKG0vH3YrENbUaAbhqEdlhLHf9i6BoLaZp4MF3Ps2BH7habSb
S1w0E1/9u4zdKRv9QEqNd9rl+GcPV44q1hVEg8BsRrzVBH2+PPlWlKTTJJitoS3rxNiC4hWG/BhM
5x0xGvTE2NZHxLlFs8DnrY5Q+0zu+ruUKQjjDNEIot2df7rgzOILeRE558gWAFflk1RAGjL42o6W
L1VHcuXHpfyMofApb2BfLr4RsYaiH8HZgyFUBcmDfuvUgtwVST2Mv7Z/TMK6Up3swZyT4U7DSDVP
hIyCBoj9dJwdF6/FhURJFEhdC4cSMxo3V/giKZl3I3s16NFyjkF/auzaA8595fObazddIfD+LEKm
7TlVMcUAuopP7QCrdsc4ZezYCFeuWJ7VfX7LZmq2N1hNtF+fmckJAEq9huppq5Epv5DYqBu6s19u
clBzcAJAStJHqRbb9mCe8jioeWgfG0eLelaOKK4GJa7LCCK8hby0ev4O4sWTcVN7nyBeRyA9f4mt
b8J3X50fRmEdLlfHHiODO7ZcxrHP1Aoe3PrPcTPlr6IFf0Q5GJyb7NthEv4HiWlaGVnZCfiL4fVg
Oc9XrzYeWsFQ8FpSOxzR9seWyeDh4a7fgFz+/yD3wJoLoQXibD5hGredum8Fak4hKRcX7HhFpIha
zF7UrZ5guatmI5Z1/G52W7oF+v/Yi0J5J0FVDktdhECSPxzBbDi5r2gMzq1KKaYzMjZ2Uy+B7xVr
desINmNbAabsr4Y1IWWKDPmDBhRxxQ7W52ZYOXE1YoilOi1XZiis16Ma1AkO1/Ztr+oRCsvIQ5b1
yUGnLuJe226zHYU0hwmGqCAgjIpsLjUq2hNcf5I++rlMqUQ4Z5NDd+N+Rq2Wd0Ll8HDKwn14MAlJ
xGPjruE7xTiR5ynFgInPMCmKRlOuQ4zkwGTCBxJa/fHBUdikVAPctVN04Ii9lgXDAcyZABUmtvB3
w3o048vSu0N2NHdFy9o7mJMBo8EcLTogtqWHhTlOPts+9K0ovFwTbCKqhrRgBaPrOkMkslz7qCXm
c5hx28SnIHHq5STANcW8jxv6KEHQ3KXQDtOWIKPj+WiUmlO6gZU1LFrCL15INUz4iLnxbOZresDd
GCy4zkElvwvJW4VJd0IvqvECoRmVfPh6xRuQrI6LRdQK6fmHwVMZizKkaNwvq1aCv5zYYoK+CVx/
IJUf1mRDl/yipdAySBs/SLf7OKk41JxQlbZMwi8dDIg9c8N3XiipNocS+lR/iUQjY3pvOiXCmWUl
yttaQCNiSsWnCamUXXPnM50HGVCFvRdwokeBYQ5lhLDdujNRJa5uhSmZr9yLuloorbpO9f/01Kak
tNXHMdJVBPngRWWvbjYkz0jlT+1liPDqj3vdK7hqqo23zLvoyhm8ypOPOh0NaA64EuxDhwoHOqkY
te3KgxZ9FdIfzjo0Gg8OE8fXppkzCZBsyfprDXXjXVCvX2x/nHxqTEuXNTuJXnhojs3gnLLbK3qU
92IGSdAAC9SV/e2l0iz5iveerD/YDM7zOTjmVW7ZvVQRXusjJf37u3y+iCizgrIiVmWuYNUbAr6A
Xz7OBcwO0RnV47U4FqMn4Pg0WYicFzTKv6VWfkBgDm4k3YbrZSeqL/S+CgpidWO1WZ5BvHMxv1hj
Km86jbisDv0e+StluRyrBparmgkPc8713BUUXKqjU0RXl+b3TUusXasdgU3Z26nJPJAUuKzZh/vu
ZWtVlmvLvaDaysLc3raLFVh6cbpXoD4nIG95se7NoveTsYz9sD6S3YlWSjpjDSOWzUh/BHazAK0L
5wrysKwE5xnDn65qmx7lTrxPNiTFqTdUB7jIgic95h54bNB7TpXgPTFZlksxvuyzb23Hms68k1AJ
QroDLdyhHRA+fz7CHyWEYd8kD+R1cHCB9pyjKQLPf+ycZbK3s+QKOGyWswf9HbRAg1oDwAKOXBEU
hnKP0AlyP3WAUPo2Jc8V6czZPR1/gO4bKO6ZEkg6HOmiaHgV1C5TnjpKE+T1sQwcSh7XOwMMGbSm
tjR+MaIFM7lRPolzzkm3gFEx5dWw71XMNcCGEniY3U9gtNzIA49RW0dug4103GdfQ0qCreaJ9Aaa
SBB646iopwiwFtnzmTMMI7C2yitdm2mONiWMNuI9koqJN9jbyrgKyWLmypSJxHQTJ7fxg4fBBulk
dgvgQ+xE9heEKkeeqVcXyS4XnBGMEwZg7fXD0rQx9x6No6/cP086UOnmVrJPSdUYvOOihzD+/tf2
BYIfEr3wv93s7TXFA8ss3C+mtVhB4Nh1tAFSRpbR+zGzh9697D6xlAFo65eOQHddb6c3Zd3UFgP8
LCCZZxXy7h6SErEDIyd684x8VCW+4PlT4cPz6EbAWsiybyySfm8BYluSYbyNZqe4i7Pex2bOda1j
k0Zj0UawvVMBFPhGIMthpcucEV8se4YrforQTOrpfzS1VDCbTW2pi5muhZLhbjR6v9NHu8INkXjx
Ue4o2zwnv/sbEWr7Du+TBvb8hWab/C96ZcyOi43vsweAlDI24FCNIFC96FduORyCBGeDOqH2kKRs
AOPXsBFWLI3LrVP9tPo+XPQK1iDteC/kbpXg1ZLjTD6mXkPJDEIX/iaGkig5qqb2LkPc1zxZrPss
XlJY8FapZMhmGwThZRuHjG5kYvJYYFlIxP8UTFWFDW2xgd6rQOgu9ryXPyYJJfTm1wCnMLNIzzY6
9yaq06Yy2ocayR7wIPQxdPXRsqm6qFGycdbWGhUOlLL/eG7HRhCs7mSSPgBEniw4jJeeDC2qXwu8
os+h7USMp4YR/hKDqZyFGx1wKt465Fl+CDGB288UEYVX5JUpu2sq9N4PJo8eMf+ySIRKhlePYv8q
/3JcbxGOaWH837BkzauGjVa92v3l5ZYgZF2XZZeMa03t56OB0Gef3Na8nW1z+IKH1yQJhiMwZYEz
+NhnTddRc+rY5jAIRXwvvkfq9AaNqBJ5hHqpscC7OFjZoUvk+fcQ9XSmm6DPPy8OElQVAs8j1ELP
PsyzAcS+UEksdFDloy9RFgZFn/M4DCvamOn8djiaLILo/zyZSUMCeHdlcwwEaeGUOBluCxsOBZ4i
hg1dbsrhk7iwRtL3Wqn9u0OGCWRdL02qw2c1KElAVkDpVy0jTnA4o6m2AliVyc/z0i3SnmxEOVl9
ChH2hc86twWstx/npqo9vZFCkDBvkI5hYFsJ1WHoZ9O/ahT/eemkf8PA4AJk32CUOsAOQdtQ79mL
zE6Y/33jzGxkq7qvPguEWcd+ruQqNUJ2ZXIEqK6kBWLlBU9bOPcWdcvT/VljaWrJl1EpCRl9tNgz
3SXx4xv86FbnFa2P8/Ei+WSknk7yanUuY8wejLHDwJrGM0y7P1TKGGxD1O/9w9OVFIo/yW6KZbzO
c+VjrmxRXSTTLr3dP9Bj+pi5pcr/H8tGhZBGXJnYth4fH9L5KLd3fMX6nmeP4zVYPOEBV1m49w4A
kZBriH8gCAKcCPjQOo3rw7nKKJFm33EIxziLlKb1Iqj0vDmMs6neEdT3hqzpUTiBSNCFrtIAh8Jg
wE7ajzBm/ep1qXWDGJfmpTi/ncD7cj1OXrmMrown39pBiGdEV2tJIEFR2BGXJ0r/6C4r3HEiSIGR
JC+9JMocivQdzVjc0MFRFx7tRa20zO0pS5XXpazp95rEY8RslV5V6zYjD8NqQg8ppmQMITVp4uCa
S4f9ImqxRaEzx8DL1PoBOM+m+UMgzN5Oxm1ykCNTbyIM78SYWvvUgAFWkM/Du8jK3v7X0tZrIycZ
wwYEKbqPJwxIEth9nMMzj22ssCVStQbWCBwtUZI+dVKyYz+ipc1wv6ArJ++Dnj3jYVog5aQ1k1jP
25AzsSHMNbO5LJIcHuB3DjeiKppYO25fNV12SbK3h0f3r9HcX4xik/uaqKYgpuuLcrQuAFVcV0jS
wp5QFgDK3zvIL6pj3xfkGMVKHgoXjHaxr2DFe7X6IANlFqMNgrXpcRDFWkGhwxuWL8mHY8GUXhmS
0BPuC/OS6UDeRyiymN1gJEIFjEEngvkWKgbhtBGjD/x1K13PdwxKaHS+pH9aM15LXXY9adQFxA8Q
U6ykoWcaAPf2waaF6gFyRFfhK4UUbvjnY+Xlq09J4teeZqgayRvzbRSUZAtcNvDNd2E5x8lT7udU
+wf0G86Bg2MXeOImnmuWnAwRE7lG2MjJglMs2ANtkqqYs1s5BdYWCmdvUqgvVm09faZRRM4AKKGg
a6dZHe86n9A7pt/tR7PCPB7w726zy2POc+Ty3H2Zo6X90JAbUdhDII1vU2ZB14EAbcBEMjMJn1uM
WhgNdfB2zrptO5k5Mnj0zvHEqpazNro90ony/7s0UOSdC7jwn/MNsLng2cL4PUSIAk8tsC+ZIltH
IrmUk1Sp+kdcI7WXmK38vOKOO9WTEXyLtL5HIgZNmFKAHircc9bbiUSICoa6X8SPYqrm8ZrYYHfw
63P62dtoz+ly+gyDtNBYv+OAFVrYj/WT4+Q3Lk7IciEnvPmDByaxtElotuf2lYlSIcdweBFoPHNY
rV4nY87erLhLb1s57Q5JW2p3ItMREDZHejssP2mY9w86PS7EttZKP9truLrEYIrEaYqkyZg6MOLz
Dd9mnHnKRT3plYcsliUH66WxJ+KS1jPhi8o5Y1oWwkJ0wXjMI6WUPydi0JC9+mWuWwhm5sihct5s
CXZCsOdDRt6IWL1imz5/OKSArbMt37asXUFO/owm4zcNntpY+tchgPSgFUmSjv1rMkzl2pL/sY0l
tj7xLYIPXYRElemgdsUNtYPQnuMU83L4fcvUjKr25JIPvs2MHvMPVLk8GtMXPaQGY1fJ0+Po/xw8
WjCGB8mdwrPWjh7lD3lnnhRtVe9s2aKiPk4lCj/kBMnESifg4pNyyvhtFyjqMkwCH6A+Emqn8vOG
aI+5sdFc0kb+3w98xSbuxZ/nEu7iMiob8Z07tW5dXSXI8aEdBgjEWb5Ih3Lt0+/bELMxDBOd0Td1
COTeMH6kSQMWl+z4G0D9fWRYREb2bTaF0kRhNaefSHOAXufAN+Fqx7T3Uz3xcoObDOorb4m18Jkw
6dYCC0QkYvDSuFlH3vJoPsKWdTt2MR9xtpAjNWowVmKxAsA+UtCd3dREXzAurGVvulQt2131ms46
N7rmbvvhQ6BKU8N1PJJzlqOR/rGWJWmh/MQ+l8WucyT9ppSg0Pb2QgAXSeeU/jE5ms22l46stAPU
1OvLuczLIMjRr5/DmDy6aj1b1uazpv11UFHKAyzNnLW8bZZsbH5o7EqIlbWUEeRB1k9I18hDjlja
jK0bECoZNoTxKr4jNWOl0gOBzlkaIG1sjmZOByvH3cl4pYPaU6HEbQqAZK1IeDuXjjwsWB6kLllW
KtqhuviYtTbPaXQe+/m1kP0OCbQj6xy9l78mWmS07Ej95ATM2Nd5XB3S82WdGIXbqzSIgpjjp+rQ
BwYPjOJmEgiiiop8OL2R/JFf/aY656hZJSio0/W6RD3+bGbYqv9xBxsn4axqgtm5+sZjfRvYBhzp
BtHd16CFyjhTwObBdJ7enMjtcjDHk9Jy2jTKlkC7XTldDrqhsRsXxDyi+HLoPNv6C44T4aXG+bJG
JCLQIpaMdop7IeSBOrO4WfOjl4k4DaSPmzp+y9yZ5X5CyLEhHbJ57vcNTcwI5q5gLHwff3UcPlBv
D4b52Erh6nSLmRpJYk/cFVUWE+KFZWDCTd8F6VhmaekqzlppRaUhLjH8DKJ/bdaYmAnBivWhkiV2
fbUlL5JNo0wKuHjBO5V6qSnqUyqsMW11S5bvbvHw++vHCARjI12fMBorIsV8BIuc0C2GeNrmfQbO
9gyKjZZUhrML4WafK2tS5/IRyKKo7m9oCufxbj4GwwfO9x3ErBnpgsdufNKtf5alwtCA9iSkH37u
EcGENfvsDQoEU7IU4EPiBWJ/yNlRW0BRH2wOxhH6bKy/nypTGctog/vLZqTyCOx6vF/OtKIQuq0Z
2JXDf8VCqKdo4MNPGlWNrkI/XwhkLgiTY0epQjqJ00G3l+/p1Tv7wgMhe/EOj0yUmhVdoBoXHW4u
q8fNUWhvICdYt1OVxIg1y37AcJNOFFcdMuwm23RF9SkESq8Kbw5BDvs+ahYBLUX3sQBs90VBJHad
A+6Opn4URf3OiYOqDnGKdUK1GdQtcdSZQBsnEucDKTey+kdL0KhxtrVpOCj1c88GZAXtFpSzdSMX
sGGtww8IwP41vJ7pzGqAXyjGdKhWEvOeRyk/koJRIkRcNqwAsTnT1j56b0zmxWkCICPYW0gonngN
lYlgjiOQ7TXKTxZBeqO0su2V1Oupdwun/qciJBEo2ZoL/irGAQQCknowZbSmtqjEDV4Pa+GQYZRA
lp8SAUpAr7EH+CZJJqs76VWU5CkmGGEjD1FNJkW9zg8ju3i83oU1oVx/hQc36+b8x9AApNEZVG2/
LwyAFY9KuqR7ApfqOeJn79tdyjGgP6JEBWJuSHPXWppMZF4g2eiUz0gZ8BxCgsVRhU5r0qiF0p/G
OSRsLMK/n/3SM2wWL0VsvP2iXO19AHn5RPtClijKjFn1c9CpQCBSG7GCJJOA0H2sp2LasEqPzxYy
sSN5CnDlXVbDpzj0JyhJgg6Up5CT57brBr2541+AKmmNOOyxbnQxKLmthEohzaWY5f/MHIoojujl
XhmX68hrcPyMchTiXUZcyWk3v1AVtTw3tLzBhbnb2QB1cU43DJbTdLEMFpJXjco4asgG7ApbFVKQ
czmIeWgdOeJSBsYNyXzF4wMjWt5/l/Rr8lNs4SQ4nYkQxVY3hUowUE9ft6IRXlj9ptunEDHmN7Iz
+69JYDN/H4a7eMRBsf1opvX9Rw9QcAUGsU7mnro1N1uPZEWwzu/YiNkbkrbpQrCRcB4XttIvk58W
piCjXSKopgRQwQOlUh0MixbuB5Cz89/IV9YM3Nz7pF7aLseW94lWMsXM4KCLlOe5GZxXuBHoPCM0
yr/lPyUKoX9L3n8t7g/GqZIrXaMDIZdZm8KscvLGLrwsAHpBtbgXV+K51GL7gWSnhCF9LSOV/YmK
JXakkWCwJZYrGU1oLxFppC0v5UVl+MQi2/hD9/E37xQNkuQct0KpdIgNtPCiDzShzWQuaYJM8PtU
VMJbAZlM4EvypbApa7giQoTEwdPv3o5BYVpmWtuz1ga0leYdPYRVb+5yoaWO+jR2fjk0XDMETRod
TXEE9T1/6RaY7lc+tU9iv0awIxd8eGlgaosERogeT+0Hkk1dz+V4Lkvjk7l7zE0uX9o41YpP1jiZ
EvBRH4FpZTkwKw/QscUrszd05RVPq34unLEi8DWDhbSThX9+G9sgOoALnPoGu2oC/wd4Kx25ujMx
MlwBsc0V4UWxa6eYma9YG+v9qxDaeBFNZAhjT8E0UfYRmwKes6PVyyU3IqFWAoxA72L95Qyo4X2a
jghQn7hQ+UHDP2c2OjdoWuN2hPmfbsJVZIvmXpVWm7JzWfr8UdwnAphnHEkzv7HOU2NlQueCtQQQ
N/QM6QWAHHJT4+yEwRtjNA3ZcjF9ItcBjBrfJekb3RUkOkd+c3V1X3GA4ivLH0o7erHOqysxaY+f
N6NNDAr/kDBdxN6wszs3tryYXsff4orL9bLucZgKY+WDvzFmetzj/EiH1dVfYJEYNPE6oNlrkfdA
4WPSZL2caMesbovj9dIhQaprKnd7WhV43im/etky26tWX6uG6vws6x6Yf7d9u/8r+DdMCiQvIFDt
UPJNXT5+obdXEUScwMCmAc/irfK1xAQaXCG4uc4UPD07hogGocBP9iFEQIjp5+XCMX5HcOyWPy7V
fjM4bCP4J2+xJC9JW74P8hwlA3RfVM+NTJOCYrrbNoq62RqLfHCnOnTr9Wb/gzym+nCkaW2F+Vqg
JtZIUtY3uhJ/H4BL2dGAAwnR6M+7+wkSq4X8gbomq+1In+FAfmhr2RCFDE6piz4nEJ0yd+/w0NCs
5PwXfYPU/1DwKkrV9MTu+tqEHvXJCAORh/zorJtsp7PZLcnNfNtjmQn0px5qx3mSm+2WTLqBGUja
rGpRY+j+xGZcqHCXPVh02khyIPF+dhw1K195O7XLCZdkCWWSwY2/3MNKNB2rWtWrg5ffT3AsoQXw
5sqFsWaIyzM7cr/fnW+NALM0vMV86rthpndlk5S+SxcBSt4mpVqgytgZpyII+eCGAlnmj6utU/cq
8K+AOUCW5LZIWGsvh4Cc/VU9IgyILyhineg8yu0BmZNFMHqyHimvo/mwJHXAV+x1DgnlhBTZ95aa
LMSKUW2cbIxtO2jGhIhZmcJEMz7SoTH+i6A5jFaZU/0D5Oy86jl+ho3Aq7HhSwi5MPsBDKWNY4VN
A9wxf9bMz8Zm2b3rhYDRjFwJebgSajRxmb6ZrmtDRp7t6xGExlOWAbo2OrcWRMy1dXzgn/lOYuqX
Z8LX51X1laewxujV5PfVDuwFaWpvUVLVUEQJMdK7lHgpHjYCBX9CeX/miNGHXYUV1EQKcsEF1ysg
rPO7ws1s4FyAYvn9qF+1VXpi/V4ErPT6u+KI4kv9+HFDENqfz/TJN2W+qwus9gMjvX+bDKKBreTJ
8ZD8FyN4zRckj/vygsQXFiOi+05O2HfXU/hqwhDkMHWmeGA98CkrjZkG52iQoLHcWGqfyvo92yr/
4xZAUrkD+nGDV7uK+fIm4vJczvl2+PElU6queDmvOu3adlBqKZdPjF5273oeRuQfK5fFRac50mA0
d2RyWpfau9Tc6SfDA7ngtqxOB9eTVhAkPtPojr5O+1OtYq+r1nFq0t1qEc2HBTwKL55pkTDmL34s
lFLOSPk5/qov3dVl3ALkwp0sgwKucztqXbkcJh/GUjjoQEJCrEjMbLVH2T3Ohuv5lYg443dyrG2a
YadvdXlYXPrdpSkuSyaZ796kj1Onx6qkSJawldzuvF67MRjIWXnlhCppxWPNz/3LGR8k9ZlCmK0I
CUB7qwxYXSWr9JSdB8djhWg30YJWNfgLGXm7bfLnGuUvkLmSmm5nJvBmDtA7k7v7+/VZ1QMy8+0y
CCnf08WJYBJOBxq3DyIKO4YaD8w/jcqMjD6H+MKiGkFcEkSxgLvThffLSddq2J0+KsMuwXIpp8j7
muq56qxohcJP5xkXnNQbQsGUutkWTL8aLqUefdYwsTdNUA/P2GPLrDkDrZRc5h2kgQtFKav5TOI0
x12nRUP+ebJswIGj8bBXauO4CDkyeMMuzSLYcYIFdFBeb5pb2Z+VrAZOUvyID8y5+97H965lb5tI
5yKF7z2CuNtDvw3L0s0hu2UHW8LIVIPVTR1JCFDCER+W3zFKrMpV3yPbLXbuhksapAUwy9otn6Xx
AXuH+q+/X87DbTyeMU4ReVxsi/+sqI2r2jXE68TDB3t63V6yRy3467SdzIratmKqIAgGLDYeHLfC
ob2LCBx9uiuunLfzuZstg1yixElu+v78GxiucUslnuIQynnA3/Es46UBqEY+MbYGGJyZ5HDbiQdW
QpK5u8VZYuk0zPV3C5Hx4dWxKUIkkqcGpoGBOysCnff6VYleh/2TfvbxIpNmNNzKKYulCvLBq8g5
1y2DMdToHGwGY4NbGhIkDuPdL5sunAE3jEfF8jp7TgAI45nLeeHvD+tJmAoTUipuHuGdXqQE9pCC
hr5pYWJf6/9ZymzcqUxw9f3Mh0ZprZuOpEsaAuWPgHtAyD8v6oc+Z/Sw+pRQ2RUIaOjMnMR5m0CK
OKyfdZYcMHiWBEcpfNbYFCd2KtPns3RFqwK66aICFq6khHNqDXQWJ1y2NIwVzq2d9+2wtN3lbglO
+3KPZDhWkebMHj6UVYWb3MGaGSSDBaotvWMz40NqiKO3tKY2MekByg5Lkido5TiqyAVck2INzt5v
qOhSp/gBdM9rJoxLDN1W2h494D76aJA6Uxc0BKdwqp3zlSyFUMCHFLslVEIuaPhAWxvzULutx/9I
0V31o3YVenCW1hkKlkg7TsLn6dqwXnnh3X2/0hFLXaRaKBVGqe5JEJF6LmMkxo4sPD4yBkg/myXj
euGDckNltisjm0+cbh5b+rW64dIjHvVyNEl57J8H+efEkXa0slVSB3oYD0v/n9FKQUuhug3TaOqu
zwZ7i2XQVHmHit31GhWH4JWKGQrQYgFKXefk527c7AkScHtdUupciDNOhMfAowqQBfEv9YykKk/A
QbuAgAiJ9IDldcu/I2/goPKS7fKdbVI9lDhFV60CInX03TTDuPhf8tdhPhVVn2eJYvKkmQ/6+hME
oCOmQUmHo9S00JgFTsoQT/jF3RfmpbkTMUZo+YhyroEEZYaEIYbLXRwP0GWNjuFAkGhSadbdxTyT
1pbdVJT+JNLuwhm6juHbJbbfHBgtpTdP1rYqjvaLNZCv5xGbqEpKFrHUXYkhvaYIDI+4o3Avl5EC
puM0VTbdS/1lCsmpXAEtxkIJxoEo3EMvp4FdC5uOw0t+RUNl5adDfH5dNIY/Y0/4cSwNQ38RX6/d
btROqECpOFtdh5DLwQrRmCEO6+XxuFncvm6lqJaUbPYKP0NlihsseIDkI2tul+rYoCbHZBTHOf84
WB/98jERpaMLm88MWmExVDHqEu7Qo2Lsn+QSRG74AYE77ZSz1um9dDkyBxO9vHTLFVJ3nRUO+Gpp
1Z4PjJwbkov/2pta5z98wmmuLvIVFHsmGIxd7b2J+NoTjLwt58GY1EY8J4Z+al/sk3qsgyeoWA42
1S2+0vkF8fbBImWWKHlORrnT5LYNwml0Cs8QJ2jLt9ePMGdFulKpNct/fqmFwSNjP7NxVc81MDWo
0sX+PKeDNjZv503CQuTRFIoPVgKdfOjmaW9qKHXSQq7nfCbxDegThlhpFgN2dRgNyKBe+fpfv+23
sHT0rc27SUPg3MIiOnh9PFl6HRBqCMDAn+0Ibfv0Gf+lg/frsdkE0x7IV0J2RYgKUR946fLPcybH
MARLZQoQr85IvGWtdgHmIh+qDBRPtHLwkFyqAy1ywF89HgTIcXwwrgFxOnMqoNp+JiATFoeTXjLu
MC2JVuM7x4hVcxlpiuswrGP63TPjzU19s5l4jUovVYpZDB6Ge+zrZI7zItKzuCXsvvHGju9NXtcH
xPC/hKsGIqSZ/0qmjsLt+OIRt/r04aD9oD1lXAaxFi+FZ0o5booKnkJBnwxzm+UpaeN+VzWjTi47
PSHP0UTOUZ+jM0bCbH52PMXlg4yqbsXLj3U125RoHKBPuvMBSJUwFGiDXG5IsguK8pqoypQtXU1/
hP42r0TYy7qKGxn9zdQmoGX2IhIXk1MiTe2ZIw8TxemzWqegKkzIRQ7ihNxhjykpjXx4611KI5SX
o1Lmrm5lA/AYlXM961i1qJHmC3Xv4iorwD9su+ybdQfI9YmLT6rNktO3pgmQ4PG6BpbBApaeNqCI
swOF72VPsTRJVfBeHiH7/UtgWBEqrUa3YHsYCtyahtq/0FJsAsne9B9LC8HCj04ZCrc3EYvL9uY5
1AihwYw39oqEJtJw2MEhcciW1Um8SCFl1FtI/S2wC+nBu/3UUDhTxnsjBkOhcR5JoyME26YSWBje
kHn8/6Om1+B36vZfsXAQa+Iw+36nMKMRiWzeX6OuBCYYrO2H/y05qpaq+ZLTjrNlcDL/fJ9fnwcv
ACanEIKA5+xeLdN4539wHQv4LMLkvSWyr/dhRJTIzNwmlBpNLDo+1poGlJkPBoLFft/dpU4uQrPp
hddITtD8TRbXIyOIYh8AW24n3jWLRR7tdHe+MnM7Ti6P1W7cUoeBeiEi6yij05aC+QpWrCXCrV/+
V2pziKcZD/yFElU5irKYKsKn2p5czWaaUOfKiM4IFD84qDFu1DlKw+8kcPq45Z5tUw1gmrbdyybg
kcZrAm6wramtdvKPVmwRbm454Te+UGnJLWGNQS97Vw5G6ycr8ilKsZaAYbHrffbueCTVPkNrFrg7
57ZhSujWJR/hWOUvGbWIanOlWb/uVE5QFi7B1PdGdWhPYxA5mHkqD0OkcN5FppfoMk6AvyczQbq3
eWn9ejxqL9rg5NcyjyMBDIsFWMEO/5bS9ysuddqSh9hleYl5rsYhwgVPwscnBQcIg4X0c1VnbhA6
XJ0IWTQJWERu25wgAUOyFG62oU2Rkz2WA/e0TJQs1mFMh+kXVYCJ11cSk3UuksoF8zzTXZUm1oT4
AtPy313OCn0AWg42VotQ81uUqA7Jq0LF8mjRNeCEa/0/j5rBKpQJPRLzX0UeTXiauMKQ0pC7lx1K
pIykGnWGU2lXGN+RrEsraQHQV1dYZHdbw3mlpXlCMy94THsAijYHaZkrS4hdDQscE+v9WQuq2l7r
P6GplRHItmTV38zXLazqkHmbFqYsTTTYYw4N82KBmVMHgKhSG/IX1FWFpa6IBuSaoiQ9Uqdo/oOv
70d/2kngvWzbJ+X/B//EoNXna3RRVMXV4MrzcxnI6+4+2VVXjBs1RzSHUWljnobmWkMFblNmkRgN
ZvwDTfSlru5hkkzz73GLYGuFItfDoI1JRTpOSWbZjDDgWWh3A9N0Yir2LGOOrrX5AiGAKhkRly8F
+ndp0iigcckuEvEQ4LXsbPNYcMB7khCEC9Q/cfMpILbUzdplMT1WbFTbf6NjqDGHrsd6dJcCZAFF
kjdg+PHs4ihJ1abaxWYwBgkoY458H2cBl0shqe+cCxdDsePO9WiagkYvoPYjbusR08qfIBb3nhEs
IKINWdMDmHFQ3yakVPMurLrxUloXvN5igGnl4uL8oRhkiy/AD9P8SRdP0WTDZe3DGkTtNNAEJtCh
Imk1FjC9ayfp4N9a6k00Edh6vWYwYEUgt0mFUEL7V6S9PkYSGQnE+PGWVyOciocNX9l1AIRZgzC0
RfkbDEdtjoXIeSBcoPCNd3D8RwzlY/lg5avfRYHUm3dysn8o8h7dI8qKOe70DrDrbNdQszLepvcj
WbD1UL+Q4hSItIfwwd4mCf36wWSfP5gWag8Egnp9zSxGOIt28n/tbDOEw1Iu8rbi9M0LjIChvLfi
Zv85MrIZJ6SUR/L8uqTi7bh7FfUcDdJlkT6jwgCgXbv1dBHKkuK8SMcwAoHcc2zQAt5/VVQBQVYS
2pxwjhGZze3WJktYareMDCyGnfJ9coRQqJ0iBtH5/gcYAH7fQktIrDyP14h2ZXeQ9/6YSmx/6Est
+LRBKdvCCpQZlCVDKOWxaXxbkC3Sj274QPHf9u0AaewD6pKDmBUtzCo6D/CvHUgjcIZJKZKrfuUI
TtQVKjR2dVZW6p0tyU12GB+zfGntMmOlyQVHd9dVPdrIDg/7omw3AHSX9aK8H72fLEuPTpnmMdaX
66nJs9b6vMeQ9rAz66v0Z+PuzV7WYAtKzS5wZnJ69DoIQX1HtgmJKnYjcchHnKe+pGo/+WdIQ+lt
x+BNkEJWZia8JHHq9zokYeR8eC5JxlhwmDinJ8EuzgSqmhTkj4M/Bq8wvndMsRwGqh6O1bNr725y
FNGsvKKztd6BtqUymVNCM9bJHrbSrHdstLS/JcsYjFh3EU2hL9allvwXVboxjStJ10KrOQflic8X
aIbusIhYbBWptTJzzpxNL8r8U9NYsOCi2O+JyImgMv/A45zEncUYTaeqEiP4vDzMOEguhrZxnAhw
S+ZiSTGSvC8D+4b9qy9aPzFb646jEO+8zK90FOUdQ7+DEYDqhym6BqBrkmDZv6o/I/puSfWAhz2u
qZ5ccE/D5VKmZQqr4Gd4WEMEXDFxJhIzwAV8bUCyJVHHdcgJovpT+TIt1Myrm7k5ml6+0ZYwJvAj
Z98dUqaS6JWgo+cWHbJiKsnxu9cDIOIwrVlfSW8D4zSbKVjfpMdWE2UkJKvLYFUokGJVgyQBcZYs
ju0GNU3opwxVfsSrQW0N0HYLE0xNAnXC2pOJPPrvs+5mHOsDLaj3mHpv63TRJLvn9XMfwxQEkg9B
KuUsRz8ZD/Ax7k41IYkbFOaGoeY1sfLUVDfaQMImsK9V6d4eHQIMv4WtmZ/sO8Kj9Z+djpe/04pi
k+Jp/V0879et6ryEttc2bEBbY8GUx7DTHAXpTrX/Kh22AUdhNiObqKoQ0nKY3bhyONg99eBUSCZK
rlql/yPYRK4qK0brCQYItUs+BcvHckywGaiBAVQ0jd1DAuzOWX36EmlrFk1+Ysy7VBc1pmxPir8Q
Tncbd5Ig3yjxFiEWuTuCvT94Kb2Bqsf/BDW48UFUBZ9mqgKJJTy5aRkS3u1i4WL2VVRSqW3mGroF
ZtuAOktmVo7AOxPFf97lc4kEa3FzkiSMAY1OVe/kpW/u7hBHQQPsHDGV0MPcJmvlRgj2OpE1Utn5
GJL1WoExc5rSbZYDnfeB9tJdyHnHdXHejIZSYcqH7xoQH8rp/9PThJNCHA+wGhVQA+gZQtWTWYMC
v5bMSlQOdlMUF2hcr3Wqszh/vnQr9B+RkKagkZQcdY9eCRlxwrXs8hOXEUGw52VXh0Wb+uxmpqot
78al1sYGKiTwXLUbvbeTJ0Al6ETOjh73F4/0C6QeA4+fv6RZ+TuAEk49pgf38d7NbOMCM3h+vJJW
+UAkM1WXXStq4Smgy7H9WU8zcfVNyTBmj48IsnAmLy5fQygG07ju9fcmCoUWaMCCBLrYTnnI+NaV
+tA9Cel1xYFXi7KfHYfQQS+GFa3Ewi22/XntfxTnNeDbkVTMrf2MHDH1P4grMKGntDvjowTEsq2N
U9Pq7pkwxPoIhwl+2znrUT/NJvhA819JPNDwrPv4RI04LoL/D7vg4GUnWe5jaPGBL3HzOe/H9t3p
fLKPjrretN3/SLBkn4Q60+pgYueu1RL//qQD7rh+EsT+L50fOOSEnvsVHqqvMlpVamCXCVCrxVDz
f9eEtzwCWfvZSFBC9uKqOdOWTH0skLpgKRgCd8R0V7wKPmn1IpFEEU31wGy0CO6mYlccJ3IlTVHe
TooNjvadpy8skis4iCNkjiOJuVckFIpCRXxZ1y+60xbTp+P5ANjQOx6pQBJYyD/4GemnXZMAjs7S
iJ0H95whgkO1b5NlsBP7UzAvRUTg29AkkTmZMFMGtwKO58jQy0U98OJv71eBT12BvSHNy1/gVLVM
OvBmuLckjRg7k4q/Wr5vcYiFR4L24qaaPecWWUJhepWlf4Gwv6NX3MEB37qGSZ4RSBERsjNBmUrd
9uDSCWl8kJhLEBHikC+eF4NZSqR+HNou4zNNt85zQVRjKueSfNvoUO6CwgNMqKnJWpivNu44R46J
Qws0soJbOzXwwhsQ/CNDDoyYVq9/8m+pbe2nE31zXor9vk2p0jSXXjVCsqy7qPFdV1fcJ1DPtVjN
AgL0vrSlb3YfMFkd2WPfU/YVzHZ7gRhjYyZQphM/soG9TbTWyzpwVitgQYq1Zojsb2/JXZ6QmHjb
UeIraOEaPIms0W/EEmZLNX6G9edtA+IqRglI0sbwTvmEYc7DS5Su1y/VkyQHfE2z8RFwnC7hgD/4
7YTdTBst8r/EEzdyDrlSwzYgxJW9BmsXWrjL6T0Ptn/ZX1SMTAjf1ly/vgwdoe/VRz8/AWriEItC
nwR62CCyHwPOa9JSCzwmajmGfFhh051Q8V5JwQZA845WGkCTqfwUBZ8nhGZIXEKYJO3BDfK240BC
zFYmLp1f053PRIGYZ66S53J5EmF32FsqUrPU8o1AZaSBhuRoWr3F/CxXVB1y5OXijaLrSDxoIaUv
Tvo2tRxLE5I0qiw1kvwGStt0B5/YjWuL2UlzEu+Giu9CM/duEHO71Xko1vEdJWMXnGeAXbuMUM4e
46qZt2Ipkmh8Yb+jrl6BBHIavZelqLoXD39eqObN653HnAPJsYuXuEJr+wkUuXtDcV7YX3+txvmO
Z+hxgJuWGzZEnnkQecqcGGvmmYBUv9/+/S/zK8w/aNRen17+X4pqu0Ho87zghYCgYCMn/+JqVY9P
A6i46P+iLHtdp6JfWAFLqwnF9i4NWR77zmbHXA/4pZMWn2SRD99pcDbZlrzXrI8WiF6CdAR9u/JO
pcP8arkzpdg2+XETap17wPpAZLpZFIHYf4z8VKpl1njTuFAt6HwqcjGpH+6ePqyX4MDPqk/oBNiT
am71DGY3sfMrioks1WxHnlPxIFYUowLnsGTuWkGMemb/FINO5mf6qWrLIs2w2TV0xfbctXXL8lms
Z50xzCjvFnco17PX/Y03P+7OyQEDeQANwpB3t1wJWk/YO46egszWJpqzIgioaEt3fXway3g2h6b0
LbfySqb3HHrOmWqZDrQqsc2r0meLL5mg8uBzbz6vcOWd4bE8qFBbk2oMshyilMDrlqNTTn75Dzit
qS6rZSWN+Hn10G1zSLKsTc26ByHtOYEsc5YJjyNcPr51rmNN46UhT96To8xwYw4ewy8K5gQ28nwh
/eW49jGK7tEo3qZIs3a3pB57Z869EsgHDHXozfvMJW/Uwy1ZZ53uB4TsG0EBpGZQMEUnG19sx2JE
n6hNHXtzT3OsT0W7LWnrjmRTvxVnnZ/c9oTbPcNWchhnVpf1Jor3AALypYj1EFIUqiL6tWkUl5am
8wyibb8yyCwyCgYFNXFhbpTD0rHQMoXSZy3mnEY9IfDWWtfRF5a+Z8Gb7GcooDNf9rsGFGF/dy2f
x5lQL89Qv2vCDgIAF1Dz9di0hVH6G0QnhQ9d+gTDRq/3f9r/E+rL4DWKMaYJTWPOs9CwXPN4tRPV
EtMMHyi1hm1ZLRf4hSxWqpp2BJaCuVx0T9xTtPTh1sCx1N/9BFcMwktz2RStysGmCjMAcGvxWDdK
hCGZHli2RJDGL7ZQ/kYNKrBwaSVw8DoF5fs0zS4Vo4hsGcYXeGNhjxta3H7hauy2IEBeQCZ1Lqsk
lmhmukMvBbjnCOpqKoABf5DwPWPzhEzV8wBgbfr7tRvU+jCLEEMSCiLOzjCOkAVjO3rJGCmPmnhb
ARbdZ63iKm85c8pUWEZl0PQ+f4OB4zJO8w03W1zc91MsqKGF2/P3tegYkPuebS8xvMzgF96y13bJ
HbvEPpgwGuMAZ18wdJO20oaTAEwSiSoGlcut+IBW/Lt1AKDiK4Jyb2AIP5ZtseKFKprvy1Q1NPeW
iHSqy4TLcKpdIMf7nTnjut0p+V3PCpoCARvmw90yWtFcyua2KKsq54CLGmttNqVDRXRV1fGWTAjA
TmiQdVkC+Ox2TAnI6fCWNgHPOG+iXA2nZSDzxc5OKvgRUSKoFevkKtxdhJfkAbFag55Gr47dxlwc
XR0S5LGZOockqjOLrgiLWgH0iaKtt1FI4lu0KpPWq/GNm5OaFB0T4TZdE2XALaPwEwi8HUgkixIo
2nwag9vmERUIsbQSNR5tAFx7/QNCOGfPItS89tl4pcivTrL3Fw6Ybflax7CbZbqD50M1xQn8t7yx
A8fXgmFLHgm4uQCAWfJo2TwGs0pQ6KCxc4XxURcjqHqf1yN+9APzd+cp7yegT8YyunMwQtvPd1uo
70iDjV7BcyrjFcwu70spnHO+iI5MJ5R/CUhNERtQ1AjNHVHT/R0DBix4Nsm1y9V1RTtjo0CGWypi
sSVFxj67/8E4Eb4A5IG3SRJWDuKS/hlWDuXk5WMF44TD0MvlX1zwHlq/Huty/N7Gl0F5k6CJckOS
vmEMlr37GGgUzMnXGo110SEdrPOdBbc28GtXQiSzPLB40BXJUvuT7jjiY089I8lSQM6frwzmGVgE
bLNc/oaLeqIRljdTc3fCTL3Hx73F/a34CMh1S7HBlOcCAyPuWvDDu+e7v3Z1otNW6AtsIHd6Munm
pc987VUuJjB8KciOrZF/7CE81SOC9pFg2rJlEmPWPEkW1zVNrCfRsI2aC8R8xCdggP+CAod7pKe5
/eFqz/gn7Hq9J+EDPhNBvdMyOz2oLHjZCOXQkCCljjkZwJ1AwDYkwZ19jYkp6cQLP8hylfSdjBtB
9aumPH9NSYgIyLhX3C6GCF/SCq+AIBgOaxMkv1+rIuRRjpV7Vnx16HMYAksQrm6GKXvCB2wT/nja
91wb5EhjvPAbtdY2MLSLLBMhz/CjNFKEaIoHrEU7AXS/y3Nns7UK4LksYhwcd+Zsc5yXMf7Ub84I
5tcD874Dzbdg/FJorF5a2PUk+1a1+f7Sbogmg/Ui/nX8RN9jnKgmy49k3onkEB7yrQG+2czbmlQa
fag+MKqXqs/4Gxsjxj8cJtZ522arNpPqkTNwAJDcO/QyJHNWtXVHh7RfltsZCeU0MMpRLylOuD9q
kP5M6NwSb82GG+ShEh9LccfWZpl+SnC1g3W/G6LiGgQEHdS+qKcz3h7+g8i2KTexAsHxjukYmH/d
BzdbSnqeMPPZjyWnvRzSY4LMd6gQqWn1hZT3ZvSw/aloIhlyKJIXlHU9rc5QQEMaqYK8p9x6enWh
qKBLLlXYmV+huEnK4lDFfXpHIsaiAf/ITk5fi9rID1GLbJSqbS5+o+N7ez2/m4lFU8HimvBMhsSn
8u4c3jQZxa1Pg6cFHDGa8ZoBLnkKmaGCyTijWZ2hvDZzE4QB43sNUFO9pzD8+Wao2chUa4VNnes2
6JA1S5jaReQElC08bpBPn2hz8oE4xhXkRm1oohIlX7cEhKogYCdO15aw6NmFPYJ2NY2/40IXY5sD
vagzPFdPb3azEfTGqio8dbL9WuD0htnwYAvqAprjq1XCYQ8iA46jLn92gpSuM3qrnVm0Yn0oOwDB
2Y8uBk/6/6pedBbWncOTNEvR6YQstkKzPp1TVwJbhl4tmgLJeDhCoagwzboWr7DNe69ChvCLm/0s
R/iF9Lb4QGax3DtvbRd6SJcQ/WcZCnuHW3AGSS8ToJ2G36PEJBLXscLg8XhmfgFqeWHNQWxK/uZY
cq1R0WLpGeHEXqFZIl6BKk0GhLJPLphwcD1ruBLuu3+7V/sNTU4JMmRnwL632eQ08g73Vb+6NXf7
K9B0W5Lm5/G3UiZl46aNeOdhF5yk4HQcv83wd00xFGHOhbYwrGnpPTWuCZBJwobPmBjkEvVVDlup
IcLvnOFeFNbk2WEJkj2NOnnR/+OLgk20BfesqMEHdtGgxByBdA+XAd2qr1FOyiA3T/c31jXjwYf6
DJsbn0utf8J5LgUm+6q2X+yCryotzImglCABmPexV28piXbNpyRDoP4fSIdUvmCQj1i43+g0yb9a
VDedgF1BhFSoyW7MmF+JJhOqKXNDWzPngeL7prbkKltku+NXJJvar9FMNdK0C1OW4UtzSrMj4K8/
AVUAxMkhgrtrbE4B1Oj3hxvtv3SexW9fMBfOw09JmWcVpIxXjyHPzoeOQ3953Xqc4CrdeTu2Sp7m
teJngLuexZblMkQA2szws/JUdnyUXQ4bMRQZ6PsA44aEAdrfW2ydijtlD6RjpGx8vXzVOnlj1A2g
N15Memic57Xtx+mnYuRBzRuf0BukViZ+CTHG+wXo5D227FJjKyyefuCe9FV6ABqUBJsTGVo5fipY
WhdDSIhCT9B5chU+MKIPr9Uu50hTCoJHf+GYA6uHtaEyYZwV+eUZIByob+GV5LSUbkDz8RtQMdPB
GxSiLEl6HsuadO/7YViEz3AxpvBL244/EeWCVrIHkC/kBggFUNpS/r64iePzmRiGStR/aagCO2XD
u9msp/4MD+6VlTHnycyRiCG6z2aM97vhpE05nUXv/cWSKM+z1tWxGqV4Y1LobuQCxSaqpOHk6Ai1
IixVYW4g9NlHEM1q3xTC70eHDDULRRaGYHBdZTXaIm3qR514tjOHvQTQ6qORtt5kD6bcLjcgpP6P
ppq66xGfrV9Muoy6pqJN1lS9tkkh9kzSMct2tqmSv73Hju5z7VP1l6HyoED1OvenU3ySk6udHwqN
rBQRicaW++u7Keoae2Amz4Sl7mRBh9YSsNxJUOsIBZjq4vt7PyjxxCiNvf75HuB+pxVLRLbra6Oa
EaOkz6ggdar+Fulgmgn+lbVJ3/EEv/Rwz0m4CuewNXOnxi0lT0J7mNkvZhuS4y8xP88lUZtB0IKB
Ma1dSNIIgYhAmeP7VM3Uzz8LqMj2885l4AbYsV4hUJhWGiZzMh02/GFXR1J66nFnZXy29NyK0k7L
XseWA/mPwnEg7n3UHhDyQPvCPz0wb0iMUCODMk68WY6jTUShduuXNYHdfuYNy3WWHWXozrzoDDrS
0g3zf/NSG0N8hq2yf0FYa63k5UFA1qt23ymAB7R8wzr7ZWKlVaSlM/GYh5566VjsCLsp1I3Y4gPs
cNTCG7FN3M93SJ+G93xAZQvFQUiIseSueo7tUuDUgUrJyHy6udhA5TkuJ29WTEdKe6iXSENnW9rT
/H5+EAmv2W0tWskXDpjj2UhdqeEolWh6ddIPQU0KmdTZsX5OLHotjTJpzwIGg21Z6hXOVYtrQhc1
HCaFCxW9CZ18+A4ih7L7Yx/ltzzCm+OUJtM/UYSz2e7XHQgWd9Jasijt86YXboCPfUdrX/Qj1dgK
x5kMJDVDSSLz5LL62rZ9nPamuNLx2aYLVFxf9q/UIWn3LdgKepMX2ku4x+YxDKX4UIFPzwR9IevH
TQ3QLRB7R8B+jUNbqbn94yNhcLxOpB+cz4p3+KvpV3D+DBgPmnGM9EpBSc8kBIoxslxke/UF7erO
mNoLI7UyCHVCY4EPv8XLsAwB5EL+zfM7cmPBKUPqUzOHd+QCSEh5uHLo8e0XFfDASnlUT+Pyfz5O
JTaDI5NptsrE106mVJiZLCXLZ1ry6S9531Tvnuk9lRf28uaFG/d6kP9T+EnKILvxqX5pfFG154mz
zzUbX6jUw3Yb+I5HmBAIvGT8maXyGA6kpFSSy7jrKn3C+mBQPEShptuIm4VZ6m3kLbKkvwQexL2o
k2KJqRxOyUZ88kea6U1xjyQYJnUzsVIUPfe1N1iEHXPSx6HUU98otorD3sDtuDTWJB22Y6b8rfYU
x9nG3sDJfdqTX2F0phtdvOgun7VQhJsMaHaUIRNaVfAbf9OeWwa1pdNy7UNJLutmvJqq3/RUlatI
kUYLGmSr4K+keuqY1RmAc3c3K8rd+Jibjn2wK8FSHDwTWJbgvFqKqEHn+nC8Rux/q9jSE82HSMGI
F33yuTpo7qizfp5dZalv0u27Gz+XwbGS1/KGQgS1uilzv1akkd9WC/YTXBCtCnP27G3A0MWLGc9O
uFdJwHKkGzpphnpHU1jo7bOdQTaMpJQSftjKxJBqFqa1Uq+TZkFOOXW9Utjjhq+/zJiJDJ7VG8XH
ssTdo/egi1H1q3hegOQLOciEoH5sHPFg6H790q/OXSL7Az35RJ1w58LnHxA3dVamn4EShmkk/VPc
CbKEUpR/dlR36dlQpEs3ANqj9I1pbVqQyZEq/JiYYmS9lqea3UkDDh7xxV2XA8DCB15o7xOYm2Kg
fXNgTxqX0wkVXDLFeLEjz7BBHS3UeL4kYzXqowqPGXcbCvBx/NBGWNCF7KiDm+Taz0uMZpBgiznD
rcOPU4UCjCU74TO63RFu1lAcdYSosJLOv6kG3d5Xjg9KZj2J1y7/pnyIOUkV5k4VJ8G390SkumpC
4bUfBLhUbHeENqjBN2Qb892+vOvN0Av30Eg+GlqNADhm7+Sw5BBEMGYXwtgSN9mDu0lT6xq4EhE9
GlHd7svUKf+MHAXdwNN+vefFcGnDSvHK97GdkYtCuwU3L7/mFLco18Lrbv9VmondQeyQ52bq+odv
wN5UED4Dqia++pO2fPNlrrZNxvRPLCRoNTaGLOPaUgkU9otzGSNJ259mgTP9ZYgJkGddqM158a3Q
JV+L+5XOywt4rhgvyBHUAZK8qkNK/GXQynj1R0WbvrJIya8PQKmgZhLAhcNqFb1R7n6o64229EH1
IxXyjHj4Ec+3m439lMGJXGjRhuv/VQ4Ba8nb+68YKKLed5NqVAeSihyWNOD9+F6ZESz4PtCpngWK
t6bzXRvRin58kKiknQWQmYP7eOhk2qXWCTngX8B93Kzb5QJN+MuZY3FtUJQXXcARYlSj0N3OIRdC
9hMCYkHTCtrDoo9pQ27ucOiIJSSpAEMFybiDGK22lH+Mt91BFbS6BwAL0Y3+/EwHJqHyN8QNGnrE
oqGhlcgQGiy0EFDuIzqGAVeBGPqAVDqIYDdkI1uxDNU7D80K+S8WVxOY4G+v4ngt+NzciB0Dv+My
0uWz25rn+qrGrWzeVAzYfod/XbpVP8/cFvr6DkMcdDqK+1Q7AKmp73g0ZdKpfEKhNpvPX3oUZf3t
s1OtnH+xjiHBo1IzZSXNrxlRGtozgbWos8TdHi+19bNvnUSTe5/NZVkilM+O3tKqTyKQYu/8U+dt
oUwccld4d8ge+e5WKb9cZmqCii4klIpRKocIHWNtAtx90iR+IR8JZuCZ1LsEVzv0SkIYls0SdE5K
Iu+xe7rG8iMb1tk6VhMx9Q9lpDm6ZVdgpWD0tZ+tShIw1k0jJho8cATIiN338kSAc0IXIgfgteM3
OzUksBXJZcvDizEgmkXhLJOyiBomh0pVQqe9m9lWvqwUG07jbW6+EYUKrwysB6Cgcf2mmas1JN5k
lq/23NPWneNiPnqbBCgML45mEybQewpNcBEg2zhboiX9VBOcwt99aZSxlKL+jex3FQ1CWg3fWEot
jt5egUE/goIn2QnwMh4VHDDOj2thINRlXBKflvi0nWnVatVEDCD98aBJNsr1udwi6NtIgzOG7Xxl
50Hfa3NEebAJNZdnPfG3fJqDFz6zIGAWI5AuxUDirqaXrTlWkMtjgADfDX9wlK2KmpTJ5au8r2Sf
0mBIS1Wwfnypd/4uELLOCdO0vvhSt7Ssy/ChwLJ8zgZ2aibth4O4tKFJT3+fa2wfOF/YnJWqjC8n
YmfYV02MAWcjBp8rvI/v8TMYzd8JsvJ5fg+OqQwpj8wbWHrvuTevru/KSOhZ+PzCGS9+1CHkZLR+
kEbU4pc8MwNl5Js8qxfhCTX87OSmTHAKwx9ZPMN8sqyA2HUhGXnezcZjpTjttKfC/InWffbc/GIi
+JGuh0KSpHh7hM7h0YUR3FNRfOtfVNwwLObiEWDQbkS580bFbpYw0RZqpNZLzZb/TdoGfiC39l8a
L78UayATgBNCmgraL/2DSes7lzK81kXEVvYUzsfDvwrPK1XdVuRFAXrbygiDF/ZteEWNqQAIaHlr
bEgY+ofRIoshqGjGp0JlGzBe34j3JZpFe1xUP+xbzH3l7S4H9TEnXM9hsRZd1c2cMf0PSppbaexD
E1PFbn63iOGeIjxaEbHJYPB8yXBNqZV+Hz9YU/ZRdqDVOWDYM5xUCM8mQ9zoApD8VJHT69d/Bgqb
0/r2M2EH+TW+SdlqYPS8fIpkRwpJabWOy9Q9k0I7DqCQdmXlPCZcRCvGlR2LuedkBD3SHVXquXKk
c3HxdZWCjHCx6dcvB70VM87strx6mfx4dtBzS8CQTo179sVum86VhcGvNLfL2m1TXSLdIcDx8WQd
egaEOS+4zspdoSINviq4BJF+PFXnUYnDxknN12QKh4zQtKvmFCM4NsX0+hxG+93iG4UMsXd2CJHy
Snw5h9nfLR5WFG2VuI4yqXfWGLULOTJeaWGicP2LmwNYHyFWGt4NThAh0+T/r9oZ+pnh6o+dwoHT
aH6TjVTvAaXABVGHoSph6JVCDHUsowXtQOBSbGsjkPC+d40e9jzfXtPGgzOaidKauqR1NKGtLuad
UmMjVNpvC9zbr8wXy2EWBhKl974bgc9fXqpt2suSUgHvh9a8ew5oxou2OzhNo2IdQaEDgXBGDdC5
BmPEiwoqs8eBEwQu0l9o/3FHgCzS6XIJ8A1py2yfuXJmX4duANpeLysdjjGF2Zj2zUmcr8AmTrdn
SFRxaoOHOy3FxxCa0REgRPm69fXRDdlkj5nZsCUcTwYkSbNkqzCAcUtRRs66vyf0rrJ8v8Zb47IB
uEm8wB9JeD5UbRqSH3wuJ/2i6Ea4xf6BWPyRaRR6Hyl5raiYQmursw7oU15ccHAYPojRKPKvATXz
ePNBa2PBB9fx9QxfngSVPdKEUYabAeZmpupj7rKFHCEn5sxiicwURBDc78rx7YmBj9h8wLMVJ1II
EGdJt7uMZSkmvqoy+uxJS5vXefhvhHa/YK4bSeIJbyG33gn7+x/nbGOY6RNyT1RRv7W2jSvGDUob
VRIDUS5KmDnWfkKAcuocqQMrCDmXMY17XQ3GDQCeI5VvxB6TUwWog8uDoIKHseZWp0xzVEaUd1EQ
lEsejqJESw8eTg340gGBqq3gnmvIhTltcq0QvSOuJ0cbA587qcbH9Vd5Hkkhzt1JlOoWEsU72qzf
/NKv6iKTMzFOBtA9wex2fdLu75YvIMMFgU0FMqt43DAUi8k+mg6q5NaGBM7u1A6IzXf5h4WF60tD
c9vvrtxxi2SWRVHCpJEjWd4D4Fv1B31YlkXZD7fquRBfSZ0TdxWz/DuQv3nE+NoMv59j7Iad5a4O
21AHucrzrWY4QnfjdT3iPm7sD77ODS8q+qZmG31SfKF7iDSGKKf5RNyxud/F+HJ7KyQ4Y5lwQHDN
3uwaXYsI+czIGd+ZgF2dOzRNkObrh5SOqpD1gBgmbK0DlwzXm0uCezDwAC3RPVF9TAJN1Mp5knHg
rqIC4/u7UEtuGdH5/rMJ09VUsRVGFVPY3QZUICPTvdqnjyisFvsuGKtnE8bX4bzjOzl/RJAhwMCm
fii1gc5gimNSsEWkahDiySnTrkdK5gNOAz7Ym7fkKxhTmzJ80AO4oYg2oZVbSxMj3G9Elwe8VCR4
reAB4ya8GT1JmEa9KVi/AGhJR1BdzwsrILCZLzY1srDQ7EH4T1e8XQPdcZsIfIEni82ghw+j3AVR
QF0VIj3JkJmjwLUckgA158od03ITMNTYQNfSVHi4ES8fkz71t9Ey+NkuZuSObvsDPf31f+HMbtDp
iUT6MGjxFAtbzPsmep5TBawpMF2XjeEIP3TNpOj161G8nOiW/wqeFC6UOr2uFniMiMhfnoKKDF7D
PslrPuqJJoLwDDUBHKQK0hocMT3JYq8BD5LJO0e4HmzB/NpoT6KLQVhw/ZrE+G2c2TktU5rWFSCj
R8Mjd8JQua/6JTLFpbGcctKUV1pkYdNaHNpCuq5F8nj2ZZ5G6ZqZ0W7xsZCFCq7+Ey4O9eVNKWW6
hJ497ZxdRfxMCOA4R4bT/71pH+IPfZk8YnFDJjwExx/eSZJZwNCxtKEwWJ9EuXCRSmvE+NFttGDe
+bRsrIxbOObVAx0eHtSP3dmn9MmZnUBr/CYRgW/8ZIlOLa8gZPREswT0a5yPpfduOlsOgRfMZnx0
ppfVoc6uufjJmMK4pz29T8Upu/wVnm/6bL6sx3bJipfEgc7rFJTwfKaPpJpRJ8Whd4GKDCFn5tqm
arVBrHr5eu29/w+lCASd4SvOCn288LhnPDuMwP9G8U10puEmaywQ45GtdLuvPDWkaY54/kq+4JuV
6xP0AGtjhmpBpYulDk3M5lt2bmHxOD4iX2T3XGrS+HsdNFZSXeih4bUBKTi83GjlRb55z7KeUALb
aG47rFt8avl3DVzKOrpfLK5JZNZLP1Sx/7ts/CPgNFnS9+IWiDBDThiKACIme5BgSNjAv0d9Etuf
FpJawg1Oo/d5IzUS0wv1lsLIgkq/SV79rWQvO5rZYJqROVSIpCRecwabbYF44vaqTNm4Aw41GCT8
d4s5Ca4dRoXNttNjHj1h8dqhgsS3K/TRnKbemEjQIpCeN4I2hni78KC3SFSEqr9oqAip9qxzzWEI
+LN7JDiOw/HkQzbRufWbUFU+xHSO+s8nVm9x/r9AevWnv5S+dBds/pWbypHD3U+N7EnlcXmClJZK
JVxHZOHaZu4q31UHDNW+GnG7K5faOJjJASwk8z9R5PhKC8NvqoKJbbjcAoSfGFJqaTRAGEAbLGLQ
T7OXjIOget+nFY/6Mdg7eGGdN6jNASlmziKIBom+m0gxl7aB/lWNNiZVtKxfg+zB/TYQOyY2BECj
bAExa/oKMuzZSE85d5wL+YARWKzUVz47DPkBf1mpsihC8eEopfH2xBeYoxw4rdCY8FWtEYVeqo3w
9/xKXyaiM6USI2hMJGMShM8zL9s+B5Xiis+io0dkSGJpMFGYK1NScQYdC6/w3MpSvzLyk0Y/B3QK
7lluEggv254Fc73hksEMSjkBPzjqUTYMryX96U4QvEFSneNuSC7Jrs2PPrBtLZp53undnyCH4Sd3
JHiGudMM3WvvsTRiJN5HytzRmnUYNaNTIxEtn0WmSGp644Qg7e/2vMedU15m6G5CQEWh8GhD2shy
EQcW8CVIG95V2WQq4RGb0DErwOpJsiO2bIqoBaMiQXSougTwEKb6H7thnICe6VrnZFYn6iTkdrBa
W8nSXxSA7YaEqC5hvgAeRVz5yIJygZjV7p6UMyuGWkJFEPWlo/98LXNRvPVTUdWaqlTrpJTG3T5r
5kiUF0FnD/WXuZwE0Z9zfZHrZrFmpCgCgYpEA0Aef5XlHlPkbuISecA/HUkcg2Xy4dH5kMxb2iDk
JK473d/BAIQ3MvJsgyZxOhR6q0r3RCRtVI6SdrELGcrPck+P8yDNzf26xmF7Yfh9Dd4YSx0kNG+l
776m7W7tQL/ix4wZ0AbZXnKHf0YNiki5CiJDgK6uPDIKlijTBwkuyEX08bdeOzBXG/Xs3qQqdZmE
KyV3cblNKoA0vaEWdoXlZ4Xo+Hn8hp3x/HcIbiVTlFIG4kWwcw96iNh5EKMGpXKSX3W8F4YoVT6E
8Wq7+2TqvS278n7+0SC1JPrP3J2kX+JNTm0eVZ91hjfiFj1fqoVgzXUaeltAukEuLGxUhmz5jiT2
7Pu3Qbcrf0K+uapqGdbfdhAUBVDw7ioVOKjbkZ1sApqq4WDJBB1OdWxtx33+DWTFI+zLKaivPp2+
NALqn/EXEuJWjBf3o0QHXw9dW7Gal92WZ4Zp6SHD0zQRyo2ZzTViJBkPixHJNAlELX6jlrSalNwQ
MF5DSIwkuvOUpXOfx7szVUzwPy9jwfB/7r/NHrzbRQzYNJUdHa8+9JGHC+fJZRddeBVF3D+CuKay
V6l4ujZZUi63vHBQuISxWer+MHt/obz5OateApAtJg8Bhok5turbN9HGu7feWtpNQLmIX83o5alN
QFjAbS5PwB4rF3FCinGMJEzxCCW4Bj2cXhdRaVM2VTPXEaBXw0u4Dp3faYvZPv8fOlXyz9xLpbAP
NsbVuS3O5sWCY8Y8nLFMy4+LATF2WsLXGPH1lycRBs0/db7l6SenS9PT/JRmcC0ZgclJLWdMqiXP
OOFl1sHm5Ot7eexq6EsK/zq9/AKgZ4mI+c/hs/4ZQn7wEQk72A8Js2VQFgPoiyrEWJD290w2u+n2
Sg83VQntk1Gg+jyXLJAdGhSpt+6OJurhQE+aqKjBBeHs92IUpLOKdoiLoQMhHKlq9rfQFnqmReRY
LwUJ3mI4ulIva0KUBGaeJxno6N2K/9bsNhJF7CuaA7ap5lnCO3ye/a6XfjtyvZm1yL4QtefX2HEj
124Ql2Mgbsz0dvKzbkZsXF5wnQfvGHH0lqPg/oug3mkmdK66/bV6z2xcotoDE7XCB8ms6cdkXXwV
ysqrc3Vvwx/2jz+T84ZI/v+LDSTiLGt8aYMCmPgh9i0P81L6ab9AB6YkKZma759woXHi9p4v6AOZ
4p6/pJ0YOaPT3lb0Ym9npv2gGNe775O/1bcnr5609XvUoYVDl3xA279h9976ZrqHCuhbbvxdYmJT
CQkvZxne77SQ8xIvXma9bBQFpL0oRtDpom0XVVpK0TV2J7iY1QHIfCmYTxYgyAZXIRjbnzKFTllr
gjCVmxQqSbA1wjB5Mh9313P31HCRQ1i/69vpydWpPJ5Qu2DAiVijunt5BIWFW2todpbSMaPJvIuR
gAcrvVoMnykRO8nRPKor1BkRC8Mbsf8Q7IVcA/830l2LdL6PT/k8sb06AkBgDzopxBVBeXp4vQDW
Q05dSpif4CUaJBVhCIW4VPKV/mbhHsRkl8ZtWkpaIZB4uUdanWv3HMEgiKTZBfMdziJUdfSqYhT0
vqD+AZDOAa12b0h9CQ6nGLfaGoJC/hpGjDImMAiEhfXfvThf9Kq/+wRuRyARPE1Egd77h11v0v+H
h22W4WBqTJlfOKruGBfqNOBjVAXgw6wndatyNNuFZy8FiIJyeAMdlErGf1VDNT9r4lM6GJoxO37r
UaEgURSX5KRfKUcpj2F1zc9xnw5M94JzW956zxLp6qzzXpVsuBg4h5MBZOUicvQ858nz5+tc34qV
ts4pqK3Ju6Xk9Paynww8JVmQPRx3KI/ZFjIsgEK3Y8lcJRqLG50ucyiRcAAnou54STSzD/ibGrTY
74DpgR/mao9WL16vgHfAZIxAZRzg5qcyoKoNHFDU/3hBrAZZsW0aLMesyQIvX4FBKoqMFCtQ7SLH
t/dT2/FhRxiTR0CgpbvPU6s622TBXF3syXIEqxdoEO91v7q0rsB+e3/pSwz2fDGxnNx7RDSc3atv
6SE3izf355wCMyxtEJLjIBQNRVdYBu4LoTvSxdsBWRg9ETjqF2QrjHpCAEfMix1PjJ7Hjffpds4G
vIGmWx5jPaDcV2N8AYmaW4p2f/Nw2lRLa6nD8rju5QbZFh8QGRwZ5BTuLoMrWqZfBTRaIyhf0vkD
/RrrXXgSaz9nwqbg5RXUfP8dEouZBGYiyFh74Jse/qRLijaYi4eejss9FRD+VG5mXf6gAw1VULZi
9G/VIqJJmmfZ3Pr4Y4Gh+ce4Yp9D8F4FPYlLh27oFolEmcLozAkDfmCLkBGdyge7ao77TrF/6pbd
I2PDHv8dXYF/5PEPUHCF6cIAn9XC5dX9PdfjWNddpE1tkY4LXVpRd4VKicrMSY8WKRq06wzwr4hO
k82JFd8a/eNTfD2jWfWs11iVMeeQDp+aw6lv7eCyQOY08ZYmkxV2gwFGxNvw15tMa89N+Z+c9INr
nuZJeXGxgEJ+Fov4e0Yt57oyzMAX1vyKXapOCBPaGyROIHp88oe/7C0xrnsD4UGSfF9BlneXx2Jv
CSxM/ipp6RNH4VhGFTKPGUVASn6lRQzagO9G3MvPW+8j/1N6DNFcRln9AdkouVpNcTqlwt42Lpg4
jDij/hloqnBO81VIBL+Pdvbf9jG0XB58okYgTiMuAb42VE2iEQS7zth86f3AQKPGP4iBC1aU8hex
vlvGpiTAA7yo7GOzYd4W05csCNTWglI7U8EBynS8xhwYmd9IX6OWjln6RdJpQ/xWYO5jTXuRsXN4
LIvh2UnqMc2ZAIRO3duwYRSQMNJ6krl6QJ8jeS8o7FkwzC7Qos2C2rLcTjo/oYNVcj6K1vm0sxYy
FW23Iutz9Urm3k/cwN2ISvfwAg0EZyzxnEk7UDrFZ6ArUrtlctk0Kc09WLGfAmMcXeGDPayoyZaF
Qbn3it8n/Y/9N8WRAvpLAhRi3IOrSlZ4HbJvVSBVIQrDCJ+rrhkqxkL8WdGHfn68BzdXYUUN1fK/
Bb0T+t63q1A22SPh5e5cmRJvfSFzbGXxuqum7HxwOmADPImZp1k1z1AVHbQJefR5aphcLnxubi/v
V6Sbdf6Ns1WE1BD8acsNz84VHfA0n+hsCCwszV2LQk+sY2X7OFmGS1aUwekd1mWhSSJOoGszdBqt
reBz/wzJuqXEYijBKam4f4tJ8zAnzZNId0HnAgLD1GGkN5JXV8VP+fa1d6xyM+HTUd2ocFIDUmwB
ebWgeiBZyr5lWj4bcSswOpzIWWh2dPsKC1166i4UUvszDMGSaqUcwtKs2mFmK+11KM+0eLADC16S
wzQbyQ/DIRWbkw92m1qkaKasqC4ahIsJ6TUC6NUvxFvhakaV2aUpDZm67seQ4qrCQ6FvO3Vus9rM
Y+stNfL9eY49c5xVwm910eJPOYTeFvGrIPjfwaUL2f3d8pxM4I2q/NAUgfE4+OuqDbnSTyzhR5UQ
Dcr5IGKlz7VJPqo5liiZ5CyLKjLxP7vm/g4SyFN2MD2uD5AvOAh3HGN4rHdZQwY+y/Cu7m09GRlO
64fZjz42vvMpZPXstAUv4LGvvN0IORpBsBrwyfd7e94FE/H7yjFCvB6RJ4GUMmnEqavE4einTMhB
Nq/02RvJIS0bbDlAkf1+rLSzyA+ch9Zw0nI/41vYislkjThYSmI8sT+yrKFA/3LKF3gF+CU4V3eJ
rR1w5R1su/ptuWstn5Ru3m+FhXObo/GE5GgL8RRCoxabJx4BFg1sQra4RrMTIlHEvs2DB1lLsnHs
XBN/1RBpH3l1+LoRHDODuPCWlfuWBG4smW6plew+Jf0vPS/SpWRstaOJMidf9IDMXVWVQEofq1zB
jzN1MVCHEfwnqElwPXY5YBwQGfNeE3NOFyYb8XrVbu+/1ap0N2gGUUefyiZc6U11bJFT8hBhfhPF
QZ7RMN9oDWpAtoGrEvuMTCcz7Vfr6jj4qUoKj3DsTI4VCgdrkR8/xS26GJxRUUDhdMdLcSuV4mjc
LimL5oAzVRj17iAE6xcvA3oYhh37M8q2gMWlsplsOz87qxtGhtKM0wR4nGWGI2EICGaiqMA8N1cd
eJdxXdwJJXEDq+OyMjrfC40W6rmpNDk7B65trlCAg/lCSoyZGO2wIeUu+31WaR6fGjd7zdYbnW3K
1obrrgWXldfUtyHpeYXenpHPuU4XivIJ+MTpOW0TUZKM583V8Xx8QAWL+sNRqsVgzA1PyN6NQzOo
GdfqKGrVm6M2gE6HP34wEv9B1rJDQPRjNTlsHVw25tRazy5qIWu0vTrYJg9qWzlTtNW8qiP9yhLx
dY8+QOyz1ZdoATUXho+A3G3DPIyn9bdUpmiPCfD7WbiDCX4pqLhtyw7Sk4AhOC7cC70XnWSGh3lJ
MRHFFrrYvrJpegO+nH7WX0Vgprb+EcWnHnFJgp/P5UeaS/T2nadwX1adg18EVbEVAayDWn9ZQPMS
GBHzbdid/F3mrA4jbVtRpzIBM4rM3AXdQ2kLKAPETE2RMGkjqlXtxGV9H9+4QnNDCV7LFIiTXAgG
yTw2iILN7mlzeciPDeWvaWZ5LIzKI8ssu7oPCjXzLQAWQTfGbdCIarQGv2vwEndfXmtoHBYhxcQp
konlQJrjpPjnR4l6l2z5m5FqouLF7fMh0yqxFP/4b9BWJRSz7bCoxx/eCdXnjiGwm17stNdOLtkm
ktzGub9tuUgGjF9eDOu8tM5V7rZ85IdkCh2bszJkCk8WRD2591aF1jXFTeZl+riCN33ckhUFYJny
GVXZTgb0RhhFuQqBZMNzg1FVn1asDmINUsYo39WKHnvQudQBf045kWNwnsWXgO30vp4BOuQogox3
PP0UgvVdCxSER64yB+7zvnCAzgjYKAWwDXmZfKfS+ovkLLjXfwT3lMS6d6beAMMKxVOR9xTQ2CXc
qs7QQeYzqeg5ZECfQ81uDYu8F+YKNW5M+m9CUvM9fpNKPdXVjEu3fieSo6bSF5wjGHlC68icof5/
SaP/kVP3R7hk+vnSpf2O5bTFdJfJmmyLyPVCqI7N2u6EjreGv3Mkx5XXUbr2+u+5EyY1UG55S8xV
lhEYOSjnfy3uGuwga24VNKF1GZco9qYvnEwy9j9Iaer7lkDbFB1p/M2x4cnrsHIlDMP+kwfmaC9J
qMFDVFvX3Rkuu85r2D7oBFs7fk2kA7fWRFumSVun2uH4DpRjj56E01KdAcOVJy8uwDlTvKWQA4dD
5m4qXnoF06uj28XFb2Fe4Z8myKBTdnsohL9HMmpPHzN+ZvfmiUjnVgZSE/DF2H84pEVe9a+dnBbX
XSFWd+PPpBPA3QXEyB5bWFkNcTRI10OlRy/JRR42VSjcyPJUUoJLuvkhq+CU+GNWFz0j82jdACbM
kekiPcBGfsskyiX8FALB0abx25M4y1ee6eCTMbgXmSuDNMhZ4cs1/GmYnwNBV0miNqf2PxgCC7Io
fHfSHMkKaQ0AUKI17nSoHsiuq7eWx1nTRQX48fzz+HEUbcMd3Rw9pFc3XcjkQyoxzdLYgDef+SSG
1pVqUvZVEtSfKBGYuAouU5IiZ+82qXrEfXruCeiQI3OA+lxjjcSR0FBPQGp7vBCA7DnXaQC5rXY2
BDSYLI8QokvMCA5eywIENayuXc+WdkGbrDmMNEWvwfB8UE/sJa97KBKE0Solrf4b7vM0hcZ2w3bh
j2hl/4p8rnS4TGVkwLUCIbEHP9X3Ughj557YKpcriZ2nPtXJkm8tZAcetpFiOF0DureK9sMQfpHw
f1yoo0Sa4GkRhG8bHIwMClcJFM+ClnJVfZQ9jTHBzAmNC7Y1RY0GuFzjo6ddxLu1UAJerQ2aAQrc
mofpFIUqzb22eki/dVdvnDgP7Xr7vX3fwtnw4B24wM5UknqMIwX8HUe8icmuo0NixHpMbD2dYKDs
37PhatvMF7S7IGr1UNAlOB3cEOlMqRfRW19NZW2FQ/9aB3kgL75RQ91QisciNgLZXWjS+s7mq7wm
ZyBeZCWwOWJ4yMBDLTmEOdNDY+VhYWd9UE6j0DYy+efK33Ulxifi5ThNrgF4RnSbIIpFaviRKj78
uobcnsmlPhi0VeksfxstdpF/NRDGVS/sAp680VFLVAdBXlMU/hioXbtBvRlNzpBcjUw9pWheG8OD
6H7+kYunxsEnh0ONLTJytUIMLqSXS1m8H10x+qIB2qpuMTJHZULoK6+R79fu4OQ1vRR7cE/NRViX
KB5de8bI3qxZ+n7cuJ5mrhpUNJtmCLRrKSavxpsCZOqGVVbK/SdmYpWDyTuJ2nChtVHelhN0tzM5
FsvByOyLTzZL/hpuwI7SOs5AJ5Y84K4XraTAvwDb1Tup01N26QIHdGx0DCd2jGKCf+CImRAG1GyF
AQbACUXXE0iP2y1IXy9c+dQEXjQBf14vOpBWehTVqqY1ctcExlP9wkLNtPhx1Sk8E/KHPmMZtXU7
vcympUytUUUeMa1tAM1fKsYr+m/AmP/ZZw8yqmpUC4x/cql8p5NjTVlFRkMZqFkd1q6kfBszxYdQ
M7kYeoZF7dv1NFVHl+s7MCdeVbiHBUNPlVZLY8/hLSKNe8LJSF/Dd6n1kYS2eDdGyegvmH+aD7z0
cu0DRBErsW1kQwPRrLZv0aU5NphqaCKZlF8bdTmGCJQjCY4szDzMMtAUXcrYfT4l9nlh6+Umq7Hu
APQxqcynS9zIAZbLapWmpjzn+q4rJuSvvuweStgbDD+ntrtEOg450J5Ch3zoXGfI1DwZJQGrfJEx
SuojtLw8xI9KXxE4UDVI0I9DO6NFyq4D4jfV7K3LMEpbmrynZSKKfpIATn/FMHoXHXQtV+RlA/tI
kv1QdTtHfEYvmV0dlN7fcbwz4We0WQzVfMbag+CwPI6wVN+BdgI/gyXndR3kNiKsGuQmIW0FniUh
UAL1CmAf1i2rAMq4n1sl+murb7eNsLkYKmVQZAy/c6WYbeyfD+Yu7eTn90qy22Kt96ujE6lqTgi4
WayEBWuTbXNMLMPSkjj+XZscvODl40j5HqBLH57UdckRnB5aAp10CVjLUyaaKgq+XD9pTaUWgItX
udJ042WEHwfNVO0LEuQosedQM4rFTL3foR99uZFudr0rsOP2LFDMRuuiS4SYGjm4FZ5tw7G6fP7b
Ng6f5g8YGzcGFe3pOLoCbT6dhDDaMGP+7iJO42WsxXelm3KOM9V0R0OXjhaGz/aWI8wCaya/3Ntz
k8nRa8sS6vZZgSgMIarHD4olp/8LiVJGuWRFdnDT7MM2CdFeKl/wP2u0TcjuebLTpY7cei0hYS2t
ueHMjFOMpx0jr27c+bWhBZMgs6aQ+RGrOwG9p35O97aflnXbuquDDkkADFIwX2xEXCtO0uko4d2W
zuB54kjzuTEuTXeJmml6MHUe7StCBs9DCERlk8b0mLFriR/U2Raiwg/9hbmghG+BXqLUkbxbasjt
T4r6vVVhQp0hPIosp/W5Rhjd2ZaqDFR0z2DNKj5jbmbGowbYpxPANGRwGeTE4Odl+J9aRMtnoxw7
LglYSvnQcBiQb79xaflUDJixM0sCwxSHGfTXCzfbMLJs6bvNxkbsXXMyHZEmgTHt5x+SxGXjs2pE
5IPDhdqcspEzCCD8UogXgPDWJ6ss3NwhB3xIu75LKtYIlnbSa3eL78TFZNwY78MB3Y0+WbZm6IAo
OQlgK8LGA4vTkW7FnxFQryAmI6oemNGTglqf6dh0fu/3nhN50FzxZe0c6JxlzVRIUEFhGyfJNVyL
esp9jkWJkvae1kGWAiSojvgQ4x3/CVLk1E0/F7fha78dCqA3v9JlmVF3fBie4LwaDB+Vkl3Dqrui
SYbZKqDMXQOvtaZ+tZHJYIFcl0EwAuEpuUhPCCWqnAQG2zvsQGuczpwTbqa1YsOg3hdnM7Udors8
AXbQZENmM8zncA2xbrmFouDRhzOadXIb2sLnotNM1JGvfpuwoGlQwBiH8aiyEW5gkIOsDVOw/VEf
UdqSPo8mYVhFLXLdNyK88qmfENkYNBLTqPc5AejPxfm4PCcY6Ac6OnjusEJmjDWzoCM9yY//1RrO
Oj8RUR5+fY2oe10CdtCR9oTqO/Alt8NT1XY5zcdpEgzahbPtCHuAJ/ppKi/qAaek+Hvsbs2o90AS
ART3g+czuQYBINnCXm8RLkHgVLLUMtMAD4hb57A+f5bqKmDHWue4rbJp3NC8hKGrkZ0R5oHmy6IW
Iw39G2J8QL+mvxmLrvslMjs6YHtTqjx1qp4YWKuKPcAkDTr/dzc1IkYwdTsmCLPgQmQJQUslnHgl
ExtLwkMZJM1nW6ydQdSHFMtZVF1A5zNDqYNIECMQwhN+pc7klYlYc029ST8nA3XTxZptovj+Q6y6
M8nT83rltvl7FKpoKTgbuQGTrn8U8P+bYvB8b+/PODl2EgnFHG2XTIxy7KABp12WddYIaHuHFggd
H/r8QFlmSxsqc5KJSaobSc8HGWzpV0A1kGsaI0wnu8WaIt9kHeVKbExzd6WNo2cZjRz1Th67ixUm
gxXgKcBY6egaSDPBYGTdQrH5qk9woQwR/oKfwvLntLF3rZwV859e10n47Ujsq9dhyaJjZPfldX10
wJ222nKKYZFwmeZ/Nv2IMd4rnuoM1ggVurRmON29S5DOgcCDt666b76S+o7Yyz8tfGQrbq7It8+L
QraTElewYbuGSuN9c6IEdk8lsjh5Iq536MrwPhOertSEqwB9yp8OMqyIaVc22R7E1RobRfpd0JlS
BOQgknvLOBKLq/xsMKb5c6CDHEfF6+yRzE9+VQkBQjza4yCHiItZYW3XVOGMKx2hQmzDk9dbEh6j
9g1R6WcKBvZy9ep7t6KD8t/DEyBIllvIchUIqe2tLrrCdAnIqdUvfLDJu3LPcPXEadHWYien+jUR
s7WOK3QAUxReW7VrFs+kb07pare8Zi5sk8y+W4jrQz/CpxkZwDZH4hb3gq08Ng5gCGcIrgWY3ayx
3bYTIdeJo+HZofh6F5Sjz05SBUU+9w62N2zDyZxoyvp1XVFe7pwoFctuQehnHdG5/WidH/7/IE4L
VQ8l/RBiewV91fNRWK3BPhzGELY45xJ96il1wR7F7r9molZbglkFTFmE2rRGxIqUvbL6pIIeFP+P
VooJnRtnDL3jt31NH44H8crsAglpJcjSjf3AQcVar26XOmbJlfz+URcaa8/+N36OcjiTdZzNm0Nk
etFpyVVUelUyrARa1ZVXkK5icQmt1UF6R8TQG1PGNYXKFJyIHMPIdhnf9xqCo9//6oh/B/h5ccCH
inj0b8LFgHIF9PWd1+HPN5AfcBQw9TMvDNvbD7detmLi3e67niNBcYvCUdO+YiDBfljSbFdDBJM9
YynPtEs/PCX1gLEZA7G8BN9qaxOi6qYItOB4pZJd3GhcFF+LfgmsnT/MS52xKpAqOOlzkA5P3p56
v25oR3d0r74vhJzhIcoSvRnRr1dKcwBskaZEwoiaNn+Jy7p1yN7KS5eK+WrtJ3v5sLzRNwi9SIvK
/pcLpf1RUx4HjtWMHw1P0TgpwfdFD38Kkli6+qcVTOzvedtegZNX/1f0FPkv674P3zInJYf2JWbb
4glJrju63YIv3dywk7gcU4S9IEOQUvxbVRnL927xfXATUvX/Mt0lXmDb1t/LJZPjwkhV9OGdd2vC
70J3zO3Nqb6CYxAli29OfntlJy6e7VlnopZJskgm178yyPj98Mf/6z3R13jIFP5fz9km0hqM41O2
5ZRcsc2Kwb72Im3M6IExtg9X+q8RazpQl1PxsZ30jZ9f0z8BhJ2hfeGh48tl+v9eo3edd+tX+Yjf
CjelPVoWvINzLdAWATt4t/h5j6FVnUcbmr5OaLemCZYy2rfbc0fvzX1YdPEc13zbNG/v7N0L8+f2
o0ltSXxa5U1Kqx5hDdRvYS6RzNKjwUyDj9Ww5qQyvKhCyOphQKH5daiGzjN38HJw3b+QCRDWqO8D
AIXYkI4TdffJk8QAR1VE/nZ0sE5z9WM4rlKNiRuJqGfSzz9egiCRIbe7rKu/arWNzlJTWrJqqcL2
FqTXSmV+QTLH4t6OPz8e/lMH8xqmv2M1yATT+t3C0fckfsJ6MlampF1SYcUdOadtjwoU7S2/KZpe
8XCCHZPwU6uEBPV1NYQ7IASwzxuUsUVDlF9BJjKP9krOEkExgaPAGnlV3wfX/bbVrX24hmDb0TbG
N8sqkYAPc2W6s4B8JaS/JJmeMWpqVF3quKO0tkQynVN9i3JnWsLfFN5OT1y0ohQiPYMpwoEUG/je
/Ot9rcOKk9JBXvKJaIDV8OcD7lQ+MWYbBh7B9dK8MGygINy0gvNB9zcNcGwk/FXhvl01Bp9KmTC2
mQicTTEN3u5+ZyZv2IYudvfBMkiTRSWspRbruCqW9eA/BJMNImgL6Ad/lOkdJCHt7Epv/2qVtThK
kr+3HdiLCWFmgIBSrlEYb9nOjVs+ipwiwWHBnf8aNR0Av+/tyj09D9fH6jJ+iwXtFqukCpFM4w0n
N3RTg9oi4k3gaFkCIF50mVsT7fQITTGIgDX//ll5xDb1iUF/k4ccFjANSca1g9AnRjs4uOQnjXDH
FGFl94zi07kMB2OvxJf0DxMpKer8g4NP5xKolrWDTrD7uEs+BBOVbJ/fZ1DAJn17PltoRA1VZyCW
42uj+mV9rl3tOs4gT0zYocgpPBOi68DL8gyCUyLY4OCxd9pd/KL8GRc0jYL9TXTWQNn2qHEBb2DK
jkBgVDvKPM9z8vKiBE1KrSWBxj9ziaVRFz97SVqj6XMXk8HDI+T9sBL1minwyC+k8P7iZO595HRN
s5OKnbaoVmi3cgl3G5hCdMjtTlo0M8swNYUcKqBbdUpPvOWLrA0dYjYFCpxYPme/bE4qmxTtG2WU
hDht4YVzV2GFDCAdIk/cWxyc0UPK0OdBFhD2vahRElixoa7xfQu6xN1y2GR9NA3hfR7r2xxB+5Y3
pB2VF59yoFZcosVe7QybDbXa+0WnbCWXgH0Cwgw1kKxqBx5XLbOlac1qiIGVbjMIms0OdEuUAYRl
ERlgzuPDhu0Au0sdJIIoaezj1IXhDK0Z2zLIPlnn5Bphv/1vdvppW49UerExHJ+olfGVmI06SU9X
OSdowxIhbHCTqrqlYQMTZTQe/I+O5FwdRzFlkxNqEHIzC5Lvo3SsqvureQqbYZDafNSDqZRpZc5R
RvDSxKhQyAvxm5uS2rbM5ZRDnl00c9XRHld1nAPBkUTM9acfxRT9Dyy+aQqtXxq2GmPgz59ReYAg
MpwkarbGmZYItXTnowP5X0pshgSvVq36E/419V0FoSN1mCGHHAREgJC9H91XI/aS7gIiJe2Iz/sP
oSVlHvhlsMtpTR9cd6KDcLWhKkOZ+TpngOoHErBGJnYhlviM3WjZnmvzfXNq3QPPPQUWi8HYKLZJ
i4HFE0FdhgmU6iIpgdLKDK52cEwdlyNYL4WXLj2u+mp/kKRFs9UQoSwX/pxTaJlBNS6svaPkdxdX
nNGpCip0LwaYMUTc90Va6pB5rAQP09aYJxLRUYFPDDF0kXyhzj/zt20Rz6ZPGATjbAfF7IVqm9F0
EkysIoXftJNGGbNsgm7ZRJoUSc/XY4SVX+2DiLfkzBu++5e+1iA0TaIIs8m582/Et+GKQ/BA9+EY
gtPe1OWu5F6fupaqHSe+4NxVCdK2m6ZdEzJkmNn9LF0UgibujWTQxRk7QgE2/rgs1NZvhMv7NyQR
lXavXY+wO9Ak6GHh7cDjaxHiKg579vC8VAmfW2LgBQthJYK9iY3zBJyPQXRPW+dMHIIQNx/zDRK1
OQ5PeX6vhNWhk/zzkMzmFhPbZ9djGplY4UKizWAdtrw3tO7bsXZrNDToV9N2LXfb960ZTxiMH6A9
SB6C5OGMabSVCSIrOlanHtN3ZCx5S+HOjX+mKdnUzMOF9ll5LPxcQNaQQnyDgc/sjrTPfyrqxvP/
cQoYxVSwDDc2zKeZaFL9caht5fkjVokv0uv1FFBSGzUA5cxrRZLmsVn/Kp+LcVA0jfil+fq9mj9k
v5GMHe6zj5J92smuAR3Rv9Cq8e5kJjz2ADKDA1k95OkroTTaw/cRfcXdejnjNVnuKJd0VIULnGer
NvLk0nxc22UMq52fIFP2jO+fWhduVYn1bBLv5O4U6g2PhcOCHNkHcoEKRAPc/aMWFioxfdiHYgda
14SM00m2pvS7u9dF/LgOm/ghH+/8y4RIguf287FWjsyYjjWfoy7RqHgNa6ycC1Yd8gJqSwAlupPf
Sq93nu6Cb87RcGGJcI/iYQnmOizeS6cbtha0PtFgGi8P2oUz3+LJMOPo4pGHWe31S6RMXoJA0D00
B9mydyY2wCDSX5lBWuDD2E/95eT6Ub02xssX9VhUh6sNphqFYSAWFJGXQMggmbqqKHoXQPV7G3qo
50RyGeEz3ZSIYSA+iL/4xT85gsGJv4MLwAdO0E2HCC1Ia78BGsVOBkK2/viNB5fI3ndk8tHnPzw9
S/6KBYwZaZDWo2P99RSTTpx9g1tdz6fadn37CXQpwt/9nAe8fg1TuDyzk8425jxCnzzV1wHrSauh
nhe3JjdgCIcsIOZldxe5B1e47ls51/7bjvhc2E1JTpcIzdIZpfff5Lq+eD1hAhQbmE9XvdOrGSW/
wNDozNm6Z0ky7qKZVwWxjecy+/L8ocAavCDcnVDoIYuc26p+kxUEHdXnLGZ6KxP21th41h3WdKoT
vG2C/puTsH74wkVUfJkc/pi+bQG6u7jlAbWdggwuVaUZFGDLebSrThJLCs/1deDzEYjuDlYgZO+W
tvkQ8xqPqFjcjM+i5a/lDsRhB6sQ4oy6jHW682F9AqWOmPZriBm9JmvA2ayJiCxH+wLTFg4bzqME
XJioHtQGLgOUAd1qAzzJEPFcbMLq6Pa9QiNh5Gcc6G07XJelkJJFXRtRxKu0A70L7C1keXog8ERj
KQXyAZC9m4W7uVedW5ZjnCdODaJgaPT1P+viXc0nZgLmcK6LXxsrdfZQ5ahpihNWymM7KaZ/9hCF
EH0teQtFrlUY2CseBlOR3t4HUBkb+g47Xy9+fQYHVGlV0hGbDDuv9lLsdmXYtPq0HiTKOE+BZCJr
fC4gby9j+3ipXsznuosMYykjo21rHc8LhuKuc1AxVo3pikDzJ/1ae/cMiJ51XoJ6b7p3RlsJUVuU
SaFwjj4M6YTudjGR4GcuIMB7T/rlMD186tgeTjN/GJUcdvEtUiDMdwn2aKW96jvbvBUsk96O7Pvs
wQZYla0jOn/kkDUBR/Imi1AiGFeusd8/nELwvUib8i3aCIHfJSrUBxF8CZBoo9nW+siArmJsGNIN
Pq9+n4x8xQF2P8FxD0l9p9wDDBToPmAhl2SMmNqCq6ndqMG04by4Talx/67Ak9Om7+ub/kkOHE8v
NQjGXWXdTpBBjmGW7Jml1vzfLX/DZhGCMyVO9h5U70H+Hi30NRy3ha906PnbYDB3/cfVD25WlBAx
zNZCU2ebU0PNWly4aWbWVOXq50IFXXGq8PFANgemM6nWhRyfXZCKeG1AbXComHp/6oMJ/NUjNygd
nRJ8H9+BQdFy+WYNmCMrjmzQTrc0qqnRoRiuHhpsM1suux5uUpUK8CzTZq2dmK12W9RFRQ9ijq+Y
HNiFUxotN/RFcBzmZuePX6IKD/MA0cH82rsVsVzmGGuply5qw5Nc+OrVGkhkKMVnGuwNx04fh7Jb
Pw2khZ96KgZNv2HzTvDUlfiJGAbDYy87B89hkEbydn5JjTjHhBo+8NIKd4JzArmP2fF+3bNTqgm0
RLCNE+PW46kni2oYAPAAVcigJZ/IP08D792ZQ59shAHRWGvzqc/XrQFYu6bP0z6RlOqYwWpH0yhz
4NFScJE+1m29PZNIw3YIcmulN8QvgTOUFkUZSBurUVehytLDQTVrACe6P4CVRj49TU0bFRWLf4rh
0aQLOzDchgM1nNrEMaiw0PdyV+YU3Z+iBpmAQ2jDHabplMUj2SRygYrBBVyaEl5voSqVOJtPKxuY
poeEa6H6RcKj/j9ecEkKF2QMmI3oGRAN3jmX824hdyKBgwEt0EHVKrTFsik0PeuSY8RD7aQir1rV
JpoJkLoivp4mkA2udHtfjsc1QUoABj1/J+evsFaLufXUr+ZS/UCydC14zKM7KWphFlezlQeCGLkx
Bhw8mWIvh9ixXOYumkiesZNazy3hhn/JCxOBkxlnTqoYOm1StwRK2Y9BMWOUE/QTdRTs2p1Pw8zu
OYbPLFWfRZuwoXa9TBQRjKXU16Lw0craxPAveGxFknT8znbD9o/2uXBGYUe27x7XW9QatyAI3Lus
4rNxf1EUpxHEEASvXod3LpzfoeswG8SXwlWzCvQqOECDkqC8p/GyIGc3V/Pt8Tbpmm8VFylxtGOW
HOODG8ECXtxiHrNYR8qmUeizRW25ulY2PRoKwIM0VpcI4AqCOzVCljl5tWPavhZSsJknpDzGIXOR
CKLU103edqAKxgFzd+KWXDpw2vo9RRk+72JyPuSCAJL4Nrrb2lyIRjl2fMxc2ucp87MS79O/KkCJ
sy0YYn26L36BMqPYzlOJKYs8Ytt5h0Mq7JDB8skKQjUqD+AXQ3nrpFeI9VyKa1w9BiPgsc+CNh3G
Afud+qCcRihBCuUqEEe2Xig8S0+J5t6o14OMEHXUHALMyN/pjESWO6P78wPphlUYN7LDIMlhrluv
lStfHY4+Jyk8qirgi62CaVys3rMgommpqZRbfWfGKgbOVpO4k3iC1gjl/aWXNQE+emVFdX0aHRVq
KfrdbSas8AmLSyV2lQhbTCmPhrAfKJWFxchVx5g8qdID2YpRBYlO5VYTPJDrLYt1ufefRukXSzDF
ShUZHfFgww2jwtcWnfMKgbyXALxpBF+pmRx+GfMj8DfyeCmJiMehK0dn1YY1Aplk1nNnr0C0NnTH
ChSp1zU7LUm1mIQWoxt2+ycmUJXLM5HY2bB/JMQNu7hhPBpgl8Wc49KXH+RsrjJ5ZIpgdjKuri2Q
5Om7pJ2Q+4QA63QRZ8L2p6GCKAXlHcca4DnB4yPE8PJuC4L00a6YJNFqIL/+CViSZO7s89DT49BK
q6n9+0G4ictjLrfbc3GSxIz0ixQ8dGjh7HNLoJhim7ym+KE1qr3caiE3I/ndDCPSoScjl/gKHPjG
N5U+E526uWzWOpr1+itBLeAKLsvtvREZX0N1hHhZ/W92XmkHialxZHrfCAz7RPjiFIzniYzhBnpg
/gmp3Kv0fAAyGGQMdnmvFb7+DrxcBrxWZc7QI39Fb1MwVSuFdoJW5RomoEw1E4+lD3xvS6cu5LOH
lhC+xFbW6U8S6BD3YnBRlt6RVy9Bl2p/SFEAR7xaNiJoax5o6Gi/uhaxRN6cj5zbEHOurPXO2Ypq
AWZFb2ZXGlIBqUdCdckAYvADSfG7SSWg6XqIlEFRTtgs6llppb5qk3MxPKRHx7v8yaM+/GIlxA+4
oAEUV27PCBMcdXYV3KcpY9NlZWAZIDQ21qymCBYiim7NP7DLNeAs/imCYwNaGWb6ou69+/6SM5GL
MBET/IA/poiSg6qD0HXSxqH8hS6wBLhxuKeMrkiA3aJqJeawO+Id9VQpbABpGJ+RyjG9z2Ob6bkl
q6+U8cjIuotXwXY/JBpXVZXf+sEFUfEQ1Zazz1EgbSeXnwSEzpQY8DJzeNeCKLbvqyuqZZOEbtk9
LSv99f6Tdflj77D8LhgnWuYzBreZnDgK3B9zrL8qLzIvxU3+2Ppd31x4Som/rQ15lyhcrk5S4qHC
dnhfM8OZWu6K70INtuTMxyr75QIK/bSL7OUh8TQ4TFhYSjY1dLrhv+e/X8cdnc+iz59bLiLLHAs8
wX3I9M2b/iVH9ce+MpxMQYg2a/YTaZ/mVOfpsjWtJJhDRkQSQNOA5QKQXlNX2T+BZL6mDT1db7Jt
Cndwmi+QU2mqYlf0Vu+dMPE7yeCsFwXLBQz9XpGnd9hUP4prC3sfJsH29XoHs1N8VVyzn8G1KF+X
HklTw9mBdWBRgG8RTCB7CT6VE3AY1Y3AxWXsVsLjL/jmMp+L9jCiHGzw929sPKeWL9p90Un4gwjZ
k7nHZs6YZ1/dphdC9eDFawTGa2ue7MAuxtbf1DByepH8RssgmWdiah6OokMGq8Ud4sXu6lSlRozz
B8TILgdwXmCqnulvd9GXOq6yrcb8DhQ3rq4ZsDF64ToB+NYpnQDjHKkWXdnfGFk87yXYwrGk/7wX
rEmY3Lxhj/5n5IBeBb6/fEdMVoIEsNAaPppTLc6e3dD2MSG62lBVvpHnimE9kS+3BhtHRRCG5nAS
qzoz++jcNHKIpro2fT9OspNQXpj/kvEHjoVDmJ3pLerXYDdiAo/jXkIyhu2xMXgWsulHsigXAa6+
g9MqMHgfAzf59zkZ0NIeQ2dR2s2edoS2P+gbqbcbtHIGDfeVqYwTBpj+8BjrDXtz016z//BVTuD6
Fna1jPkWEOS/GbBuHQwYL+/CKH7cmh7tcTjeUuloXUerXzTxxA0wIY/3IENuoIHbOSDTGs9PgExp
ScDjSvXZDQ+2hQ9rGSk8LpxE83z5BjtHVGcMo8G39NwaLClNMp1BCMJnferv2y8FuNUCOgem8DHo
e4Seo8xeLT3lNyIYETjubqHz+Gutw4hHE+lKcD/yjxXLUYLyTxldZvOsjDbpu2mEMgrYDM55x7PR
pbmpMqljAhR0l+7Ck15qyaeqaFOJKnRW9MVZ+c4Vrc6MUS2IXRlDY9h1fZ/e8aGwzJoqmiBhCwbe
UpmuMtE4DbftZ5lTyK8l74rK8d+eHth1IEY/Bys/1LJMD/sq3UhFIlckg3zForJtdHZS5gFUiteX
qJmRImMPIXxH/TPTEtuboygucnKN1rN0+zkEDkeN0xEs7bsTZ3Yr8IYGntCG4QIS8SMLfHDBODgK
HQTTzMtcIKW+Di0jYz6HVB1eI5M1i7MrxSnhMhJvYeS+6PL+XCX5dMqpoVb9Zl5ESP4gcFCP1cej
3eiTFMGf1dJylW4pqQiL8ZgDE75QHTQt/nXw9tOJcVvphbzN2Lja3zdd6TMcJzPetbLM2z6H/XF9
97CWnPQY/GNhV8i/RQy93CBtFE8ZE44W71yQhIeRT3yAKEYB1Jzt6z6MtqVwZFWKGm4+7rZWI84C
bR/XNUDH+QAp1TKnpWm73ZOqklnlpZnES5zg4E3M8hEsOcwrNGQ/+qaSgSZjBwSJ16G/qi89Ac5f
jcCd0n7R6m5risTg4zFhKfyo8KeQD/62MIZCVh0Ea2yxpdMMwlLmRQcFgP/sabjjJAj2ohjOjjUb
Ylc9F7gkrEuI7WzvxfE9ekvUiHC5NWdhCqDxAS8GsejtxN/ZSC5sbfuZxsHuo31f7FBWQv4seAGQ
G6HE/us7pq0Z61ui2UbUL6icV5tBCHavp287GMpW/VzAlgh0QjBR0kVmCckel5f7NgUZOdFBtPLO
EPQS3B905JU+iA2xZRf00K9OE1Eaot/RQ6s2OXjQqCoRrIuG0Y97tcdvtFj9EqzazYvvZfqjSj/K
FJd5b0o2weaMflqncXCdOlnp5YFXZzhAL98ubhm0y9Mgfyicqdj5i9lgolDpRGZgC1Z69RrVacht
fS0d3lQTyqgJ2B+ecxw+Si3wkZxNAwkV9CsoBJEDP1DTnEPNF5ixRE2r3018YoRIlJqhPYmquwSV
Xz6CxoIEUuO7qp2BnejsVK00xpCrQInj8qqSHuPieutN3FYG6FuwlVtSaM8UMWi4t/ozpKjTR8g+
lz63ttuLRNgg0zG4UdUSGb4xYZmtI5IsVvtOtnE0GoEna7qT4LcEVtHbQMvJkBD0FEAQU2Sos/H9
m/V4b2aLd010lx9EevaOjW4JpB8/LMI9K1Y+9936dEFx9Mf0FZPKbqsbcyyG2aeMxVM0HqxUH6Yv
BuWe07akCXs5DJRXf6HnWfSE+qqlglmGz4YuphvGEroIDXeocXLumsUdSvedrRRBafsSh6I0ZGWs
9wvR7zN6hbRPTh1Y1hpK5uaFXt5W69aErTR5unw4wzHzt0Bm9exHj4gv13gTHPOk3S/uUaYgc/mH
3sbGgPfSX7jHAyFIKHVpVWKYuSEwzOMI21qDDUUOqDB2cC+o7AmxSDw0kc5Rp6P5FFhplLKp+VE2
Ggr3/QaoMBisjkK1CTZkDlNoRTzx/ioWpYqmUzuvFt+KBBxsxte3Jtv+gldQxOlTeoTkVXuAbejp
VxxDAIV2+roRt8CQEN/9xcIftXvOpc0SpNXnC2MAUs3mSIM4MP9/bQN05+18S23JwdOslIurjz2W
+/wVeDZ9qj9xqgHu5FkEvd7rZrIRPju/yyq8AsfpT1uw7V03qxiX19ZAbrNZXvWwGHglLkE++gg+
dBPgxBF/WLVI9/ehDErZyzmNkVl46gPDwOJYlsCpN6i45jzfDq+weN+0YExvfbm4rzU9asx/vl97
6JF7WpnvlbbZXBaih7NQik5GhqkExtGn0Pjj4S5GYxwq3402Ettfane0gLfunlXp/tbliGUwBXmi
iyHe4eHVmiaUGEU623SJ8F64uBVD+Zt9HTlg4Cl8xG34gY6YKUIGocuFsCoxXTpRdryr+ZM2XBb4
J1eRORBLh8jYx1XeVsXNXzz8OOv2ksDHyNWqIK7mTYBTsLOnJbNXzTm/AmgGmlW9MaZ3NPxf1kiI
L2yAffBrdMfcghuSOv798tGe87PSSHCJCaxaKmBaWUe2lzyNzKDGVfGAoj08u/HAg6HaLWFWCtLV
38Y+TpZag0a/RK7AT79WSDuXgsrWX2XISme+sB+OBkKoaYs3HtujzmZwtsEeVlkAbuiKNjCwaRIW
pM79CfVyldjmMMYT6radqXTrPgY/vZFebmbccM/SfRm/+MI2fHB65PHLJ2VvyV1qKEX0kY03Wu15
I9xu86uYp0KsE8XLjXKVg2t4Tg9SHAgBqYwA0es7P/KZJi92oPtyyB3D3+PxVzIvYvNv+lKsyUyM
vE4R2qHVUspwmCM5SUOEDIdK8Q93KlZtpKGpO57e97hSPDLRg47+kiqHvTkN0ZdgU7CJi8cRpyl/
CRDcv7OkWYSa3a4S1el3IQDE2ygGB4qvHxrs8gtnfHntFbc1qn+fPdT6wywZy8JK3vB4b6WoIXsm
CJRD5tHja3Bz5CU4n1V4PR2oBk8V/bQw3RIxYfYWXhcbAHIPAbs5m4jEzzIX/Wlc9NkeblHf6M2a
H2B1hOuAOrKE+Hr34KR1ivOmSAfzehhcPeScUmxIPeem8VKqJgO6sLHv6croDZm7nwAf89OQGEfE
yDgiyOXohnH+Kw4Qzs2oVssMpUG6EaGHyyT4k8TSgf9VBuaje7/MTO/eVz22a9FxZTuO7EZZzsQY
lxY5F971tFxYevkQKCZJTAms0qd0Gxe1q6DEnoVChiGMaHV0iJLD9VjVMJkCwB97mCVCOH1AMUgF
veHXCzwcLKkXptnfC5RfCfr7EyrcD0Pi9IccFcrRqcCmTbnVgMq+bF1YbS7GLa5gFdFnR0OZydP6
gu2vA8OwzUAtz2ZRh1fDMmYEUPQujceVHUxDxlQ8ywW/430lXvnUDNd3Yi9Yg0r8WV4/qHAyxJWF
ksoL+BTzjgUFCU6QIqZg3fndihQq1ZFG/cYNsKESpXh7rFULtYeOTq1AWgHErnl5tdL0SjLITMfE
Cc+BpL3a+TBqRFV/um1avZiwYa86nCat4WrdHIVBjy1pcskKZL9FK46GCpaEhuwp7yODCeXRVD/A
kkbMxAM/hdnYYO+Cb4Pzz4LiQA823Q2AojK3+yIv3DnAS5UI0iCHyYnnh8xXdZuSoMkd6rWnRwJ9
EOpV7u8pRILz3DJeryQyn67epfgskobf3IPGJoMPxy9wgV24QagPshNUqXYvuI+NNPJL8SZYlkgg
GVAEzflY9hkXeoMUvulAIBK1n3lLOC3nTrFLXNWmJP9cmeXa4hXB84YjZ9TXcEJ3gOhybRIYuKbd
KleGBL8WP8HHbqXbEeTfSk1o1UniaR5vJdTmgcGbAyn5u9JOIK9g39gGdB1465dQXQUvZKJ8stv6
kAjYZeuLqaom1xG0GWVKIiovzc8gCnqC4i44ONr7U9Dy0XQMedf2794Ha08083wMH21v/IpGEDnd
B0zE4RyxVMvoRss+uEm/WfWfJLQk7x3G+jAMgKvpP+BcEzdYtLM4+qO3AqWkChHkjGEnnQup9nX0
glzbS9I2eChtvxUYHEPpE3XAE9UAbfepZf7rbn1PKiy74z6g2QMDEWgKXwqR8yUk7SUYgAiZ4pMt
GiFu4oNEJqPpBXFpBDTjxGXDfkc20kFm4obJV7p9qqOUknEw2CK2piwfD7KxsFLKtZ355I0bp7em
BlhE3+qbDI0XbL2MfKQj3ix/7mrN7jk0msucvUdSTGFVWIIwxHUNXNHWhpzQUS8qA9New69sCSCN
FS508uOHzoLiNzUaKLOOesLYCfA17YMAUsIN3SSMirmPxNFWa6XFGlkUKVUsb06kQgH0NLTJkfov
9FvydmLQu/sBw/JD7InZmYimLMLAhXR/NGsfYVGCHiLv9WTzwGUqjCaLXBNnd0AxkkhN1nl0i/Ub
BxfDjQ6uuHBFUlts3wW/IFgOCBePIBmBsuItO//ITMKDmzv453KUFfyzC6eQTlibnOQjuLyp9fH/
Bq4d2vporljAjWdwqQSNCsd9kGJANypPrrR2P4B/aCBsEmhFHtC/5F9cjw7Pf+/cUIY399+el3MR
D6UYNFFJFCofnKMrK/ChF2AzY/+fDrPujKXDU0U2pKnbTJWDYwLaYh/Y5mupj+uhMNAOeD/D/mxg
fBZExGX7NCg2oxfelEmoy/pYHJgru0mQuQE/b4Ap0xkHBa5RGjYRSaPK6/ePpWXRbu6hx/iUtuXD
/LhgGrLcohSz/qGnwIVRytrZ9tcnRJK721pCv303ePnsNa4Z2i8qlertyZ/HPegzjoKhg6+VXlPz
Jjn6s9qZPw0tIrgd40ynfwkFMqDKXak3mC+IJySx91BF2Lk/2A73nT45Y7RW8EJxzAK6zC3pgpxh
q3KIMW3tyCRCg1fDcsTNm+Ng4f8kkZFk7/H5CDfpx5NvG99WvXW0XnwlPyyOBWleZk1oWLl9RYSx
a2HtwLIoUnqz/WXFuckCQRF89IsYGH9hgSOhD/DnO0OnVUzPwY5nONW9hnfhabOTj6+TjoRqA5/s
5ouHkQSHXssFH23Z/n6+o6w/Ct4HzXxS/n4JbAAUeWiyoIFm4WIGCNZwU4lWPkxLlaUevbsIZXny
bxt3aOODwPtc4eMKVUQ6ccd8KZGr+XUrAQ/ep1Q6TN7RNuohMeSCyfhYDkl4laeju2J/1EZu9vsJ
vGqAENLLySnnqwlsKbUXQI5j6q3REoa2xUNymSDcUlW6q0AWuknDH6gqCACdC/ockQ25xnlFEs4L
zHoBApB1xG9ZrtpFYdKFCQ5cz+sz+CCSIjlBTYCX5IHklqR2xQHPQtthGAV3AQ2a7YJXdKzNfoPo
Zq57ZoHZxhfiAT6KcDBPZSXjJd7Hvd0IxHtE+UurhHkQN9nQ6Rj0vP7XzNrGljkeMzfo+bSv8pYb
iiiUy8gIMZEANSlZLyjeRJRjGWSMvUPHn6tCBercER05l4/k0VM8mEwGdVukzrgD2f71aklhp/zX
ScMkNnEV84V2DkhMHwtrTX76cxYqMrfrhZqkYd4Q9GLSW1mMtG4IP5QGFwoaNiRaE8QdcwKCdWsr
mbRDSi09Bi19xbuf/J6xxzpQ+KSjHoEOZXb8gku5aHPyTzK85GTj6VDVk2LjpHZ1vQlIhfTjKijz
ktH8flrc7/AaRtMScb1E57/X2+G3BNGsFAc4BlBkKBY/yYoQkTzNt4rbXKkKlRd4Sag1FzT2bc1K
6i9r/Ud8BPDcg764vNZ0f3vjIFfNq4w4f9QGyV9Ffy/k/+kjpreJLvTQ/xolgIvre+avn/NchkEV
qZl5zKmxRe68hk3/4auewqg3WDcssnXZ592TPmt/FgoxuGYXOJHcF1UO4iWiVNlR7qLkBSrkl8mv
jPaAkXUO+JdlLIR+K0RITqpORKhZXZzMdMDNCMcBV0EsbSf5skhMOM/iwVLDRCkaLkISDtbKUBTe
XJklnSHWUFxMqewxEQOnENM3avZJEarjrCDGKpz6qSgtjLqWNliSt8+KtDXEE17ngCvPTl/8eOpd
J+xApAIdlSqmF+zxgT8NquJheJ/+k8ukgFkatPTuai0k+oP/qPdtS6Q1K9lMDpDX6Sdf0J5xa3RA
vj8fFoDxj8usr9afQk6mr2Ph4X3mDt1UzVeynWJwHL4YyUwnC4yUn7Rv7tFTGnwYn3s9R83Fflf9
8vgbBeKA5H28Yv9XgpdwHx1EUzKWNcSm76clU1hUvVaUUuX9g656jkXK37XRJ8HjmgdLYzsTRjM7
2cAyhUWjLngwUNI6TgC0DJi74b5DZRcqlILbsuGlfFkgY80Mfeeg4NxGzKRS94TZnPDxif90TS7w
c9+BO99XW2wwrYumrJhqa0vcVdmzWPzjY0u+byDSBu1MXDAMag8NVa0VMZm4Up5WVpYltHTMO+wS
bE/7Opb7sAMZK9V/ynTxq0biOEk55Tw4IWATzor+h2rfu9M3NWf7N8NHbmcTsXS4Z/m/d+2C0f80
oLjMj1dJ0v9ruOqIo+TMBj+E7AN4TFN8HQt0EtAlRKW1KIETkviDxjHrSooVXbspXCxkmfhrslIV
+2t5hZGHjCPw1CAeYRmMUXF8gQFd0r/II4OpNp3gpPJW/NmT0j8H3zoZMNsVpI/AM0gRcUYBwMBX
+Po4JMdqXnNTKaNb8lOYZlE2eFTRTKg0RCNmXUea60EbL4Y7AsSCJGRsg6U8NDv0z9TtHNS85plg
831gh8ReMEu4V3/wFVps00fLNGOfQbHqzEa7cm/kVRu3ZGCqHYhcGcfGML7DeErIzxlwLgps31Yp
M/DKFbbrETpwoLKVhIqJvfeWHMe+1h/VEI+Cu1Q3NNvh99lulKDmO3tWccQTZ0vQ90V0DHCRgcLy
67zutcwoETZiiu4tvFJuNFqCuZL68YqSq0+yCzeVoEcinPO+fDcwl+AVVaZ9TymGv2aA++aaad73
8o6CoWfMTHz5zQH13VcKAAzU+zy8vwXLkJ6yPUc06Ms6gbH22lmDPLgw9prCdOOC+GA+vzVkH572
W42QJhwrTkAYCwhk43frw5w0D5/7vn8X/eaTGmREDOv1aAFGqBoyeCKVD916g4At2GkdN8qyGHCx
S0s91y6FdbqeWoSzFW9APyH7n3/ASSAJng2fwOo6EeZ0JNGyLOr4tzUgMS5XDb9wfWqtvr8nkKWO
XcstXP//kbgWRNGNqeLRATLGJouIoxlSDqCvjEMWL4UwhfQZBBLPQ54yFLRkrzsbi3LGrLU+OMc0
CKQFdaXSv8tHj63fL8Foq10oS4F/Dikvh+h7Cihx0f+TRQTirRA3k2JpTbrm4PBgcittEXC0t/38
h62a47xwun3DqQU3eQXZGMk4dPlqFtpeiyEg/gINKxH3UVBYWMiUatfW6oMm5woXXEPUir/e9Gag
a8Oq2o9XI1lotJMGKN8OCH/B7jZ8PDYsZpXBGm1ZnLHLGXnrebO4aUO5cATJOuhWkVXcACjfn7zJ
KHoUhBPioxX54zMFphzOlKY5BaS/0lMmRaEmgSFpWwNAAWLaEfcEd175RbFTixCxKxscB/BeG5FN
S2n6ICqFHFnITSyZmXro9wGtHjfpqI4mSVRpDwbBcxWDsyB9kDRnnxRw18x7R8Q6v5FPKjSMFtb4
d5G7Uv6B7F+l2Xp3ClEpS7b3ygKx6wvG48/pJirmHsTEePX25PmZVwhj/lgvdeIRO9umlHwl+OpX
2ZLdXwOBlMhz+01unQJ/KikkcrbjkWoISdL64Xmv9YBsvnzQkSUKyyhUeI6jtFjbbrjOAqsli4NN
Fr5qn/lQAf8dlOJlhUNa+8F/KMWi2NymP4JjjzvfKL89nRdjWaPrLYS7EhG0H27OylUrYNwafqGg
MWpYM6eVIvEHL2IQzLN4p6SjrKxqaSjHZMXz2R2BZFKORueVeOOpzyrMIfsZltH2nRwfrOXZu/my
dE/J2fwZ4EGYE0uqvmqhRWHFtW+55/GWeRtITzPYiSisQoQC0IyYeld5dQOJhWv8Yt/kTPBvkF36
bD84QIOHQE9AZfY5YW/m0CFc0BdLx7iRbQBLrTXfs0jI+qAOU/Juk74equnJFsvpuL5MvK2UHjdz
XX4ytYiRecJ0YczziT68nSoKPjbI/5IDOgb2DiAZVkowoP14V2W4dtFABQ1+AYyo3CcLp0+7qj7D
9XbqLrQL8jss5IIuwgxBaGgWL/oFHqnbYtj4VbzoUePYAE/pGBzIr44eHtLw/qP8f0x+zJXerFkW
dSz6wryo2c6c/SxH6zGZGQ4AepuOcR7mxa8X4btmzTJgLvWkPeA0J1BuhJjj6EJS4D+YUgo8APlD
AxfBOIhbvFKtOQPGoXBndccYD4ioy4hdCmcsIvvPdWHiFrxFA09SlmkW4LEj6yrHyVnpCXTcYYsG
kwNZfjJXZeAKIpmlc5knTHMznfhB4noQ5Is1Aow6PPqeolZeTXLhriV4uXMPfROG33RCKKz9IKJY
PjWxJZxOTGJa5Sf+ApG77lWigHmRE1P0FWJsRfT2At/h6XdUhg8m5JcxIt9Ou4qI2UCw2R5C87l3
FyDy+eaLxAgXuH/2ncEPqikhtHFgDfwolsFONwUunVIEazyXPdrNHNy1xRcynq1RaQ0rFiLCj6H5
wkcWK5ipL9paUhiG5k7foMmC3tm7NslbJeXfntD6IdEDIPiJI5k7b+1nd5JHYQfjIWySFfLOOO4T
TsToUbLDGGlS1wlSDq2KT9vTA9us0oXVw8CpDHZLynV4Gbvn5wKemkcolVn2JI3X0mf3o0Y3eCmu
bMHrq3YbJN659vrgHT3xHS2mhVovSifEQ6/jR833a28uCfMAGbgoHPe05lvNCNk2pdjJS4cV7JWr
C3434DiuhjfPf2uuopKoT0t82F7nb1e36+CQdOnhGk+aeOXmcI11ScfGSLslPlRAXliaEmRqsxVB
gWd7s6/OD7l6+kZxodfSrT1K/UEGrrygYNADgjufnjPe6i35cKJubcYcHcwMO4LC4y5P56DvfZvR
ILvSPrVNobq2NxN1Usd4C/qnTKUjctVc10/hQTg7kvsDr40XGRsaaRh07HT5ydGfBIhSJDNtVY4y
VZkPJtwLjsKNVfVWDu5A2VYqv1x+Uw6mWWyXu9UGaEwIEP0UamSZid1EHGl5L0mGfU4ELzXvI7sq
rki39l2pkQ+wxNBlrhA1tmxQI+0aE3Dfga4Mpry6xGYO3rUnn0bZWxfpL8mZXZBj0aEAY8T4Fode
Mr/+TqGhJHBc+yCpCRt5/0BP/9nAXud/E72yHsvBr3i8sVzOhtEAP46NfQ9vjL8OCYKjEFR5WJSF
X9gAJO8VAZ/XjVp2pTx4GmIJ+6pZdblR5xicd/WC1Wg6lLGw4LCBdFWyAlPezOGx78GFnFrCPU6a
QUyNKj/X8LgCR2zd4A8uH2OnOQl1K+jLG31jpmk7nGePTC9WRvmIwsdYX1rJszVEeFsCKUqhuCPV
6KGnzbwy3IXfvHHYpsg8bMBaQCh5LuVoCC44KZsdBxCTu/l7tBqNaLBw59GtXg4C/f7KQTtMoMFo
ZrwjGZiksVDAucXTVSs7IRUabgyGXkdNcrXmXdTwGlco4nYNPA4jr4uWV2CFJEI+1xRWZzrr/YEH
3qxfDPo0FgyEcVyKZOwujt/Xh8LmQ8nvLlRyXxFHyWB5QnJuv9LuAHJeRBpeJGzZCYd80HItriN2
QOF4QvvNnjHJ6eKG+RCy9a0KwkYPbJlfsIziuRUKWW2uHi0th39WdLTvCjEnm0FyllT/gAN96lwR
lJRD4Wkmvhce+HOhJoqKCp+55ZFhwCMgeOUE/QvnU+hVywCYrEBOftHUahwl8RMcusnvOV1v8bJv
pDr9lj5/Eff7cyWB4dsc5q3zAa+f1R5smm9giGilnnIPKBM3WGAqR/PJDUrsaHd3XlgtBiu3hGyb
UWKPrxEZPKNb3V8UU9wNCOBODKdoifQBaES7R2FZuLy+xlbJUO0QzzJK3MXxgODU0MaiaP5qqwuQ
f9uchBQIfAWilFFg/5aK7ruUIcCmmhQlpMipZDMeBgoNymv7A/+ZJy0uLSTpJADQMy94JHIfDyZx
RsM3takSE8i8pizUlMGyFw6mslAWGrex3k3f2Vv7IJxsln8F2Z81ktoUwna6O4D5leD0Lagv+M9/
ep4dOHApSGXWN4iFtDlv165nbxoVeMiigVmEpWhjRvtG/0wuE7yyks6dUqJFjZmfXIgvbGc0VoX5
8c840udHgd7XHoPuwsxeUcjbJCFhBthmxuzWyLBZ3yDxVlzai8GsXbGyAe3LTCDt2CyHtxbQ1DeJ
5c5wjDA6NxUHK/5NQBCPfG+/mTRhktSbx38wv9MP2ixvJX98GCrWC4cj/eVoleK+GfY4nWhcKhec
7d3K9WdXsNHXtdJE8kJYzrLSpzIR7cYIGhnNvomjkYpywKruKb3l+qzNMEg24BFnKTygsgTz/lpD
Bm23v/VRDSusn1SGGLsaluL0EvzuCk8mJsJ82Fj4wX2OBAFX0DdNexcKrIVYk7Jl9qZRcVxN02sE
2MVSVAiG4WHQIDy5nHYrlXUbJ5yoVEoVDIxwYOo5BymTTM7WutnA9hU62XL+uiHXi0S6FErLFsL8
7E7TaKWg3dmLnICm2DJ0RhyHTcDBk1Hif7eEIbIZG8gtIACqLyNZ13n3N6x5zySiDbfY/GEqIBdw
SFwmPpXpx8hSGRBnjogFm6ZJkKTgRMynOxxpJ4nAtKHQuCJIDy+u7E1vLBOKI9aMMhKIG1TXnDTj
m+ro93wnTtveE4AuX3JbgtXzCV5AMT4fSaQBQKWSPNo7XfpqX30EVAhL0YVJqT/mm5foKm9j6HEh
GN2Dc/J8Ngl60SRYOH/udh3Db1yRLeYnjO85HUhbhVruMYtKP1d1DD2SmX8/hF3IQKDFgiUjzebm
yY1gu++uhnMmy4wDttaRG2dWfV7stywj8G/o3jZowHFT0uMfcinn44+vLLwSXw7Oqc8xLlPdKSpJ
58dOEeJhz3cDUZICCkGIKeqXdJBRrJ0gQmjTu5Aiy9UnUqCImTiafNEyn27F+d5T3Z/p9gUerZpM
2zfT/Gq5HehSqOytSGaUSl96CQSrCd+fFKNutBQjYNS77szPsRmgblgKljdgUwXbogYvb1bsrpoA
hznrf0zz7ejcHaYId1Bm7bdb4owoCtgttd54+EOUzDWHhzvAzgNB9Sep6LUGgfVQcslvyizZ9GRL
ENSgPXiFgwAhPwXElzPVrwHDKRhMorCq1J3ckF+zL4oHmqvrRE6nymaxLye4ZKibJ6cORQP1vUY/
tT92+AkIL76FSipbGTvCof7p3lzzr+S+ndL0JhKwPcjUFivyLwG4joM8FKVT/4uYibbDvmhiegvr
2Y3YaOEUmZSR6Ue0/94rCLeXV4IuQxaoMlpENW6zo+Wk/YGHYN/nG422BMoVuaodBGgRs4hrXEy+
DdoGblLn2o4YJcai3ufSwEiR5+tn0w6N9A9D3tULIZtfsYcLxcyPxBrZrI5Et/TZ1puYEsFAyVby
NvILmpG1YT9QRTIyVt7wb0GKxVWwbGFLWarOBxl7QodaWad4W4PRwNpDqqi7s8VvHGa1K5EJgwTA
/gmRpMGgoddjFE6IRr8OnLSrcN30HLvGN7I96WXX7xbU3pF1SlqrdgKUV8D3zD9DGVLwmNYCh0Bj
ydYGvHvNc9hMHFxapxQzXran8OMuvd4sZk8P/a1g+/ZONW2jMm2dvRB4clirUssQvsfTRPmIYn72
Kl9v6q8Zbzgfff+J9/bnTDEYkcnnGI0ukRATiqPges9WLTBeTbHbsFBhoZOsSM1e5+Shr6g5Rr2C
nn8PHftPCLEsc3braTF6vYbkBxaEESJszF8HTV57duH3suJWb7qv+tC7xddJ49sKxVlRZrURbVmD
+NfOiN0oBpwl+VtNgu4XIBVoRsqD9R1XX5KrjHkup04Akf5fCulxAKiovl5bOe58n93bYhYlhZ7B
i8c2XctCZMMuOCOyl0mrvog/pESTo1vjtgCVaL6dm+Vvghc27DDZJpsQHUwJneUXFRSKAb3H3i+0
65nz0hc/AHOS6A3gn5IHCKVZR1V15Vist2Z5eOljNjRDc64dQLbTZU1Geti1g7XvskHo7+hOTSwY
/s56uUU0FXy6ARC9AIHldd7AUUjBfTy2nDm/q2kC/rj/BDZGicQlu0hJLZJGHNrUvQK1cJwwuVYb
nuKaw3x7aw9fbojWPEFh9lGBYG2TXMNm0+Ag67IbqSn5Gy8JtVikf1NSEx1Z93U6uewr932+H/1l
yHDVRbGxCUWZhYLU/QFS7l0HQl0YlZ/qe2U8is3L5pftaGVe4U/5oD7BwYP0aR3GpZDSOOYi0Hrk
cvZMHbJ7Oi88cf9Fh3DCRJgarb/hR9vb3d+2+Tbmv3V1ui0wqr/yUYWf0GNJ8krJwdhx+Im1oVKa
ICsqo7gHQ99N9wJqPX2z8+u9L2QO521msNFeg8MysZ+ZSWeMylSekF3uM8+19/XxTye2GOEalE1a
gdgeg6Pw0yGtQTWE+wK3uAIkrMnqCWzrwmvDbYM4SNcPTl7Lqfr3sWdkoqUrWlT8T4uYxT+pq9gV
aDdqcpG2JKivnNUVGHvO2im95eucbiX8DjAHc+2VDCwo30Fdo8FTxEmol/jKfElVq8sdjvtgd2tX
kmK/rEFjTRJN3ftj1nXB0XEheDczqNkhIW6xtKU4spp5qSmzeQuaj/jW+UHzJeNLaUGxC4mBZVyd
jZRxVvM8DYqp/3RVXB15KBXVRp+R92x0O3pc3JtQEyFq7rw5QlMT+Poxnva5g8WNG1AQ6wIqlBNf
9SZplDCJY09fkug6vgXxdUIRK6zFg/2raHWI6d1mm6ysv+dtWDVr+WqrnsFkIsi81e/zAcY0JntB
WP10AZi8Pe4lH8zx55vA9YC6Ky67oWX4JaHDIBSspTAODgACIEiYIC5685JdgO2YEVpnfC6xNimU
SCXfmcnZFzrn1OmugUdUDsxWJFOdxbnd5W2qUkS8435rMfkp/NnLQeTZTygHx+/bahqpUS13iKDI
A1TaLOkJy2tZOBGu8/CFRlCF0uHHYwwBQcdci/f7/XVKm6NhnDqjXI02frnKCAjTfc4MeHUxVO6D
N/rXumU5PXqtb1RvAswr8DdnSR2rxy/jBKyUMJHTHVtHQ6Hc9lhAMIUNT0SSlwg1BRQ65UAkcvT1
4FJvFEZ0JE0Htm8c+m2qRk8EPAa/E6XUeNdvjI9YdMp1DAbHbo1BvGP5++G9Q22Sc8YrdjvpXAdc
a10F4fm0DUSMNssplqbV5jd/Q/4ShN6x4UfmVYQGAT5bcDked8mqFnCUtJ2oZZ7W+Awq/8VVQVew
ch6pn+EYmovLzdkytZ17+n1ej7XMTLLLS+jvyFFazLhp6fs4FCclNPqvG+vQv+MGFtqgiRhpcCfF
kNE9FzDZSoF1Ba0OImsNtGbHcfiFg+XnZ2e+3hehZ51MdfTrzP/Fvcpj7nPC0KKrvcE4sFvkaiDk
iuWJe9UdrlQsK+VZrQLW/smrZWYWB5+cU3yITBywDZoDzjjUdfHMFJbQU30+1R48ooOsXXemuCGk
tPL1bCHzuFX3penQdcNuUONE2l3PSQD3d450egxCySDxKu5+4fMfrwwSkolqVh78GV7uag3Wpc6/
MGzZo0JMJcS37a6wRblYhKcaydrrlzlrFb/DQKOsFgey6yyivksl0ur48735PsAWMzqkpKFwbn9B
5d6CzVBNpgXfnaO0Tv2L2h+DWQtNdH4q7QN27dWZNHC20t1QO1zHyyPwxm/ZCYI9AVCSjd+rh3r6
xfNszworJYhq6QQHXo2gavqUnNjMKe7jJcFZ0DGi5ddvG9dhs8UWNgmHUTTFWCYAsNH8DCeL1BhV
/H7sBFQOEVjMYSnO0T2rCRypA3V/EaDvDdQSxUxQgxiNgk/ToVlXrlbRGZIzSqdc1Xf4SKboKXXc
GXLk/moxAoJ48C0O+ffg7SE6mDypn3g3gHE3D1zYp7n6si9i8mb1vkKKiicY1NDEflGt4pl/DmiN
cMfguPuCo9Ar3uBHmu2kX/DtoYSJXQQlRwHpKbuSwOwXOb9mNeBywyUsyEtcjp2VdYQ3vs/sT5AG
V+H65pdAHBmQTNpQphmtkK14/3zhAN2e6ZgKCRPHUtuCYpgxOvnK7WuAM43aE+zilM5C/pjRalOf
+qzEhvAAQuQAsXEtxq61Gjt6wmwL77T3qhwLqv5aOkO0A2YvxSD3WPmoQawNgFQ6hQBjgTFK5c1J
O89qqaSPueouuhyDYwRRGpLLjJEV6Y1/ltkuxtbtksODaWFxNQGK22Jg3iz+vORbJTTTRp07uTEB
d0EtqvuGBG8U7FBawMBU6EN6Da/xSzrccHbW0/7wKdJxn3VC/55ibaH7Y9v5aH3uVbwLlG2r+6Rt
Mprk2j03Yd2Ux19kw60aGWGT72THJGosvs9BDjcH6g3HPmdpu4ZAhrZq+iSGfbc/kEhrRWZ6pBVj
kK/UHxUeBwrI3AuLsxCoK4uBBLpEP3aOvU2DV7VgqUvPjkybRsJ+ofPNB/QBfiIYagPIuoIBmigr
K04i7ka8DsKeUzd+881EQixtrZ9J49/vzqTXYQYKOgaM2e+3M4SHdOTHGnKJ0tUPYXdHKAvu1i7O
q9elyy93nzZqdXG3gbbzGinoMPtE9RYR7oK1+YiTcYI5fcF8s4WfxKGNIyNxR5Z0DzeNypfYhQ6/
uJRb31o0X3moLdsF/sQTZHW1x7RAKeLk+C59bGpQ5NYPioWwKrMDzWvMazhMZRAq3CqrtDeBG9bs
hmxthb8fezt4/semOowZIoYJ52/vF06ephn359tQo3fE5P2aAJV4GtRhs4tB93vLsfMQ3w90kWma
VelU5wT03sEKn/EKq7M8PX2g7UJOUfcGeWzXRiUuo+xc5bjKMtYTiNMWN8CYt24QNN7w5z5oZcXI
hSN4LUAgGHIvPOkidY9KqpvqVFu7PHR9ZM0ZIOCGeU4ZFmirAqrVxxGJtr3Q/0Fki0gZz1i4rZkk
bRlbSS477IAfFJdu9UUtodgQq+jhTvHTdJqBlHgWSlquWvsBoe8tRNs7gsl0a5pco3gFh8S/y30e
8+5GvUwRLoRhVpb+/4SqWHRu3pV/XKbMuA9KNQ8qG18VNt0udFmn/UNKXqrgSnif4esg80hFiNvr
X4fbVl4GZObGJxRnX6REs52pl5D3/EHq4j6wQWppOrmC1HTej+FidrXiUnWrtQ9LZkv39vqbR4rw
dMo18F6vdbAzeIuKOtyRLzlviJL6+Bu/hQBRSwXPIJXe6s/bk7Vk0Wwofb5UKUJJrKz3WhAX6Cxd
Qro1ZvR2UYAvHoLPbS367BpddjS+uk8AMc2MPc3hBOzVfB6qhd+7zd6EwvlQFs3xanDuh9ZbvMTa
lMQh5Fxy53huRelDoE/WJIYq2MWtGr7M2p1D1Ay/lIJDtss10Y4rqgj33OPPyMz439BSXqQWxe7d
TSQD/STJg90gZ35KE+opvt3fPlBpZSwLKcIlqztkVm7JExWcJ6NED69SBZRgAlS7Ia5lcQizGAU6
o6zgS6Zv+EW5kujVIpF5yKBnDLrnORUACkmso1vtO4XHCbGPnyUavhlCzSg/nX8b0dGXGizMdJtk
4IghEp75RmFodcEwBXJKF9hshkB7L4VCx85WUM0SRyUBX0CWPSZLtaeRo4DeBjTeLTsNUBITcGne
38baR0ojVyD89snIUGNQJwKhuzRuK3Aj5Rh970bK7oQ4huGsiRyxyQvAeqYybzxJqfanRa/k4oS2
C39BRUZJu+SsbrkXv9dKRgOAcxyuOEo5tD6So84fpuLIOOl3qkJApwXtOVRoUPIitvY6tc4mvmZs
a0LeJTpui1MHFBgcqAeLdovnxb0fRBRNLa2P2lb36pt+51BXjIK0IQ1P5h3p9sCMVd8tlU4eyaP/
dxZ8gDwhQpSyudBXS4bt6ovshfeDv37BTLSkMHUHztVn6P+/jvGgJP2+tM5V9X6jj0gfbfUSOWx6
3DXvRkOfpjyC+tr0HE2+tE+NbhO3AMPb7YYHwV3N3OaTXjESFq9ssgfy58YINHXQJQOr78wrXINv
pnOGbCMhpQuo4S8tugLMbBMhfptlRpYdXkpB1gALCSLQUF+HZ+tgjCUYWvSiwXBoFv2GGFk83Xt9
s9EVnjj5o0AuocWZJu2tZbB/QDfBMYKbNpfdMkm8up19CAKGrHhY/0hjLoUOMgcCnBZ8FOxoAmWO
ZRazDTbiXl3T1xYGqOSWnxcsrUkZi2ZzsWTm22ZDWx717nz5lp6o18A0bBM0OCNSqoFom5OY5Oop
TdULHd2r4u3ojemEJpmxH9aw48ecCVn763lxnE9Zy86nGdpj+uj2wixyO3JGqNxI7ECNNYCpYKST
yusBpQkOSDfbWHxlCEAVlTnEuI5DSuUyuq3UPpEfVmHS6ccar+3omaqiGbdxyG9q74jsX7bve9vb
vwINbajsW6zWJIODWtpjuGiUCGlfIIIfQu8rI4UUpK/3lqbKT1Oh4VPtkLi9KamzxdhL2V79/mAs
uCz/c0m1ZckzcopBDRKmy5lzZ2N37BObgAjQIDRT2Lm6co08Ev4VSmV+CsrX8bKMIH/mNUYLPVs2
CZ2/u43Mnbz+Q2BEcxUizieYDbw1CFjXsSCYEoq8rm4zp5QnqX4h6x96oDcrhMH1P4D6+ibxoNMS
bViPK5NZPO936fP9KJP4tJnkzZ3NRafFdVFVRGuUDEgUpUMer+u/3ksr9ThhDpm+r3874Nm6Iah7
Q84HNvhqsZaOrqplmaGXENcd43DkuBfbuagQs8w8RrsUS0reyPmrj6ck7mXfwT6pQZjJQ6LQlxXg
mI2QNdutzUMGYMokrtN9cO1tKN2hHDJ2v7YLe6zk2mo7cczrVmfNHiY/7lG2XMOItcHFRkzTEIuC
FiOzCwNI//mHHHA/1N8YpkjvFzPvpWPfogmCPtgpkjk8aE9sK4ttua23997HwY+A4PygM542TK/G
PqzN49rkLrqUsRQ/U08fedsup/xfd80vX41deEMrIielFCD+KWXF/yBFhC6JDrZDl+L4c/2P8wD/
ATPC6qWu9prJsMkZ9uR7+S8iWgGbtp9rtff/ltkVFKB/DwipJ3DhDnzlo1wNZuaT2JA/SCGHubFl
V/B6aFghehti8b6pD12mI6YRBaEW3bXXq1mPCOsP4UpjjNSOSBiKk6Rj8m05/FG0sS1Z5kY5h32Z
lwNSrhtbPS8r2cSUt1d2Y23tCeSodJ1JhESdskei+afjQbK6TGu1ZDP7VSo+AwobrgLqb0B3bvxg
a+s4VEKsINHXSPGhoBo8JToqihnMW47UeoPtRf7NTf5EJi7tU+Dkbp/eJcGfurVp5tXJzdRh14Xp
VjIDt7oQToE+mNyLqnsL+WMUDX71PRon7w0BUjgo/DsIR4BWURVQ493+HZB6eejlCzL7HseIHQDK
Y9M8yQwrJFkny+qG6PEMktkahLc8cXG4Qcs7atqADxEaB21kR8qFE5k6F0ZQniIFXTi+BH06liFv
VAV6gOVjN/6hdEFe4R8FsiZf/arPyPU5TYNODYy5942N/cz34r2sQ4M/8iqxg1Zmu8CFpz5BDkHn
DMkI/jGaeya01U/iMoNH2IHbQFe8uZyI4Rc/wPsWE9gi4xkwjahMBya0+6Aj+9gYNkoXEUnNG9f3
62WFmWwsbmnfScNDyucD4/9HGTI0TWFJg62VaZuY2T2MmI8DzP5YvNXYB0mJd911QjrgPg+dz0mm
+Km0JD2AVqMDfL97iG/zf87N8Phyt9C9ohEfhFHGStocmf5e/JRWgZpziA/QKvDj0vI8yUjQ7Um5
ly9GlS8pH6aLfherGw5lUiAumTRy4jJFPNuTpGQKXdFl1Fno28eqo0HSSHhKtL2Sqd/xpjp8xZNm
Q7MqvRitmMHLc66rRkq5gTqw8kxKSInxPGY32SKy2VRmxOgK+ha8H04Nm3JhLOM08gA/VDtmgqEf
BroCEMSDDr2Ee1+ChimKPM71fLePHeON5ileHdtcQ5Mmje4ECHte2gdG7Cs61YtM/T5ojJ3q2wsp
i7Wzvq5lHk2idF6h1iFQ4kNoerKhAsY5Blq2WIl4MYmo7aIiA7n0lvLjF5dgA/AUFyJ2mzeiKwUA
iCjP/8IAoesowZiApZOMSErkww3ggo+dkaw1oUiOM1zVKa+jJj5aqr2Om/F/eJ1zgHD9itn3y89W
jnmxj1hrA3cStJz1e9YqJaqurvMhU7UmYGj53LxZKUn6JvcQC59BA+E0RDus/4s98Mffimfatnm1
QQoWu1yEQ53vSe91Ule0LxKRWfzjvXCx8gB2qB3UKHhEFpt1em48qqyO8Io6W3VLaVhqfUyPpR71
/abeUyDzjCJo6plc515CO9xO3pEpV5JZ1SXkJVIgAI/Kub/m1XCs7SyouUU1EWdi1SjgRtt+H8Te
sxWsPeOiPAf9pyTUHs4/E06PvLoU3hmwfLTQhDbRTMuAKDw3MHy0Z+HKdtTiPZceEA6Nu2KvNFL/
wdHGFbR7qB1KKPA0mcIXn79blzZh3OQjhcvx+gxkx2FzVhzqasR76+r8bpUIdSMblp/fEMfHpnzW
wHDjEvmHvoNIVniKVSdnql7uk6V0gWksBp6UPgkQoNcecAh84ZfMlewiwVeZLjDTTdE0roVFZm11
63upE5rFHSHDg//eNcwpJxUxZhFNlg8IhXxPJN3yqxT1IRwkFbLj3aDGbVyPkzJaRrLyhLzezXNK
oIbluuN7PnXsLZNwv+PL7LFDD5jyW1b0QRnntyBHjRwiFBlfcv0Mrw8liRzpxp7uHl5axixcnrhA
g0AVwlmUILEi8FWvQHmA5DYMBz4A3BMCTettluqpRXYbhrrCV85KJShyxuExThPNA/8TGEEcMLNA
3pRcGmmo5WncxWllLM6h9ttKvKiYX3kCvvL9BDDOdzpz/FXCwg5RntHPlHtsWrrheUL7oKAD7j3U
MPmuNTkYLyPFiLt/nMZgmp66PZWQtONIW9QxlHVq0ilydw4GBkoFFCP/UYP7+gCwxwE+hpaYCRnF
TbO8uDEQMgUlicVhaw9PZfmDExkk+PqobRsj4sQUkqFKZxLoSm1F7sf3EJtxSdTqi88uCP5nFqac
76UT/bOsr+jFBsBxovXKQdtqBpHV7EDDumXcoHdGvCZljy7BSVNh7DyyEspotfOtpVUeGteDDPO0
2HEY96jc5JBBlEogXASxMVkLz2b3H9AyLRanUjNG3Jor4kEKr0ExUnZUUMdx2ootNNNW/MxAk4IL
i235RZD7fNF3KZyMtaxyAjecnx2WLZdN2h6qBzqUVNoDPFYMS1ZogInR1sivq6uBO/L6J57PeAMG
SzBqWmmiYQz98m5+Nc2WcFY6C8CWNvcDh2k83wCo9XAXkr4XMTvLCDrJd8cah5Qny/yUPn0KAKer
JRPVW4GI6wO+QbxLt5Lkv8YAj1l5W2eJsLu4iSuLkdm99kisfsjAWNJWcQv7BqTSFlDCO4xlUVIv
spIIoKVOebE3F4nzL0yROZvvXUrrwy/292nj7jqdRyRRJ06e8FWjv9NfPxmOvwrQC5DXK2MKG3kp
FyHo3asfHd3zf0x+dforexT0758Q8sqcYOsDZP2BORuwrc6xpi4Nn9WJ9ICWjbQKVkcY0ecJBMVX
2Kj4q62sLsNRX+mdZj7xz73Q2fytcn1MXXFg6dFMOqWh/B9Lw39SPXuaRkrI00YYbmGKxkt9bzCE
J24ybwMkcMP4KscUzBP1jST5JICznzCDDIhZ/jQ0OncqLA07sdBgI2o5wy3grHwJmzE3CIjuGuL9
S3vFQkl8NgE+lWwQoCGmWsnbBq0gXeVfOqRLJbhhJmeLNtxDOtu32FDxDDpZ7Y1RdQ1Wwa8bKDV1
Ukv6f0xI47d1t2ouf5ekGKGPm9dOT/P6CvNgVol6YZOeWxDKrgQF6Rwk9YAJfSMcQWs+al+PKlrR
/ala3iA6HuXajP6GSw0NIEfwfs1CRR1E2HmSP2lJ68zNyK1tGm6W50d4EAj+A396pJso5BXuvx5k
gdkaf+Oa2VlZTG9dJDtzRenq0ckqIx1lCWZu5S349c6KLBbm7QlmfJGj2zQMlLsH+su0NFVDD5Nu
G3xXCxQFft0/BrUbH8uwrDeiHG5glA62dH1GVbE1C1uUkqm/i2sX1pp8ocDNQL/4r2LqyFqElYUK
EAFobzG72N/rHhqcw4nO3j/abOkFNdH7Mcfmylat8gOi0ZEBCU4r/TzDQ2r0f2DFnSU2+2+X//Xv
n5J24tBCplw79VgRLafsp6anwcVtOc9TznGPvGYUcDdD0dxuWF/jkid0/wiF1Ypc97wPb+8hsM4y
KGrYrR/y7S1A9S6kELYc9bFGLnT7T2xzKO1739oULGbwraJPuIQ0zQSeqvY+Qv15jrx6L8E74xHv
PPcLj4ubkftjkIawNK03KsllCRa5fVNxKu1zgHJSMNkxWdubslAbGSlvYKoHFZ8wR54ufp9rOA5m
/aNTfWoFBAAxF5HVVWjY50VS6zncBWAs4IrG5cCkj7ydP5uj8jEYsPIgWEsgZ5AexD4k0S4AbK/P
QtVoWncygLPYuAMebEcbAxUM7wVuWWqG9EP8LSv7n4tTHbxB3pZ2V2DHo7W56osD4SdwLV0P2EhD
TEECRjiYBPMcS7A8ayMu03m1eqBUL5D8QcE+xiGtpXC6DS8Uu/Zb/IRg0mLEFlmjy3MLhEDxoX3l
/DOi47Miz7GgTPY2FXjcsrYvBvnyh40U8HLrFInQ/PT0T6bgclbrvb5Yi1FR7D2cCm5Mup19TAhh
+LW3a1ZsEzf61gpJr7yOGbQQx+Lm2m3VKMshI+BXi4GzXL+B/VituSfBIhLKmPUmYuVgrEPuCWMY
3K0Hi99qr9TQiURQBYC6rzWcKYtBc6sgKC42tQ/ndE2DUTUGJRBmpVxYoqSf2MeWN0HeU6NkkZhq
Ggx6A9hzfuQkwl0ZF1BLUE5XnzeN5TkH7u/hfxGP/fnFKWfTfvyG6OZKOEM5RFDSYgtH+Y1M4pnT
2d/fj5HixNMr9UW8JwKO+Do31cnOwXx8+zWaGdv2fmyB09nhKuvKA6Itdr5/6XERKRXF4PvDGaqe
vROCPAYFMPHO6QlPae9inPU3RuSEDTfFDbAmEE2M3RAiphQgkxJ5OuocGnNoth8WYnW3ZcS7Y+P+
KRowFiQSw+wS/W4JoiW0AtAG1u63jTGrYNVUuPuUfxklyAlMr0z5rDDPpXNyEdSsG8laZH6lDrvq
AVQMJLU2yX2lbG4nTUtn7jjsBcVknc3aSUcJhrIdcur+Zk9HJIgblDyJO8fpdjotll3ZXstIS6/2
3KUWoLQMjbHG/kwr6ETaJRlyUCydKk2IqisK/+CISulOl7PsJPiAzHMYUgsR9APhXGRNuJKRxtKV
IB621NC3WqjsBkgqWDSY2vehxkkE89bLuGMwgbLo2UmMFBGuEYm3HFCkQx58iYZJPp2KfQ7AXpcz
H7++2Tsuo6B7MK4+LaPtERnWqo1FRLytBoQUG7FVTubuhJzf06h8XxnMpwIV91ap/1dZzCKGqraP
PAoW2ZAaYCqkE3XooBFLxYnD5uv5txCexwf6QJo/UziRtHKaPj4uU3Q1/C8a3715BGSUZBg3rSyT
av/tS+/t4UIAzX5srxIPMbo8VZrYi4yhtF0S8jKPk1ZYFjkJpbg3GS/FxImIuLibWxI+v8PPrgVP
YVaWe1p3O1cj3zn2uL4D6+lXEzfmzlMNLJtWEGSe+o/RHzOt0PzKWQHtjChsqeuzBaOrsXnM+oeP
xnWoV91SUPqqoYB2ERMgov/ArgwjCScKdVpFdxlP3vK/afiKjt6NZHBfyQiuPUz5wBiIlNmmWaRb
3tlY9dA3IAtwJJIy1NIV8urIvygdLtwaS/s/rp+LgRdw0/0Ae+VIX9+Qwd8sR8nQgUX2dTpsLh05
aU9uzCsMqAXG8+n9QyfO5+1Frbn4GEUuEFDa64SgEFTee/DS7EDsHLl0eG/0QaizMAdc1+91T7Xg
/n9D8zTcL7IlWZ706x7KjYl0etZeRQoEgUsU8zh6XM5qpa/Y9GP5EVnxJvWv2v/DlLJ3/rFDoZlv
lDtzODKZuQ6go6cJD/C/GDEEXPXQ+bYjYLSQoXCffNRF6/RGbT4wOEgBKMQc11hlHsZe7ypQlhwn
oPcCkfsG9T7jFCuHCO46pFOPKgJFayWaGW1+J5obmvEUtVgJzm1Q/cz1MWXuTJnLVeoI6CsLbIVB
zNOGMJ3WnjQaPS8UQeWIJxzMD3otoeGNZEcCLGn7M68/DxH/QcXnHXbo6AdLQ572a6+cMBxcM9Yj
o7g9cBuFWYdXTmTmUSnHxDs6CYE/f6W4rDvFrgI7WPSh+Q8pCKPfStN4MA2AJnCmQddz4Pq1cFEn
RZ7+UawHtHbRGmdJiXpg6Va5YSYfDoMpEY4zcfkJGv/8miFE9of7X8aXlg3CzMtZZzB6dHQw+cI0
smkgjD+34yVem5il9oajouHcMnt0+Kaq0hLvfaG/dQDTjMUU0PpFbnyvvoMi4JUYX52U6JwxkRLw
xhvLm9L03ucUAu4MlNfirEcpqYyCpxIb/iCR61jG/wTda8Nb3Q+pVbgpubgqXl5xBVD49g3eJtEX
lrvpu/vkWtY1m8w7PUgsdgWSYWGY5rW/+ypGxG2J/kyZ3iHTK9H1rO445dzUuCb8EnZFnEO/zP/d
65KTuAK9N9YhrzgHm2wv8pvEhSZOKCunX2p7A1GbW3mx83rvitt93pTDoA+NdEmHfG2q5jaLiKx7
ujUEEZXJkU+2me+uNYSpZHJa7MgXPmPNagWy8/sSSH8Wvj5HacI+9R1u6217ktoAsfdr4dOzF9/6
yAgL0m1U5EyUxxJfplfdD1p2tT6OJn/u4+Vjn0GoDYIyuxn0uoWqxsQxEkxBmwnRkNzPOPUK+AFx
8Z5QjYE0g/9tmkmK8d8U9LQwJ0E3SfLDm3oCj7BTGUJEoeBlBOCX0qyUD8j8ntAS2kgSlQVfplYq
3izsHAGys4J++5FRViXNkapyOeTOU+xE1jQfJo1p/NkCUtr+nJo5vV93cCW5xE0MssJc2GqDOzUh
87rFLlDS/OW6sudSEZXJslB4Pz4ACt0HN+Bl/9fmCyo76NZpuW8Cy03iov0QWFcNM62zSGvZFRZb
3YV4oQ2no1j7pkjpocF4u2Lo1kxflsG3zUNF9w6TFDNU7IR3XaUpVH1iIxYnZP6BwD129rzE1dCl
7PZ/x0jd+AnSXzmMxwBEZG4GuVIW/2foihsxqZBV8vDrIiSQjT5eNwOylqNvnhAfWTHwNOMgRLxQ
OvOsJn+HDbuvqu5Dj1Ca+WUCPiYTzdFbk7w2yzqfZA0CkMQJhHsdf2Jq9DFHcTEyDIpAHueNgyvM
rzsJikaKpSzh9pQ96nno3VZfd3E/JZGLZmhQOyvPl1fbN+ihVkluROudCcJfDyScLeT0Oi5s3nBK
KZptD074GdE/FO3gW5OC/g/4Zxt0Zh8Z0BgbCgGAB7UMzpict203YoWDMiwul3RfhylVO1627UZH
JVE48wW8dXv66Atf+r/fIH3hfFjrOWKVwIP5qA/l+lLJO8q/MVCpYlSfpeIMDlcy6efm9a4BZJ5o
ELGqQt/LhLNO7Gq2a2NnQ+rpJ9b1m5JdEulopq7bS/yfSu2/wDQV4IYDvGaZ8Mgr1BP2ZlPS1Jvu
3y/EjNduQW9EDB5jxdPQWCV9njZmHO072JHYd/N+RSlTccWxgl1EizS0xrexPpBiFgveNGg6j6m4
CILMsM1zxpPVwEd6yImKt9joIVsRY0YGdzh1yLw3CbcGjNf5r8G4z0ge/XXj5tZ27IHPCoCDLgOB
KpOXPTxjnrvTLSXyMThjw5Knekmna01aKQ3q6loKaaAIrGC7rxnDRwSwQYNAGZWnh7kfG36/tR5s
pT9ILNtLP5orey1j5p7aKRVt2Ex2JxCy9L50Fw8p68WNeJNXS71L6klrxQYlhc+B4tRy/c1J4rTV
uSIwrd3GFRcO6pTd1yFLjHVfVSvasMD4xGK3khQrBXpYFMexYO7QVwjbka07iGGKCeEozeQQirjI
2SyJ0IdsFut82ObJMVxNOaFPBV3X8OmTn81QTymddDz6MjLzB4B29U7Jz2wfzIotbAxZM3Qewkpj
5t5zh6W+AaU7d9lAVvDDRoMSsN5iD8Og2g1SxDIiAQHqMwWt/eWzKZLe0FGV0jw+qnMwNoETnTlq
Y36Fh/YChRFxGu3HSHO2DFYtLSR+6pLUUQ+qNnkembJx851SxpQhRhGfxV207ooslas+231QjnKk
OuIqX+OrWd+D1gTyWr8UY9nDlH9AJwiVsq7Z9y/MJrXDN866jgkeGrj5ZSwd8Lkniud9LpY9QvZQ
uR5KR3941vo63udZd5vo1Q9NeD9rGv3cvZQ3PWS+NOYGFpVjikZCK8/fgXaGcYADj3JgEIJHjJLy
mrgzp9lFaWCIBasL/c4o63GzCU0fIGWUndNgDKRGdCseCuTqRPEfDZW9Y97/Ezul6TtVZEEpB14e
5lXcpRAiVp4I0uGkBEf13JXp+qCPHLg+MDXDXdkZywMmYSvX17D+JGTz3hUicLoRym1ZWfG2a8X9
L/KVHMzcQl2lrYjXLI0saaR8R8HtDXsY5NKuk2DGR3vpDKISTU9xRIwo+g7oCivOmta7hLDtdGwv
DN2nYA8BIZpBCmeaiNmUm2bNO6azirCP5coNaL8wk7MfLOQpUt4gU4k/R1tZVEfxNtjXkFY9aT+X
0OZrpLRldDyj1edDU32Jhk43B5P9rAz4O1ngyrVNpzx0jTK/+H8nR7Eh1T5jB+VO/rITQpH5eyFQ
hEFKdRroV1NlLge7nm8JO0bJ6aaWd/OHWXm7Vs7+qe1HLhoXhjFaXrQsFUCY73RS+ViWn0VvRhuU
HnQsmbkgmC+K6l6Z/NxwSuA2i2Wm1EI+7D5dCSaYRnrSLmDjbGFo28qZne9QBjOWIWHcbPQnFoHh
p6DqFN4Yu+qFol0iRYyLwerBIA/jIY26BW0hEx+ViMuwcc21IDUxUOxvdOd786el0L0eMc6/hSuC
tLbrZ1rYk2f6xhfam8eKctaoEEJEVDzDtfAIoqBKxXajNrSr0mKbelXdmgqy+COXFpNBcRloxQUk
5IUHKbdUfRn1byq4Se768fxaQqEnMTqBmLR4+TkTojwE/PLpANVuaogXR/X9mku/U++f1rCFwNYx
qt3dBWzXkRheb0JvVg8v2CFzRfzHo0XE5c2Z1GCVD7LnwfYd/8H79JsVuX2QjORGzQw6fbOTvb1f
6vI6dwwgyPRIbhqAMwXqvphS85XmK32BhheX17M9CdMzEdcdtkT4v3gmO4ug04jWcuCr40ZjYD2P
em0mGE9hKVSpgOPhPZ13SQlAnKqDuuic/eMg6bDbDw3y1f/pJEUmtvRqSZCuFI02Sx5+QTubQ6bc
zG1Y8p0Gsv/37fSDGG8JSBYaVi7nLr/jzOYiSXbnEelTU7hBIh5WsGoKpE1gBEVoFvEeTj9F2s8U
YeAeuA2JxI0qKjqRvBx4QtUUNdmpXRf5ohBWP8K+FQUdwiZd1n3LQpetpkucObXir7IKYKhLCbRt
ysucHmGvh7KXTZsvOLUFe3fDKxakItfjH7HFMaApsUhFHtYNHEGGccFvPiETrlNxHpT8whbmky0u
hMCg/A5xJjvWq+1q7lVnVQFiEWwP6bZuJnXjTbLGKcEeNLmAQq5RsVoGEk2+0acDslATPgeUnnvs
iRCkLb3Cu8Nun4oEHbKs+JQKqgDWslyljuZG9TGIo7OfxH3up4ExjMoejZshU0B/WATfkiUvhVOx
2bLkKBdgW5DqCDjmYtR/8h4bQzSmkz2ikrVTfCDaC/C9KqTIckDSJYqtJ7lcVXTPN22FZfTeoDN8
OFnYwdUabtgOJO+SUU1F0xyRs+eGAg5MIn4sSsebp3xp+qLKIk2wgYZGjeYmJYYfBXz6D6jaI6lH
LZS9o1g2aHHyb0YNwiQ/4vjhiiMqNijY7RlfOiXNjA4a7D593fJItwWIyny4TwRTXMpGz53PynQw
hYqbuc1I6/lXoTpU8CkumqP3rC9pJSdH3SppfLtJ5241PJAegsyyaATrQEa4rVlWLagq7yMmAoDV
wBSBKaNpMm9oQEdt9VbHkikzakb6lzbmPn7h2O1CViBild5AxtQgbIvvMW7k8L6zBqO8AK+5AW6l
xC9gtmVV1x2exwTVh3jxAQC5s+7ramUxK9jzW2SJfZUn/VxRS2EWMKKB87jI3H4g9bzmfZtzoDom
OGh/MLeYNanOtbDnuoHBpdhcEbR8eJvSpaMEP+Tcjm3WPLXSy+5jZS7W43JL+spO/UqFdibzDmrl
D+Qp++ifWalloPentWZ7kOMt/A9mhD6eAM7ryHW4ZpEFWy+FB3rhlw3kW69JI1SoWbj2W8YJbiQg
MzEhknhzNsbd843Ut5s9OGS5evaPRuxkZmh+Rmy7dRzUYkbbzh7xcEJmqBrrH98XBvPhLhp7gX/Z
GFe6hjo1fB0pPjTb+ybwrJWk/HqmU48rGENNUqPSTYHmpFT5Svd3pCV6sXKCFXWGu55wJHjYCkeJ
F+c+baDquJLXlPw0K5m0K4KdejAxQy0woFo+tZEPcvwevsvAFDEGedx9IYxvN39W84DHBwhtPiWw
VLb84Isvfp7TN2gXn1ptk1BNPQ3vmr+H/FvmFU+W7dnKJ9qx814sDNHEnXFPJsOHjwfpGsWs7hzp
42K8ydCAnkBU/WepuosRYa+aY0r6d/BwkzPKowjfrVdpCneHXetPOjIuxcLtMjapJYPYRaFslOi6
kx5Q9LhHsVaIswh+Si9l355PKK/hR10syEU/z5lE94qNlAyi7GB4KzOaeKM1twI61xiHemcyTIB7
Ddm/7eHmEbg0P0gDXCjKzHSRog06q3jtv5eOgHlBGGSCuA1at3YFeXMCbW5WLOq3my69ZrzSJQ4H
fZIKMMW1MfiMmedmpa8nVrYxo2ZLtFTorNbdYOMt9Le6p4bTF5fXnSVDQLWftqWSFCMrgnbPoVMw
kAlFJ1ZJakK0Rx7nmbIuz1uO61KLyI9JiHjqtmTk7mFAoBfbX5oSjA0k51TRvP53wwh4S99e7GJZ
DgjIQU01RwkKg2gtQjwrsEpo0PnuHogeM7Gf6c18q5RvBOhrMOUY+OIzrg13SHcFnTnUMYmiaTHl
DhZIj66r94e8c/sc1BKWoWUBpGdXDeeGkiRdy/gEqEDJEEOl4eisfusRHAFwhnzhy1HYM28V/pon
aAvGxK1jobHFFuyByHky380fiO+zbwtWuUSOkqwM4GnMsMzXWsdpPNTtg73ma1TAyz+aH1HZGnJ6
hYiA/L4Gk80fu7wrpSn5BP6rxp+xOJoqpjmV4BGgg/PnRELyjrvXfrZeIBGNt1Qua+OuDK1kLGig
dYTsT66r/txXUOzqHP65Dn/o4Jo1+hJpmlFb/LkxNYikIErdLtdEBfDnZ7svBADaz94FO/p0HTti
8kG0vUhbSN1ozI0oVhVXZyr7Z69JDb98xFtBYBvARYxEL22C7/QO7JSzPPjzZdbdkJdqduum+oL/
Lrf/UmPbmDWGRwX6pYATJeIJ8TD51nhXdfY8QuE8PHDWEdfMMAl7dFyX8tYwiGwRoTZenAeq3E+Z
Mw30KWK+3n09deiKKIsE/aEuWACowAUfVZ159r9nbUtLgk1AIPqZgFE4c4pi58+c2jGsD0orFxet
WlnxCu4npk6tbREtZUT1FAkAvzLM+mUinI45vPbVoxpXi8STNKmtxDPQHRdX0Ma9i8oz8ZbgHywT
2+6Kj/pjLeiGnd4XfjuFSuSQSqDsSZAgg4wC6gY9Dd2idZo6rdTvwJsGnrS0ekxLHopuAajVkM7y
pvdk8HWqBsBi9WICYjmL1ju4c3UkashwRDsI+JkCOM6rA4XQNlhlN4/6Jto3WUmWb+4SefFCNvtj
PotuNPSq8RIK/STkId0Gb5bMAXFsrh6k7lWJhJUAzAmdAJfyIVN5K0rUulH+Vp7kvlhE+qI17bo1
apZGoT2DRyIi/cocjGhh3XWY88yrCsKY4OhUz2v1xnYqrmunXSyLjqJZrerJ/u89Vaijs/+k3rfn
dEKd/iy8t/kfNTh8gJ1+3/ZTHr2sVf7ro2iazTwOjXnfhVnrTR0lRh5CsF/Wio0UrNQeIFd5N1Oz
ayuw5bUa7tI54bVm+F3wAnvx3ziaK/6HWpuQDt30JcKQLdGCMYBoRQAibTtxVncLEmN+zVeLex5M
t5b1FGH+lVft1kBdQc5VRQKnB3T60egZ1lIvq81mHEJC0sll0WLgrDghTMTHpykF7eJJLmsHnMtC
4gAot26tKMMY3/O43CS5zE7GAbRRKm4rbs1cRzrxSxAAH0VF6oE6ey1IPc/VMgnGn6Dy344iPYe4
PshRR0se3HEe7lHn9A7eti+xpUIT/NQZJ0nf7LyP8yr/o2gD9XvYFGpq5la42E1Y7YcgaFrGYnwR
MopcCgOPhajA2GocaOobQ7N3HhZH9ZUvRTlywbBUym3Ev6YPU0vg2IBH1apwktmK47tWqW7bo2zf
YXy8IcfDkn2rJs5zksbnBDOIEr5hkoJr4KCRIznQE9sSSJCvgekwvlEOT/nXHL7+vCheQEsEs9rq
8BzzbSIE6LdF/gngJ6aiWQ+NW3bp4Ijj35uh5upLim6H4LKrgcfTAKZTl5I0uSWokPAwRzQrk8UU
lGDL4s6oiuMN3q5Qkkn/tSJ4lCxw5eEZzc20ON9ZS4mrSF8c0dsuLN+gGAb/rt8a9g6SsFI8YSGT
NOT2LQaaeBIXm5a2rLE7CnnWLGG+t0YWSTASiaSPMm2Pa5JBbQUeo21iBfLdv+nMYAK5T3frTbAy
lhysdDNAiUCkINnjjX2LB6xXRmmta73Sx9LisWZ01EkUH8EW14HOAru4fc41SERH71gU5dpBo6Wr
0VvjGSkQXxmqBVxdNhzPHOeeqS0xC21ykfl1M1rGxqlOXAUoXlQixkFncpoZ47YEpVDFcGVK2aVu
jmLsFEZ0NojaefLy9/1Wu/rrjFHu2PekOMU03Yk0qzYJiSJfvoXUgH3uu3P3Nb7Of8fKgQH3WWY+
VZmOJkjmhdqv+8M+w3YqSkzTcEpIcsbfmtD6ctFYquHUbBpWLTSMCo+unT77eEply1VbBVoBKGah
IQvABbSYc5aMEWB8Y2Tm936W9EqDEKS8rpl8MF8YCY5jiq+JgOm9sRMQDbMf5axkhmY0gfUrUoAk
cxQM7ukz+L71Bk9WJdkMClKSwAyldQFR/s8ug7DdsSTpokhYWSLOV85QAf2ezDZDmtDjR8QPofMv
zVWjb6SzktEAhMunhe2xvuRtQmRn+zeZi+/EWYJfzRrI2iUp2Vx6JD4V/NGVpFJNyyY5yWpt5Yc5
9mBfi6nvveCHzTatl5/ozKmeCX1K6tj5E1TIR8cWUM0D3BJWaElp22RWO3C38UG/Lwbig/tZHMM6
2lzy+I3IHv8u/GDcdvnVaLtT5AeBMiwsT3NC9U56SM4Yhr8jO3PxQE3liYMQ3/06O2q092tP0LeU
kIoZzbzgvKKPeW9zvqYjaJFSenK0tV8ymyWfUpFlBncMoXTJ6GfBEpZmH9x40hCaNVHWYnu9vtYW
QacsX+Qhb1o5PVzQOH8j0MvbbFU2e8RiQ8YJUEAaGOoluu0xvN+3diUT0cmSQ4HmhyJEkvy/aFJy
lzKlAfMne5MMoHC54VXBtCQTf2mkhsIBaCYp523noDF9qxFLc/JKRJYPC1p7mCwdibUFJSsnVpVX
IrbYfsViZDteLH1jwDVbhXU9qKJqaWGtmWnfKngE+pnRss+XR3ET9ZM2csk2l22mGjLnbLvcz1Ea
mhVzHLi1s5oYx2MG4FuhqCrPNnRhO6yHIp2PL8RyFx1Ph+GVLdVxD4PCZwNL6GE1wHNTz4OCA1CK
YiQ+6dnNs5G9FTjgnmM39/TrUL5iSVllOh4rynnyNYY3ieCLrRNG39ZzT7AZu/+8YfuxRXHgPGjv
56SXNeIGL4IgqQilsMVnAkgOmHmdB8FRt4fARiupr32m7v+wgopWrgomuT6XwlgpcBjSaK6cTGUI
riqeDpqI9RtZCK0S1caMAzLiaXlLVmUKueiB82jOfx8a5tyDddMi3Ht0vdJHefh9NnIMaS0ZT8YK
DZ7heYSeqZp01QXdYhurj7sTkvSVzYmDjOki99kywBPXp5AM4O5S3mOcYR2sCNPO4CioM4AHLLck
BfMZkIAZkD7aREITh30T8iBC/l4Ocf8OB7WtKAcBmJsOXi46JuTi+ufQJ7U98g5iPnV1zLzje6S6
nYjMtpTXpm78FzshcoBnieHiPimCFL6fDgnPmW6Jn+DnVQ85ExsGsEbUFfZl/5RakxZb2GSHsGPw
tABUjFbGH2Ew/sioFRwEJu1a/jAbYvf6JwWJBnzOOIGBOUuZtERgY97WfEtssJPkk5SKP3Hx0mkp
kL4wW/RJXn1/ui8Xe/fkju0zFotkr5Vm1WlLpqylJwZizO6cC4d6H57kTdfPRov32z9UCq/h3hS5
wysOI5g1CjrvGVLZ5fnw660n2vIUbL9/ljJ2usW9vUmdZosbBBQAnVdMlMkfmzYJDAABdz5DS8uD
ubQqoTrZRszC9esYJ3CaVeJ220kUmtJy3XgYT5wl3uckp7S1jZ2GVNL4FBhiIg7I9EYC6eN37sI4
UFTxVc0eyiMZfwsQpuHxCGko6XafJ4E6nfvcW0Fc4LMl000o+NF2KxA5Moh3kudagtm3xdxQ0XF3
jYDAMi3vtmCWI7q7+xIqLxd+xR9ufoLwZEbPxdu/6AYn+CSpr+/HhfJPKhnPrhwoXFnVyyhBYw4M
hzZjMRW8os+Ilxn38xC9wp1QmyfwqlwcqU/mB/j+kcQaYnXNrJsQfJfgqlepO3hLonTCy1sZs0Je
pTuxs9cy/YMvms6N+Je24WkikUFOj+jzdZyZQhCLJasYnSsielis5G2gP1rlSoZzKpDXSZ5gIIFq
N28SdJyJQLi0PLE6uKLKII547qIxqebshAjrJkHF8lCYCNWHep8r8HmyqtBNOzBs0yd+XindVaT5
hXFcY0xKvZDvptJEfwHB5NDgP3wL9FojadksWffQ375tHvbyDi7yEzWtXdhVJjqFfJIW9W0Qg6I2
Q7OS6i5U9AELJQppVLfw5uunyrNWpe116pZerTWEquIBtwufff8BpYNwczBxCvcqmMz4RYlg0EKw
fSTpcykJV/Ka9+v+3eP4hx61/RsrOiDqBNFzH/ASL3eG0o2PjYx8UZz7KYc3utkUAWxnhSeLgDQM
OhAhPlLYS6e4BBxz8amdBT3qTskZfzFVOoMrf4RWyUOsy4TfDEEhxYdbOEQp71cPY6lJLJTpNBZW
hM4oXZ0d4/T3pmsiAt90/WfWhDzqfU5wm3rSi9XE0LOYH9ThodhrGTg0k1eyf1M6Y7hGSmTOcUsp
sWBtc8F3IgBx/A3Y40XjLlK5tA/meEqsVdQLx2n2HIKQHEpgJGWBAlwXz05t3FMaFRFE3x50F3Ga
rIHTvvGIqrY09KvHKfG2XPy+qdbFiqRZ7CD0lIBcs3xi7z89gFQlIEXDYDoq4LkxehfZVkdPbqfj
U6waCxxgAY8c+6VPrnCA3F66AXg3vuh7n1Y/q1xxYInBcs9HOQtgCo2bCwJeoPhldgvDaA7bvGii
U7g0L6+syjEyjJO7+Hx6uzUtXmQikLAyK9/MDvI1JIjG7m0upNiryn8HgcvlbW/POkXHBsMuB2xJ
MC2dyPuz90vLmBQgYpI0TAWzeW7Hvk7HwG6/3EQdyHFBu/RV0OkTgG5Lrt0djmq0RloBJkxxvOuf
cfULqSUS6A9wzaApJm/BGYNuXDp9ym66o/7BJIt7Sf85Q5VxRhtEsUBxFnWwW1U3aMzOWYAnsfO0
zeKwbMhZWzP4oKhsWsk188JYrcv50zTkKSTin4xm/0SXQN/MGvOAT6DCyafn5VLIl9PzDSAGmXle
oanWI+PhFNEJfEraen9UnO74mWOBKepKt1XvTdt9PAWuJi+XGyfcTbEaSKxfezVZTBkdsnfFpWpY
2KjEZDJrI2kOEHt1H2FcKqAK8Qfh/y7XykrOguRtxzLvn0udxbOhBgq9VMcYjbMu3YSi8BPovLq6
zwWxQP042OLypiNLwfZZ3JFxcBlOYE2qgRPdd8DOgMXxEuDZGTBj0yn29XsIwav5qKQtnHBAwM8b
G5S5QKecD+ACzTJAHP5MoGZHkM4wZ20OsaVuPMJbnwdlDC6A49HoiuAk5+bAw6vNxPnH4wXM8rOd
9c0OP4jIr6AIdscnUXXanxAEYQdJ0AiBt98N15mcz+zyPKcXtKD/asAJa4fW+vuGJcON5wBe6kn5
co7+iMp2fkMaOQGEJoSlvLX6y9CquzNpm/g04neYDzAK9HpC0YLu5k4yiTbVfBGYRUqs6wMY9cbx
/I9IucUmyJKf/EOJEFbBr7ivgTaUcN8fKutnh783+sSPLLTOU4gPfnYJgHq84VQHRK+nS3GDytch
JoYtkp++VzZEdn8Jsl0HBIHyTwHRWLCiIazQ1J6dNnUQoVonaaneHs1S1vtnSkqpUBsvg6pxdTVv
3LCUm1vjbwfQfHn/oM6psLY2T7FdJK9PCGpJx1ZwzdyJ2k5/IcR4Op1Nvh5WL+4jig2fo5NkamYo
L6vw0ahOyGDAGLzF13gNL5g6Bb6shWrSjospGgHyr9DoXdCIJIhuz16Wkwj/KrcMZhpW+w6wF7ri
tlaGL4NUm9B18H6ArOCHVMmQMAP5gewW6uP3c0SuFpWj6JI7KEBPRrNQ21GPTmCFPav9QUeOfCdN
SegTGngQ91Rmb8i5fGXXhpGL3+cIcdNHShEtWjBC0JOudxxaalWBAN1qZa0KVayNzRuGERa3O1gW
xerLtVQrgVNDq5ixQLZkFRMfoOolfJG5CnGB83iCXfPkUcFj9/g67DzGaLFnzZI5f2mwUOpkmPwy
nHw7rlfnL9pPog6uTu1F/xp4BEoGtrrhMn7kniBOfAwfyKbdXckPfVWnRlRZxWn7LCaA4gyMrVCM
vr3DyGNIP6qt2/UCDDaqrxqdZVFBIWJKVdj5saTNFLB+LQXpilI9uZQcvLFHAi+GCjn5pxoNVrEY
NuCYZ6mu3WL7qA0gGfzqnz62xQ9lYy44dr8HNgwkJNahTcF84rgXs08h48mfa6xcCadOiGgP9wCB
aGf4UHHKIpVtRKJKlEv3GaIYay7sk8AF8jE0GUJ34v6A0WTfzlnW1VS74SFd+M42Jnr/M3O/RSlx
9Z40cCdlDIkzr6+jy2VLjrlAGPSnJkP7DnM9JPxaRtaOKEkzhp5ioaxdIzLIjqhrDvrcG1WLcp4s
OOS+PZutuaIT4hhlm2Ss/W3z2xtbtZIsiIPigQOsQ+twQUmumKL5IM7Ww2zAL+DQRH6h8kSHa5P8
eeyYCR/GSNFdQm8DTXZzYoHUeSvU2a2xRS6kyt34zUdgO6bzhYrKiLEZAbq0cRGwZewq5WwLgePu
5e/+ZcijgFzvtEJUhNzWrVLHVbpnz7mfpE67cOOdVIzlB0mZA/tSMHFR/WgEwn+xAIuhHIcKpySV
onOLpEZP0YjAFR+AS4FjBZd9HurRj+sSA695cve48qIcHQf1xdkVCdN0l07ORvMZaBqnEk7i2OoO
ZQWLRFEwMDED4M0ZTWw3v6gFHe9SSYG4FkFbg3QFfoHUGKdrNrjnd2dTVI5A4ZiwFv6yAi+F+bVB
rwqQBK2asVZ0kVQkdLPMU5l1/02yhcRcP5zIl0VJsWFDS42McXpzVQtgNmoIy4UFFA/SXWqSLYhl
1D9OWTpvaYRA3umG3aj/SnjeO2H69/5lX9lm3meYWm5BSpzOdXiU+xeAWUEsGM3THC+SiaHwym/l
TJJBsIgkWsYoqQ6iG2UGOlit9zaS6qYu03XDNy32RXI9bWyonD6KwyBq1spjyERpHz2KtdDgMgLI
XdFOE03Yh0DGEbm9q6KWAVOsZAUxGd+W+or1kPE4xtd/mtTzJiDSRGR/WgFyL+DTYcSa/uhbnu2C
PoBdSkoX3ZSdAm+Hak/783CD4Zbv58+Hktdk0lqgkPYwfeRujXFyn+eCvvYEHpTjPtAhyOvV0WVw
sc6iw1eu0GpKVfW5Cn/WdjL6BEyVVy9CRqiT3T1M/VBtxSjxc0RKfv+mLNFaeD+2yNryeaxx+wJV
M2Bjby6bwKpRWI4BBLjwiTWTEizQrqZplNhYwDrzmztUP9xCADagBEZpBCw/C3lxW5GXZnMmqwdK
y+C/VVeRA0JzPxyznwJAYI7pV7xfBdElVzRXf7tjnrT5coEBsCeHrOKQHhXxPAsOVdTA4EbF8hoM
A+WIG+GXRvBSterjR0MixJstqgLdBT/V1weGXSJrlvrwy6Cl/Fvpig7L+wymem6VH2/7BpJsDW2R
BT0ccfh3vjJf4tFieQa2XcdNfvvBlJOivy0q2DlrephCYgLIV8/dqPJ3wZg1FdY6FAVdgEbOpiC7
+lP7YcWzKHQViRAA3RVldEB1MgCFIlKtUQv6Jr+bKkpruKJHUlxDXyTdb1MPRLYNplPiAEQZIGib
pUjaBagS9hFfiCXTQST8coEoLgbBmwlImu43RpeftLrG6iJmywRq9gkixN5Cp0y7Jvn9GPUuZFgT
Lg1Jvmho72n6xsmDtHGuR5oQlVJtSvknmpsI/zs/A4uiwWw5mVB+pkd+KWhodGHr/dW+ZbhV95ye
GFAbOe+6Gsf+dBDhpoAayru01rTWF8gmoDaDBFby/PCMXZYa+PLdm6i8jhkcxr8ETNz7XudonREU
XTcI0d6Z+JghuADjMYPvD/CCioGwIwvIU4NeL6pGmWRsaXa5Ie0CIliXr7xni5SAKsRpch8xtDQB
2iGxfd14DP5zwT2zSu4yxXyz7m8r6cJDAMq7NR22Gi72HfgQPpsjNDXu8Z6ngpBVg6MlOW5eXd+6
6u2B0S6xOJX5hiyHeRf+Q3xaxQEPGeobrzCbkwopbsib/0uSJbL++rU/EyBvxQNvZC26VMU4su5P
PFbDw5vbbUJ0HMdtY3ywwm4R10/b1UGI9YUrG9CPlOnn3kQN39yUl4Kgo4n1u6Ga2TbQyJgbOQJO
lZ6KM0TwSymaIh/f4lcavZbig6lln7JTtWItf2ezZ4pRn0vF5VywBrbQ3vk+7sNP/RK0QNteby9W
Y/rPDRWhaxMhV39rNYZu6hoLZY321goCv2oowc820vZ4Zp8Xg4d1CZMDfooclub1y1ldkRb0G/y4
9olV9gBxi50Rwpt0KvQukofxyieleud/RqQIlCoSQ8ogiNYw1wE3BR18O0cGLsOSeJQhzAMmJUqN
RT6l9na/s6rB+Cp7ELeWDsz8KVfBTmHSSS87jwul7QjOrRo+HUX32nduRnvbzYpx6YoOMw6ekD51
velqundSJ2rL75MmsnqErmjUopgrLWuD8ZTvskInGw5g8WgwLan9h53woidVeUevv1J6b5nGGLN6
hR9slDl5Sw8q4a/8H9oVim3hvdwo0xsJsBZJI9VPb2xksUNpu6bWtlwnV447OTpNe1lT/o6OwCIQ
BUS8/j+hHbFJbYsriWFSGQVpjxYgEKbWA0ivCDXOKJx24XST62dj3BVccVPE6j1vYL4loAilMzVA
78EzNNPzM1QeUlYGDjRXKkAlcpgAuQiJd2cqRKQEt+cQg91j3smstM3QB0XrNaTcQRj22tsXurJx
jE0heto1HcL7bDJy2fK8QCRXUr0xuv0A8YJMzQbSKHPn+HT+nwWseqoV98NQVtRvTLUSC8qj64ps
I3A1KN7gJDIloUKARva46K7iGDXvfZD91dQgusiPr4CbeGNAHqQ9ADU9FXZSp45LJTE6oNe4QTyS
W/WwYKyO0WUym0BPkNT7p7Dkr2JeRYaAmse3LIg8kiT5Ka6R+xtR7H8XxwQrxVBF6kaVY93BTtnY
WWAl5dIW+JqLeIGOovUVBJ7sinN8I78dRFHyvXY7q0nZZ7bpG86J+IL6EKXjXsuT9aQLMIQbf36x
dTHvPBIYXTBy6BP2v6nfOFS9n3BjEJgwZ+KN2hXoT0DH4HrzmoIdFef/X8FzC7q9lGfyBIsuo+DF
9mYT1vs/WyeZoWKmMJLwltvos9DtS3qNTLdUvFbGOIoCtdLxyLMU5jpGOIzxKZ05o/IkB4yhUuoU
MjbcZMxpXX2VPvOvbk9/5zWbqo02/TItIXUiCUTnGYrQyEyNyJb59L5gsHpG89F2POMHiy9q0Cy1
M4+KueZNltKYGuAAyStrOEF36dtB4Evo0jqhf22XrIPSjumQcwc7Zr7qHxVLPYxxJ6sjhQwVTN1E
Bn3vKqOZ9kvZmtLvqMkiZkiipkRaOEB4KIKfuy83UggVKFYqTKaacHihleWMBCfsMiVDceV0IDP6
ndVt8EBkoSYhI8ETblwNyq44kTYV3Wy/Dr47itoCIf3S75DqRP/x0YONQPSKKa2WbNr0Bl5QAOlu
ydBksKcehZ78fK+We9p5Z/8rceolMrLWiMwoUGT7Vi/248J8tkqshU8XkT1svRupkUTNE27oaBwq
Mbovz47CUrrPkOXl7pC6cJHOkhe2YF8DPc9tQQHH0//DKx4mCPUOiaAHWOM4DNF2Le2PyAvy98hx
1RNoWQr9FQW/T9YRiMx2s4Qkr5ZO2U1FqUebZx6WpTfaYtjXluyBCV229RWMGnudXQXk/sG5Ifb/
74cOqFq1q9zp7noXi0XH/3mlT19muqcEkbxO4+iRIWZKec4KmIzCHytQ6x2PARDWJNlS+KGt4ZO2
oy5BvYOIrvypI6cmeoG+wR4kYuReEpfTsZ6lp3pX3/jrIGsUv1f+p1HXH6vCQH+3KnxWBTvqO/WS
lfCTLpp6k135ZZ9jqw3/AKS/goleRbdTqaFf4LYM6aAR4lGtSNQMYBth5RHhazkls8CEZLMomyqm
m0F/OuG2hkNJW/LufS53xNbrK2BLddPFn6Vkb0/3S5HcG6laZXQONXh9U4uPHCzubVxc5LuHHr/z
9xQkTmGqjOJ6XylWMBXuDEkYfX600Tvbgfb+pSTFtpvW1EvQEF+F5aNl4i2uYtNFG6lN5BSC+xaM
B5rLt1Z6LU1vwsD8GvoXazfjF1TveawMF3jnaT2jInaMd7/tHmC4H/ScvCZ4BPwt46s6Lwnw9H50
jPxpz6FrFq7pHSzuoYInjTmdL8iYBfS8W8o9gYE3uIq60x14Xg0uMgilvu1wvhKcuuZZsg1p5Dbe
NP5pOSyFAJZ/ePFEKlz9wTUGQodFqq2vqTrGoJ+Waz2p70jMs1MnvytpJ0vcVei1xE5hiuTwVwdX
jDAPIOF1hMh9LDdiaszRoD9ZL726QimaZWuYy3D6UAQmuuJG2bPR0adwRBT+dR4hvqHPsx1YlQdh
o+3M1I3rhBOHn4oF5Hs16lWlz0mVKTopTb1uy9x0A824nUKp4EW8pF863nVTPGOWwzMM7luPOdy5
/aqqAbQUympp2e+xbP0bx6agY97iOsSwP+EUjdo1vDb3Evu5BFp0ISURQ5vvWujGKxU04qeIttKS
I73mVJBVTkVmtkRFPx+BDv/oBuapGI/CWgUCYkEBjyacjcYHX+1oabbeCnTnD3beglO0SP0c7PPO
vcrSPUTW0OfMN4lnqJ3mwRyFNFMm1+Kx+pH2Ei+p+F7/RwlvvPNZUgrGVOJPQtOpsExmV8CkOVWf
D2XorvE0PrWTXAi7/kHqPdwD/GXKIj6bn1GtpHJqLZ4p6IY9KpOTj1reWfBUvVHextzeYO4w+85x
0kAFmJGB1t+jF3a9wn6XafE41az9UKDQHvPlV4B1jMzlGKRknZmB0xD9jOaKFe6xiQ9wm2/MRdSf
93oxmjieZ3/dLb2+bft1QCq1fOvW3CCg3AjgCMDALbOExHYmMK+68a4tx9Cet0SxfVwts5XB5txa
QCdKHSWE7eS7YKjIx3KA8RzTDYAosTPtzGGcsWhLyVZsx04l9NZ70ykXwa9eG37EMb8HbwYBGEVT
R4rSqUnhZZ/BXkBatBraYCxNTGVUqoO6RtVqOIms+ZdZqEBQWRSRSlgeAil352J1TaVKirnI2CGm
lXIypPbuzc+rduFCroe2x7wJPGv8p1iBJPlRG4vYzTvmPB63/5o5TzGubhneWf691FaUi1TTM76Q
Edl9WfESKhG1rtKulOuOxB+GkZKoqL1MHaXxVvSGler8w3VtDmNElWxRbU7MXYlpwUkS+L5uwghF
EaP5G7wKN3YRXqUD17l5LshdI5QuwWplzmemWcubyNP4E/0kgl6GYWBihesZaDVZRBTmbSrlClWL
fdoow7r/ThwXaT7DqPnFP4J+WC79zRae3qvamQAnnKYQhaU5LYnffoLphDIl0mbY3YS+GX36WdYb
R6aqjxZ9ZpL2ZG7f1NXKKsw41CwLe8DcILUMgjDyekfoP/lhJYzxi6ffjmk68ULBcTkTXP/+JLJT
2OX+09tUz/k9kgEbe4s5nxY/ZcNjbUrUI1aPghIekJwiFy8I+K8F0CBNrLLbPPh8j9eB5xebpc7r
C7ZYNYUt9vtJTMbniqc8TTXpVZpmG+TEJ/nTgZtYNESfCIQsjl9b66Riq8jpv3O5jiY9psF8sx8e
kelfuL5QUXmbxDgsac5X8r9ofHx01I0QGu7oEa/dQxNr8/sdpq9TZZd6wGY//iEG6fEM8GQCQCHF
MAHAnieycFwX9vGCnqmOsYz4f7THSezyezM5uObN+yvKiVdlhjbavMEvSlXkfvBFtYXEk5I4BQyJ
z7YD3kF7CFfwYBafKWU7i2PgMPZykVMDgeJGkMuc1ZdjFTThj8PKngU4QLxsft9U0HNI4x9rVNWS
dCAdPbrrstrYy9xxkug3SseQ5Nq04jNhYC8WzF2A3uOwmOCyEm0IdXB/715yn6tZRu+ddKmKw07Q
hpe+UVSzj6LHig8aXaWjnhqqgwTeipdY9lkNxdIumXcD06I+iGLYaQxdDqT1fRwB5oSlrBk+k8ug
Bzj4U87aHcdm/Zkqxcrg0bwu+Eo9k2Xwv0s41ikzAw9HJhFZlrczj6sDWKcFbXZ0fWjB1LScToNy
6kKzeu3ivCDMU/TJY3fdaL8CHPkP7wcx9el4vr/qlSiejRAanoaRlyUYDVOJ2Ivu28MQfu2BWngv
NTgDYzTfwV3QIiuctYQJRIDrpK5cF4BlqBW75+EeU2+cewWRHPiw7ti7tXkA5a6Lc/dmiTkZLUuv
wVUB6LjIhnzL1C71E+prN1C2qdD06oZavxV7aFoTNGIvZsNbyRG7VvbWiZwLNhf036ZHqZUMjud+
zpz2KawRL1wZtNZe/szTX2y5Bs2BgY42/yuAboAx/oU/4NGhVlqmGx4zZvAoWitFECxkwS2ilnur
+zPhOweBOi6y4KI4T/IfyNQpLg28mK/LpP0CB1itBYCtqcB9yU7RM1H7kFXh9Y//b+4AyqpwvUve
6LcJ604qDDJZ09jcX7M32VTiMn780WH4RsuwBRIhv0ojxyOZR0aC79YENPkGzzlmgfRu9v5twf1f
4kFqsa2t0j8+VsoLz604GNM32pqZZX4vtcUKPszs9IBuzn9ccsDPPrleO1cxWj83a9LtOxeurSdE
3k2lVm57FVN8Ah513YlkKeKX4Rszvky8UnSnc9vFJiqQ2ZGZRk+GBaY9SYH8mkJCNqC6PcNFikgA
yrS9RDqsdXHMIFz8CCsB77j9XcBftAONEU/0dHI41gXaON7fjohAUv6J0yFL6guIeridiwbsMapH
dla5y1biyec986OXj0k1XjDmMKP/IRVhxwGGRarnZ6Y46AztmWf+dQ6hMsPJKNjka0suP0fRSJNH
UbHI84FFvCcCM+d/8GBery4fdwbgUqvWwkkgpWoZJRhkICjZ7bG2ADYyM84qYqjrbKAjgn7S+QI1
iL52xWMrrKvzULJngExnxa4YBT96A/CD2athEZhANPuURyjgYJuQAS4McTk7p1MRdxR4EiPAaga5
dfkC8pFJbNaJz7GH5Bd7s5gMhML56DehZSEbYrluTh+pNDk074HaSY8citNGlIHYmeXjmm+xUDWT
pDVQ/ECvmda/v3dfcQGWjMlF+N890oh0+OS8TIsxa9dXw5mDtJnwIH+debSc6PSga4FQYE0Y700Z
PP1X9SteTjPpMT41G94lSJG+DSWtSrMuUcB7zrBjQ09nm3S3ETTqyoXYYy2t38vurK778zW+6pv8
BOEn33bhBWjcHUftXDumdVsx/iQ1jlu95YL92DpUggtpPYiGRDH+eTDQZU70hFausU7mKWSb009n
XgnecwThx79rotSbJDhocXnRN2Uzb9Yx+T/EU9mlfRUBWbo/g1UotlqUNHx0AtJi5kl6ZYTlzEXR
cdEWynFPP2QG0ExY3Xf+eE72egRiGMlpr3AjkDtoeROVZiGMVLj1Rp4v7BaUyEcGrS4b5P8om7tI
UUO/OOsrYpFPfItFFEFz5lkbqLVSgTnOW7XsI5fE6/g3FXd8lZs4ADjEZ0V6o8GqZdxhZNvsvyp8
SiQ1PzJNoWjXrMH7f/7nEVBRkKbku+ZPgBdheutYNTxC+tccIw21byAeQN0x4Q+2FW9/maCzTM73
P+5slquoH49v03zFD3/vuUn8b9L4u4ktuxWgwU5zX//KFNPc4bU9aRJm1IdikujNp1bAooDNOkoO
28i9t4e0trlJwQnBKpebuOzaOZOibVfSB+NFNqXH76XWOYvkDVpbCaH6sYwM7ZwppM/7brJx4qg2
omgZYRmTHU8wel8LNygp2LtMPTil5PG4B8DcktU3hViGYQ13yhQljb8IMLNGQmjwpbbpjFzCfho1
04DO/wNIT+aoG42c14AHoQ/ogGUOTvdkUpCGvBv5/LldPK0nuEfAR39MEpTlfNTA431dhWMV1Y89
mCEZQMHHlkv5jm6vHy+Jjd5aWRJz8kHhUIlVp1/B4WtdqERG8r2sUEuwBtnuB+n2kMGU3aQkvYWk
SYFkUzjsYrcDwYwEk6YGqtTe6W+wduMiI+vQU9fWyWpAqFnCw0/cLLrc+NkIY/1gl/U7724WIa9r
B1hKcJVjA5TstRKqqWbZsiBYoQQ7vQj1o6g+4754XM6ldWKNGhnBURnnj59OATDpsBIEy3oHV361
In6qcrMYoVWuUHDqElTS+AMGNFKk/Ndrvi+S/Qi1aikS2/vgm9+DEY+oBGCWTtq/2ibQvpdkWvfH
8e9/bMZJOaa8drk3yLOVZl+EYaK3zSQHbmGr9pkENu5TKDlxYGEUcABK/pYz6p/6+N14NYxzAXWw
Xm3T6IEbK6pd8hKMSrdrehrwjfFOOaCSYxggdj7Mhx7LJxUcyBBTxDJbetDzWb55Lec1lRtNFAPy
+1VmnJwOidFjaZLC23EF5FDzhK2WleLmflTNeTUFUQ53AEcRSRuhUFynkCgIXeIwYlQ07dpx1HZW
AxEnzihPPZGJ8a3RE8IQCd2kPfFosqx038dK3XFw7OtIJA/B/hxjG/q4D4vCHq/mSTch/2ulkqZT
GF2gWC9v6pFwbq2i6YMKzADgtK8oG0FvyXX/TzM8lzo38QrfMHtljt1s+SDNXVmv0kjCeBo9Va/D
25ZAq3jAPhG4B0MXaoho7MBcoQjyrUVVpcOzczv6B7xi7mo7Zbv+S/pUl/Tmt2lHzLx+riqw++/c
CRGyWjC5k8vlkZjXt5BBLgJZcFYcMpspKFTe5Dt3VN/OdGQ+q/bKnQGe82hPCiD94sI/JX4wuVKH
OpkvZVyTiPltTA4doOztwyHS1AKyipr9+HsfBzEkspyLaIUTrKe8uKGRdIr9X60QdOSXXrrjKe3i
JBstFun1eM+j5A1tn7KP3rY7ByyMmvpQ4+aWxcFLl04z7wB9Mf6uQ2JjXYC6f41dTVTpUqDCsZ3m
6+FBfnkOjS6k0xfIaEvSpxNRgU9wxU1EvjB/XRE88sOarX9CmtFv0ZLloAOo+b4qEW/166lnUn+Z
f1wr0OE0hgMg+j2ixgFnfw7HKOmGvcb2zo456M09X3l1YAo1NCAZtWEpp83em/xEJOGvlzilqZmH
16TYcmVnlVrqxI5sOzd+F6BZrBNlnpWd6VC5ivmNPO+7U5KfhmRUBzXgq2Jr7x7XPxDb6N6TggIt
Z76DkfCwjNuf3nw2JP1JMtMKRK5iL5cCuD7LOd0ysSDOrub8skzErlg6Xp4ImQ8cZnYEJ49hY0xY
FEhGuJthv5wIkHlwNuqNio9/ZSe37nnL4LejP2HUMT/4ecX2r2aEh3RoaKobJNAY/iJw27Dm2/91
WR9Jhwc19BZpxS15Hu2Ko44i119XG6UlnoJRpbz1zQKk2v3NZ9+aLEiZimzR5Ls1j0EZpM+FLkTE
EySGTAWwd5epUN1pVxU0CcHmmtbJzchl+YlUemK1CD3PxkYpI0UdrvrobqzfIdPF+mlGCdLQVfdr
oWJShn6DZMXQHXIY93UWOUU3CcqQpGxICM5pMq6yzwBYKCV18MKjVW1WgEk3/VYt1LjTTk1rjkAa
swLoR8yUDntv4telSHKDBXt6is5H8e786tgqN87LICbfq80SYOStEESoEhQOBu4q7/DPVytnyi/h
xX5y1utKHW3z6k3unMLX/fZQRB27s5Wg9++ka4cnZPT27ea6cTzwPoIVZT3f5N1lK7OZqTgi+q/l
vFHpYqyVKzt+qUEZhMqC8zYieSjUz2ytVSmEqrn7tVHTZ+ebe84LQevBxie/dHB/bUM9NdByToIg
60gz4cDLD3jkXjRoaJc/oU8AAKmZdvj3nRtMa5a4UDW3bf0GJdLonGsZ601k1t34skld8SdZ3wba
iSFwQ6oxCjNO4HmwBMKQmtb/Ra4zKw4gSP8/hT4OMx4a7skENsEJVUjA/2SYTi6m9HOwza8Ix5pQ
zIuTjz3wy2brtNAHbVHzY7kR/ZUzdt1xIoJzfDt9l8LxO/Fp68bbWnCOqCn3xbjjjApjgrK+eWrG
ovGJ/hfK42frdhllnaljBqTHQkF56Qr/k6kO1p9DCTMIIS6ZEHjxdH0GXgRtMXp62ns1tgkXIMq/
r+Qr0ezH7ib6sKgWB4NTYVOMrElWlfEPnoswB8ofIz0Ggjqmtc6ACnRGYkmAQuufRLtyRSLfe92m
cRiYMBlbTASh4ad8f3QVN+bXK37rZ5SjFnUE7mK5tqhBLQQhzozYalM6ayaDvEFdF+MZJl+GOVba
IH45VtZiDYoVUzWri4qPTb6Xek212aW0RozrrQaHgymtzBZM/BCefOwyzlGnT1Y9qBv4e/hPOhAf
thB5Ro2DmyvO2JYK3WnfdpWkOOMTMDM4LuC3nxcFFIgesKxXM9OhfnedzYgUy+qoE5HoCGUvKrHG
QxhCsNrD0LYZfKPhXYPKJCSVqymq5rs9KWfdU6OrxfR2LMmmQxD2XL/k9TV/fWuU6o8CK8JgnRMh
D3w1pghrY0V7fHN15bcdWvvMoaahcuCk3o5fbRxLoJSoxBl/a4Sojat0upfraRnBOHVBaxxAl9RV
X4LBG0PjGtYuWOSo7zxxwMru+yeJ2VPCwU4wxYv+AA1O4hrTrU+go+uy2SGplXgyI2azBcQLT5Zp
Buc6sJTo6i4Zp1U8PyyFUVbo8ljozSUYKpEwPyT/9o6kdTiyD5IhE0NJyfpl4KFaanRIp48jBE+i
G/HH57SSl/EKY/07IocYSNTkA00yxdw3kxZ3Q+JV5s++xODHrHq4LnfJanvx0Z4KpyvgtrsW+YUg
8NRmjUzLD89YHZ+Q7HNepXW4o3hMy0rIZT4gOvKi72PFKF7Yfq7CrpLekaC8bcQfE2TvR2xVbvc8
jvSwFThfObM9G0bbV/y/EfGlT3Kw6iB07TRJhH8i6dGIpAaz9VQyJDlZ6I6l+fYXfii9af1w3bWf
2e/yS+C0jBorsTI1G8duq2BLYq2S1Q2y/E94BFpYCqUEecv1bVwTe5uedd4+MTaCWZamodSM9VzL
Y0ILWEXnfmmcpWDDcH/g/vZbnb3hez0iocPoeYfgpYqsj4aDApghy78j6HFsnVtN0eFoNYzjPl/a
Ue9i8nOiBe95XkXsWdbpg0oXWt/qvYFABJIw9ob1nvJrAFt9FartF22QvmTy5wcIcnuCRsJS/Q8Z
gqpdDqXGfz+np+Z3avqDi78zix1QIkVA27YM7+diTKzFEF/rVoKSEM6eBslGFqyCuCkd1UCWGYEH
rkubBrBXgiB/XDGLRDTT2Fd9y8Wq6bC2N3GEKCoxanbdMC9Eexp6Ywc1/hp5Alak8qmYTa8koTNY
MuVowq8/ByRvVDlgteGu9fJN/JDMYvrkDYMNwC+EccKSSUvIZv8PoXx3B47VilSOuOqjqFwAEOF3
TIUwHYsTyZdfMIg2wrp7cQRs71KX2ZtADKRmPNRi+2/ePCDywgNVBv/gFgFH50k82lxPFpLWom1a
5r9Ja7H9s+RIU/Rl6UqbIe+Bk/LJKWDYuzYXh+BR+jjPlnI6xJ/rdrT3PktG0qQPYFjf0R38wvPj
btscupyyeD422WJ0uZRbuJUth7HvHzZljZhb2+QmOhlFpA55xkRTmfq2/R9PSky3/fQvUFK2AefN
BqxelBhAvDBgsF5TQhgIWJfYZhrAAJNZcGaJ9lmS00VSNbL2bUCK+HUrKDMprRvmeseRSC+5TVQK
5wrtk6Id+/uFSKtL5Nf7XW+zm2F7sWbqvqbNwGFe7dlVmuS4uQ7mAJmYiHqP+WOKHAuxtrNJzBok
s9U1CKD1v/dQidI3gEmSL0YjB/kvYYpk5wAA8CJCnCgOGbJq3XvFG+UbZTtdpkJ5hRmzGZCXHkW4
ju2j4H7BnynofZ6/3HXWbCmKP/KZEhVEIPsEtQ0vYwwqE9FZnlxSNEgRZWTHcLbMDsCbraCLReNK
nglxVxC88/khfX9kOH8mxSsNt1BGK3Sej0bYtkb0muFXFbYjbKBTQgBBJbtva70tAauKC37g+MFx
cmup+OXmEPHdUl+cgMzgOClwwNNzgbjYLAjGE3Vz4bOus6G3cgAD3vkrClm7/i8/FyhFPwQj3b7a
9aEdOV182NXLbF7zuB10D2ALr7LTX1urDFKiNHRB0ZWE0P95lRHEuGIWg//KHMM5jyR0nyoVHzD5
mvES364FSOeCQj2AntKQh6SveoHXcfr9MiuXDndDqiJzJi7PGZ7oCS1OqKjcpFX7FcL/vjf8q8Nu
WChDJyX95e8GMUnuakOg9dtbk6aWC1awysscNi+nUHA50hWau2r1zgTrRrnnI/Ve0Ge3w9DX+Nze
3zBt64N24jCvwDoWzsuJtw8uKg5exnNRWvC03U+qqqoq3ePne0fR7wm4eI3eIWPdIS1pVCOx8wv9
MBym2Kvn8fcQFB1d8Y2+Rstm1Mugfs653wDANfVWg5vNtxkJcudAGUBR8TivhUsVKmYOyZR9JS2p
04YGBFia+jeqDnXM8kFCWWDlv+o/nWllDui8LIRBv3LDj6Q8fIeDhabOb+Dc7lyB1rNo2kVXHEM6
ZE4KFr/ySg39BWzeiMSps7xNCxQLVvIp9qknvuAoQ6ir+JSaKsZ1Ef0mcXoeoBtaq4asjFDHf5Rp
nKBokUjOyigeirAbniUz7KppA5aTf1illsR2MXaH/5V5zYw0AudLdjHGu/biCZMC4CcKwk1sVWBQ
ztdgNu3R0z4sBbShSTSZnXiFgOUHdjQ7DMs9qTYwHRJAcSL8fmM1kuj0fXUPvpReoPntYeqxB5wr
QbpqVlPPsBecu7g1xemOQ/xe6yHP/Xn46P4nlKKxkaowGHDVLSODfArUQolVpQ6CY4gfjJrCBVK+
oAwc77UHJRLsKKbwN4AQ8iFxI8KTvGNVkpfd7kbXSScRUGed4XPLJK510WZk7zYcgL9Eidy6Yiho
hZo2puAYrt4hrgkzDxKxZO8JVPfBar4r2DJK/5B2EziLSW5vwwuMmUEKNLuL+ikSWKlp36Np672s
7Um06JCUfbO1w3VKxORsPTFONvKEL7ZqFXoWPb9dRWj12+E7Vj/NSaFA92WlRe5oeD0JM0bAy3Iv
qJovCHEmoVgGRMhNU123Yz52P1iGwktL4+UyLqS5+HAAsW5Zrs0sAGtTngGXJADOVNcUoRTesQpA
bthbMlzupZpcg41echn9cQss+yL61YQhLG1/hUW9wdwRAwDFt7sc0i6tWxumeTfgiuBrEPxmxYW9
zfzISv+N04psxQAjRnN7654n7HCOjtptoMtD5h5JVxTHQW0sxDCB4JTDpXY6J2eh6mEkpFyYF7Qj
Po2qQdFQNcnNH23sweH0DnXnxV7vXHZjYmq3DL3eZlZKEdUAY4qcPaYU7zTcxsXvFW0q8FqLHosQ
aeqhzuTY9CF9mkivu9abrqsN0HqS7fg0t3iVuhxWXSaZFgcYzzIBg8JsKdeDF3VhcNWB+dUQ0Q9j
Vru6dfxIlgN/4/bjVsgOjrNzTydKC3NlXiKO2kK4XI4kLO4a5epOY8zyiDP8YkBvLsgW9DVxwTCw
jddyGC3hdv3TZaC/f2KRkcpa7ST3n1Jj455+42ce+A5X4WYRMOw/MRw54xt5vC/fHftfimB6u1Ge
o8k1E/mDtwMS6ger9gZ0xPBdYcc3zdIxrrcwiB5hXv5bswC6D5Nqt1AoyayvfYExmm4RFXmDXmsr
+oN7ENrcNZ5KftNhCL/6WsLFrh38jU/YkXGD2pKVnNIg3HpT9rexNyPEoDy+NLqIaed+eF1UXsFE
5sEQZXlT1SnyFNB8D9pBOOWVNJ7MnQF2HpMrPt7id9lMEq0CfHGYm5PEhrSFNZ21mMu4Q5mrdaqR
Zq835v/TNXyLSQLn09ygjPJL7PaHnPsW9IABfJCc62sgWmhMPHv4qf+cgYK0VWz+2JpkBWhqC0X1
ohUGiHzu6R8SJQKs7U4tIpwguLyD+arBNEP+JSxsoWPb8jRQ2UFzz9TCQCczdgtBng4T6iYNFM1D
0Apcnj+MOWbhbwCF297kQRDEQ73QN1vuo/FtTD2FkAsrKjxDoNNxAdpjJavB+MQzTvtPcpJt1R4H
jn1kOOJel+G9JZbNmYCF/IA+8sO+MpdN3bjfA0nDzcOFeIAa/t2yksJvG81orGnB89mQpd65leM3
ScVPOtS4F1tVnl8/D51iX5Yps8ohHuOIWNo/U6ziY9TT/sLJFMMrGryuGwlm1flr6nZgeEAFnY6N
xFSDayM0fefp1wQybBYgIkjYwRz38tUVgnXwXpk0W2nMUBY52Id3T37oF9F5pX8YJLVAnFImwnrf
w/NaNdAvnyzspKbqWZUFwVyxBvKJNklTjL8x6zgm8gUk9OpIymHmtjSvFXmu3Rt/flGVJAbq6Z3x
y+9GgGZiXmNdpfCQh1S1CAbKJ6QrL5k8X2ZTpRzCD4QalHa+L+NwkH1RARFINz+10FugU/W6o56L
ojSN5HPnwM02yiUPmYi+1WroP1ThYGzWGVq+kQ2LYwLeA0q+Pi1X3Eix5JipQfMvdL7OTAdHAlfF
YDw9M1BXiCw8z+cMcKoEIoJimjYmHrndPf260MX4EWIp2Res2WMQUEDG3WA7vHkPa+sz2ksSv7+B
vMckh2QKMTycjZUfmZPU6BE+IE6U/Vx2Du468qARkp8/rmH/pFiBHuupD8adKYronHD+wLz2j0NY
aDPytldXgYRYfudB1JYtHx0erQY2xW8Ry3cWBkRr5uVEr0CQf+43j1nULMbSlE9CDa0Yi0Huf5Xt
uJtHHy8XaLfJTBfrfus/psnrvC6ojG4fI12HvWgU/XUEreMOAl/+/jikhPlqkT/kFncgMA3aMfwt
mC9GhkxDMh1/18hBH8mH0f58IFhg1ngRl+oqiuTn6cP36PMY3yYnefF4rvUFJdhAoQIQOy43f2TP
kNdIzbsTmGSmKc5DRq2q3jI3BmMy76u+ES2HBvoEu36tRMX6shjU0Dvh+LXSzst7QM3+v/8SkWDc
Dz4ekIOUBlnxkEg3DQoJL02QnCAIZYaJApjGXt5xo4DT4wS5kp7sHddcMi0a25mBN6AFqLdmSF57
CdvyzORJPIhe3MP45F6RA9/REaGOvR2yvT8zkNAIyGWwx22DyCBbdhT9AZMNe2kp/+KbJJFkJEVq
xR4JN0FACjU1o7x3piUfyfYoHkGFyGo2IzCDLHJGd27Te2nHothJVKS1HKal0Qf2P5rlcJVc5F2p
xL0WJlPN7Mm707u5KmywlySGeFK7VknTywT8UGU/1Touc2ua7F8gbHMSvn59C0U7EagGW6/iXKq6
IVQ+H3BcqTm6BtnFPJn4hhieKEA2Spo4LNeers+DjFw177RSKcDljaV7demzIiGSkn5EgYoF9I2y
3eMv4pUxzWkCceeV6HoMkJbFYoIcFeSIw3pApM3fJEOaszVsMHRVu+1E5GX8gQUOVjqomr/YoaSC
gOZL9AJ74BGIol4muzDS//6PjvwEhpDwsIk6qpEFoVv3oo/03iNd8UdjkSwURZIUKFhtWEvGkW7Q
/p+k1K7Y2XvVJLrdSqYe26l90NxB6KVDi79DkCKDrkmjD8b2chMxE9/t0mTgI6Vfb8N45QE4jhRO
axOztZzzI5WNXFWa9sDTMWB+5tDV2cNYcYJfV0Iicue4pk5FLKqQZ9qc+dDNdxDaRb6LGIFTx35T
6FRmCsvgn02gXU7HTnQ/D1f/cRDT4LdrTRvBsZq234tgTOJSu7y/+3xrjI42mUC+yRpiEm7kF28w
pPgZRNw90hI8aCZsKoRsOjXE0ga4pd2H0gzmmoofEgwxLogRFwVFo+do07xU0n03ASn3h6Y8WwpD
UH5jDAVmnbiJNzvGNCIFZSR5u/F1anXsTcXFxYboSYhGMYCWOfZXSliHpC/PvZqvvfLVJ2FehYIi
Z6HQdC6wXodGpD+XLQBD03ncPOa6ZVuKpXmQJFReXx9yke8ZfQFrBeVg1wy+/Ancy8xUlJ7wusrN
EzLdDTJtnmbnXZND6G0m+danszel35jYGPAtcd6mRv9x4VwW0k02MGPnVENlpQNLZaFKg/tAhdaq
pJYuUTq+c6jbjT2ko9oTN4jsB6+1OcFJls/tsobtTg3V4x9UmbKAbRtaZrEme/VHx60ql0ByfbUQ
yfnF4aIXRFEHlhWjYdYUs2S9QOaOzgUu7l2bZH3FRabLCtN+VNLneOco+pDlUSvWqSPlw0TgUKxY
4/sSVKC4O9DiBmEt8gUu0MiADwRiTdSNBLPFlTKRsX3ZaYqcuddVxdJPqdbzn/l9Gaezz6C+ApHS
zyDSekwxSQ0KHgnTf+pernM2KiEEdQhKZW4rTy9p6OjCKQL/4OQpVWTsw7XvfVivjdBrSQkchIP+
xBzfWawmOBQ+Z1iLw2SBpLEFC2ic3LrtYBbM8/WXjd+obr9GgwhpcizRI8+eg8NjEYlIDIMaKfhk
iiMnowjpEvgplQwXx1CXAUAFS/sPFGis37jVK37oEqjAiB74wM0l/FzwhliZH8aQL8bVUDIQVHtn
jciN7PQnuNKpvmwvyKiLDUX1JrmyYjPwva/CdHksye3aZS9Iyuwp2lOAaTXM0vQF1HyxChbAT8KD
E1ezRVCCQg8U24ieRESkXe6uKNQcNeC6wPYt2mKeLhgfbEmysdMVkAZvi8u469FtAmgHgyes+wGO
3pntE63Gma0OKhDEvp58uSn0zldk7Dd/Hfgi//ZeQC2AwpM1nsdO5WvF3riS+4wT/CXOjsF1qjB/
8O7qQEdpejiWZtvYhe2QnKP8DsxcXSmYfWKTbKnHP+Wr7lAkvRwT3GJGIAkWqmWOMsVq38v4dUqk
RA5v2I+0fiZZSbnWkFuz9KRdkdEp5ijCEVetPBN+MOfWuWka42O6gkdKiqcxgqKrFljlI9UNIMjQ
78/LehznFWnfB3PrkndMSFV8URw/FM/KaRZ8srpBcuHcUQ0CpIhVGxg26y/M++Ijn3zFzWVzc1j2
HMYhfFmmhE41Q45yFa0fkEJFhu5MG8GVqxXkmhnwuz/98dONXfqV3qlQZgDVfrIpBxVuXhk4nuSe
bMhAK3TpZ7YjP7HvMrz/FPaqeGOaPWKiKFCaTtxGZRrYvslmRnNq7LOt9bHWJKM33RaVQe0ej6yg
+nNZ9ZMcU+2wsXy5BfNkJk7S8zUtD/0D56jN9bMgWFiDhqEizDicFgIIgnl6oCQDWOwD9BCYABrd
7fhdzrGTeHoDMZZrQeQ+bEPaDCydOvAlEe6YNuYWPBWxB3LJh6Ylm5bZbwmDti95D7It9/zwll7x
nb/3qOrQHzNvJeL+HeAmzGDDawOikWTZwkERwhKPPz4pWgDlb8cbW41lA18kVkhOz4u0Nt1V8sCN
bF7fzAWS4OjfwjmCu6FB9pvMS2TkHUZMMkJOSjyas5gjw19KvBKhdpPK7xk+R8N51k5Qx/NqniZU
+xDWgk8XrTYlGSG3wOsfVgZUsbmQgEA+GcNm6L7d20/DqEyLPfJIGm1An+Y7VbswTxaGi0rXja8p
oN9nTUMRLFvSF9QPaXPr1ZYJfv31krU9v+Wx36oupqc3Ypclx0x3oFX1jz6eboKulU+mFgM0DWL5
0Ky92+1903koIHvg6a6S4oePmA4HndDABRou3viG2+ZzkFXU0S6U86xwbdhGhv+kcQwFf7Fe3/7h
mFeln3zDjeFlCDDPP7plVhkiW79FUU31TM9UAxEn31kL9CQd1+acmP8A03FvyI37QAo5gxJh0W3v
17DfMHL3ZfCiBmJOgpfT7f6o1o5Kml9ElemKUQc4qMX0CEf/DtjHg3T13k8zZ9JJFY52Z9ps/MVU
azUxDawEkvahRKXb6/VALkxa+xmofzLQATA6/M9LRqPRZ4/dWZjTCMEawkmqkRVa8feyHMRUBOwk
9Axe+JW7cEBbHe+m6gcI5/pfong2zqSu1B69b0KbVhR7S5phr4GMMHzra9jJwYTW0otu0aV51pJa
JH81q8N56ZtJFo1t3uLvuyMNxtuDNBmdbqJ6kFLg49Kfd6dn47b0DNXA+3lnv1NX8Ei0f7qhDZAJ
G6c5T0BVynEIrM1OWSJeVRUfuYYTgy4/eM2B1kcOEF96fA00/HOcqep/qSOvAg5hFB8ZeAPzYmEA
q22IuIrEMx26sIGg848H+kRRVNLt7Zs7HPQenB4iVqcpLI7jctcYcckIHdcKGR3SEgOvj1D8BbOv
rgjfOAtTJ9WTy4ZaHmwcjVfFhDVZ7KpwYxZaMC7zx6NPwjNcXAyXj/FMMahoOiBKTTLe/zqcaDy+
LCgKBzaBHvC70tZj5Ms7I/KiJnBcr2JOyLnsWDgMnb7N0rc2yQEH8SYG6iiJF/OpTgzrk9koy8lv
MGnX5KPMnIT4p9SEbWQjI1ZXwhSMHyEPIcptvLAD/Os93eA63HHODG3KmVdtmbcye0AC+S1zosug
9DO1hTNtgaHyFcm2JAq8xR1Iewp2jleDv+4apK6lQt8+IQeF3810vMtbdd7JA7TJCi1yaVZIbkFi
OMkHyVOQiNKZHjnqL1RhMuILEFFEmNHVc5qfXNZjyt5upAHajU/d4uFvuvyPGVgWdWPx0aRA0mxT
TdIw0bv1qE+AZu7Xq6RxYywltF0XmdCBDxf6DC2a9O69kjtNu5H0VqE/S9DxFLGpyOAevgyeDNxW
rLPCERAp8o24j0RMeSnbCIuiiESDQpAgrALqdRA8v44MRNNdOnVeJopxAy2SnumHThLBoZKDLRmY
1CvOOK2Kg/6SM1gJvvev3YFIF+D5YlRQQzGjIbkm6hwpnsVHe+OQRSJNQZxSnJtTbboDqMOLDgE2
FicXE6nQ5P7p56Ohm2ORCvLVKRy6boCc1mhLrxm+HgeV83viSP4wIKKsy5+AdgSynGzhDCvbc+lW
9DbBnAczlYTa1igfexBuYZ7WMkcFLBodAQJEddyHRa5p8sTEPAXok4hz2VIklxxl0VnXryCZw8kU
hRgbHJIaKkH0r7w7YNHy40q4vs0XE1UHJRaHRWTAU2ZMPAixo9WDvWeuVpFIPFhXzFqIy+7sWJUP
/oRG5n3i8626gG9+lddZtM6+nfctZbYzvlJ8emXbMgZmaGK2ePhkocOmGCnumnEO/HOX8uxewDan
3lT6mUVDU9JujISBN+FyTLLQf38UQXm4/21eygDJkD+qT2/8pq/JMY19J/gxbSErYDTtdR5vak/v
gNba1/e8L91wKRTCA3+cAJR9qxAzfiW4F+qaZVDt/QT2IGekeZ2WOUmAXLs/stfhZtCs7hlSScND
ep02ksTNhv325RUpfRlu11LEnYsPPl5Ilzy1VvDTpzopybMd4PDWcc43lZX6kSB9MSIj0Oh/AkTD
ho2rKhnyIolHMMtEbmo/1/FK1AwsGJjS07yp+KJIig0Y/1NqVJUCDTCnpJ0rN+E9D0zr6gMZHw3W
BotveJDDbf/+LE4pHAPNz46uHyNVAKXdSAMhCPsVO9xFnrTuq4Kt5vNDjTdEwaPDeBUwtgNI7W90
cFDkp4Lj84NqT4ljTY7VWZrXGVAizBNevGX32TDR6hCfuLbIbYDFKtcdtGBXat6sfKtZSwQjPwXH
X5MoliklzSElcCI0jD3Vkwi0ZKTR03R6HYK7jOdc16T4su8D8LXTtbvE/W4LfWcvolMDjJCplwsf
l0DUEHxsM5fiD4QX9w8qlikW7TKX8atjrZ2geInxDx/Fhxp7qkGHEhkxSBDFhZ+4V5uIAcXffASw
EqQNVAZbK/Yk2DX6s/k8uD8qUbCNy7ZxGsBaSg5vROAhzECF91GrvJoac137FiiqWART+o/MtnA8
SLRkqURGMFFpfoR8i2hlj6fJaywbkRuTinfXRZCPpq7Po3bZS1GHsDlqFHQXIPUdGXaXMa9O2T7Z
2oB0d3N9137iRkJ5Jx1MSbufTOF5IIgLQpEMHCBCr7IzQ2JZ8OBsCxfNln7msMzWsBb3H9tTaAmi
22bHPp9DziJzmOkeQluETynL8n6ARH8sfS/HIU3f+BBrAKutBdm0we+XTQdQUkUwLfgINqtYUPR6
/gvnddG24CJfbv19ikKavja/RdE4LekpNbcuhXMgzy9UjWWolvXL5umIE5/zsOiI6S/ie6tbAET/
WEsWqI8sIfnNRMdBjrmMzgi0ogrdUMzGB9GjY7xqBwu241aVh4pJ/q3T/sukowBTPY0QXNytPncN
NtwyYCTyUL8DgtYwZPMp8h1ZLi69PfmkztlZTRxQb0YerNBtmrH9E7ebisCc/kqnNUhOD6HtXYYS
AfxDWIVksHDoaF4ZEiGX74AJnGuAkikH8Y0U7iQw0xNx1S7D5J9VyH/LcnrbSg3F2kQwYo/A1jYZ
IIdAlyrSCOpOr8Oe3KMgSZBKzFrLlX3Go+liS57FYI2w20cw8YTqICb9FJBx2vAurpD5Y+Y7TKSi
zyDVLlBikSfN5D3RJt61DXri90TXsRcFU37QIKb5c5BIlxDGQIhN0Q71Qel9UqTYzEWVhNvrT89D
oNELkDR1VdQ8y/QnM9kZrlDuXV+fhAO2FGQyVeGbptOC2COq/Goctq4ZP45CGLgK0WaguT5dkv5X
dUhhwIRbOjZ9Zti5kqo68JSzqY/BJ5JTePxc1H2GUJ7+HXTFHkveBhDVpZmc1vgSqzO+8PsY5zS5
NlBvf2D3IdJah360sItCYhyUQbdw1sWrlXWXPjfVl8q6ZxpW8EovGBlIqX9UmC82FUe3PLYsd7PC
7b5iy9kV16UshWr8m/sihQbPvRXrspZX2L2Ja5NtmDhFifxvYDcolWO7tFlSmwADkfWFwtjxYpaI
5hjVy2SxBgePTjd8ghd47qj3CYfxcRMOn53M81CR6Wrih8QoKBMkwpUJqSrC+nqW/jZ52tUHBvzD
opPQXreOHFySL2dZkGsBkjkfp9/yl0BdzmTo/HygkJyIX21GbCUd3GLY2OANpGARHkM2/ou5Ue9q
+ly/HbWeKzMfgseJ3+Ak4RGyvhwWkXUiGuc0b33FjrF4Tu4i8WSyIvmMkrCJYNGpV5ocHQgjo3Q7
9kZmxj/7WW4rO1vAY9Zq0aIXAxJWIYK7vj782XN8uHAKrw5KumCMzuiUkPXuIzXP06+gU7Z3d853
KCjxOkuM7Y6ZwE8g53bw/lQeGGHoIdjC5pY6E+w1HVLY0XrqVyolphnKuQIxYKdiZ8vJFnJZP9Up
LV2/Wj062WZtDkooQwVaBcHGYQSJt69U5cdMUXJh6qNoO/h/QfkqxSkuyjYcTxZkyUwzSxm9P8ZT
GMEyx9J+JEftxkbAYz0wm3VA7qtB3G1iFSAapf+FDpAzXgn2QPPMo+BA+qFmtipPj/Go9E5eL00r
xymA3uRngyUfVGgy5cMd8Kjx3ivqlUabdbcfbodTotis1IZl80tVai+2sS6ielW+vOIgcKsiZ+ei
bzrCzfXf4EHJDFpV3LW+hOq5UMct4V1krah4/1RhXaJ5CW+S/mcrmfNLwSPeZzOzWyysYJnoTRFR
guKYM12DZIGJv/iWl4Li/HGtA+cq4tki16nnheL1KQMmmqqnIb8Tk6KHW3i4qhQxnvubIgT5EOBA
ct07qC8PDr0Vqj2LG8zaguKa7wWcwqy5geRmZBph0WF41sORnYyW+QFWRR43+hKvETCXnBORtMeP
DAnc9Sc+cNdaUVywEoUUsaP0bjhbGrKqMO+NjbCdawRKpyOjJAPz4reV2wma4W/B7FtFoo2tG2f6
VqebpnFGc4ZDIiGeFVsRRP4lJ7XXdGIoacBO+NFkW7qgbFx+oIMfsHbE7AURT4ZUM3ho/rqqJIok
CMnYOO0wJ7+gWBayE8czsnk/vG1yMrpwVLkTpndCfGP0apGWO09OUv/ctfCYTduQfg60ugbvmWWj
qyf2qMF6EniT2pqYyOrtERk+9q9YrGu8iATbVUdeFhVNJN22D0oOazSKfS3Q7SzQ65Nv7/w/nZbI
kV9WPPoj71ofFOhNPT0IuVr1QNlWKVEAxWl0a/VSo7B86r/6kXkmQtmDAf9Ob5Y14PUYJLsevY64
X/9I7j0NUkd8SKHLX8ITB+EJgN2f+BOkXIBvBoKGjrA07vMNHD4UOV6Yr6R4dY3ZmaA2FJhh5rbt
/bXvPCwLbDxqtUiyOrTthgjuUd6hL6Nkn0snKOZ+0TC9LY26tH7qa95XOveSV48FGdqEHRzcF4SB
u6JDi+xgQlWJAHSb3mZms+ZDNDSbyiGr+gCZPYdHy0E0cTnVWUe8sZIKJvgmduPXwb33lMKkV+0e
WCE7DuP2R9S36ss1qyMNzCf3k4Li6QIxmW8V/aO7A/BGC3nfIsy/3yCenCOpwn2rjwfxaocO6Qir
OfkkYBwNWcZpC+Ny8AhGLEWoObaClt8Vwu96F6c6eNbIZWQduGI5ouPBB/EK2FpQXI2BvXipo/iQ
CLqp4svD2avHypNBOtrUdVye03sjSJgO/seqvIaJs5kTj0a4h1dkx5yht3sis3yt0UeV1lc2l82w
tonvR4KBob96CG6LspXyR0kw/VVnjEhZWHepeBKk05HFZNfXM4mwVG3Cagus2s1+ycIFUttN97My
9oHtK1nMyeFDcP6LRcoYN6aB3xXgqRhkjmN30ppN+LGYrFZ8yuYW1bqFDU00qWU5OFGsMtH/t7vH
O3cgPSDdCiPHUBlJCRP9+P6xPIKOtelB3Sh7DACpuYJLTiFHYKA6OXJpYLFdJ1bgGp8O/PVp9kpe
1yBrjo8/wrX34e/4ozGVxvKhfw3Hs7Az0KFCvSN9xh5Qt/FlcQEFKwxZtt4sZ5YdwDcLMtwLlX7p
Kx83WqY23Rr7cAkChXHeyYhzX9vPFLUpPqZN9Q1aSeWS7kKQV9msJLr04fh6SZNiorC2Ju/21ZN8
i4hvC0gFKtcIQcLudL774voA43wiNVmOzhz9LDMFQbq47DkarSZJjmdeqKdSBtgR+Bkp4RTEqIIT
94PX01AiKN7e+tUeCcC9+uiwFsQEOSxYV+/MVLIEMZ+kfLzh7JMbxxdXB+lTe/b3yN6+vdhevxj+
bxZSmxMbFBaVvwmBP46n1/VXNwg2UjxKhfdWBHzT+5bspHRJu7hhH1U6pGPMdpk0fs+tX0zwa/M+
sNgPkhJuzPlYqlujtXXrEiyqU3JpWUvCGpd7PFv5eq+SshfJAyTBCJnVSmf/BU4BBpg+CNH8tbRz
LcIUW9bwcgmsUlpQCiQmAc34byEQc4Tr1YK1PFv9yc7QgldhKTVCOKhjVL1hPCP1fSbhVSaQ+TMK
Os5JBcXYJZ7pjFa7JEn+gMs9cxEoo4gNYGC4hdeMUQLLwAjOa3S72XRlDa2MUGDPuetSyiiEjmjA
IZ0Rvjf1c009L9HMXOCx7BqKWmLDVlyyR/eBoK6Y8fygJN2Zs+5Tbh4fTe3Gg9PnVR7lHWtC3sWm
/fwhrvDFsVbQ/KIw7G8HVyurwcKJwc+Zsp8DD+CyVeCF1QhbYS4wMiYoihoP7nAliw6CMgaA2bg/
u1F2LTkNE8BMZyIDCLmqvDkXs7cL+CdUfM6G+xjSmdPTWnmg5NkKTK6X3WAkM6UbbH64VMkPafZL
1AmUgdHMhg9tHNkVskFqn6GkboPRinQiisXlxOl1zHHwl4YmLO7kU1jrippX+FEFP8VBcf6ZWs2X
DH/ORWIC90RD6AWpFAQd+lzyMVw9m7AWbUMW8eL++hYK8nLZSwXF3/p6H8Knbh5AaPQhwM/VKyy5
gjHiDqe3cttTGPuCeINDxYyYNQPlElX3Jn5m+A8KbpooWLP019TIKOfvcvfE/SfgRGAmm3oE0IeK
FPWHSvsRsyiQuv35obeD4CMgGrq7LjxzmYuV2C4Tx5lGr8R4BuptLB+5fnVpf5raNlFHFfsD8o5f
cJCYH3bpnt4R072+e63krhGqHXvqmhRFRb0oI51V+m6TRfH/fK6M6o4JwUG8/AeLn3ULronFBf2D
5Ks1dfvvogzK2lL9hopA+eZtvzNhVZRbwBO/ZZ96tlaOSSohhRY4vq/tk8j9ZV/L8RkgXdW4YUdK
Ro7beP83umEZ3zBFMxrYd1qvUXAmhGjCeyVa6g7/Zlje1v593u8/Vc0+T6r40cRsjNi9r1sGq/BK
q3n5AJolhn7sj0Jd62MjxaN+BnN3vjeOipNWnjtDd8rp/BpdWQT08lmVsbolVyfZH+qC4qR9Evlc
6UqbSN3kbV2aEXWuZ/7+zCdiJC/Arw+Ys1AashINCeW73/7DPQk/58v2zXDLKmKSDq29TeoCY+uh
2yJNs8JdjB5tDOGSE7naBoTuQtzH4uSQ2B2u0TO+lkfZ9X06Yzp/ska7bQZFkPFjmSpOZ5JeLwlB
EDXvTAx0dBnnCO8dDz1Ak08FAQvAi5W8BzwGNT/iP/COCIYwKKVvqn9c97AdHEX/Mz5XN86AYm6d
nWeaBveS2zeFIcp4JYoPhse9s7dG37rKtF1LEbISUFrY9LzU2CT4LCCGcVUNi4JAI+Y8DLxsgtKg
jyZP0xwvVTsNCJ5e4DAp8hHrL18bd34Y17U5Hhn0ZJr4yFLONo1c2hi0HxHr+WNM4pRhsmRxK7H4
0zRm7AjXqxf0v7zeQ44ppbZaNdUinOFpXUIOGPmAxkWL4cWV5/zsp1OJrJ01Hgr6G1StGZGiMXj0
YxO+ElM8WmvGLszcXjTFq5ICp7mFMGvNf8Gmvjl2ljy8PMcnKZGcJvJZzpEcj0oikirOY1nxGsyO
jbaUkK07USLwa+EheNEi6YznRC/2lwS+492ABjAU1S+JxYZeK84IMb3zKXRe1fhn+IAEGr64QYFH
41Y2YjFvJxHX+FpmIIzISz+nhJuDlrrC8hAa/laoSfwvJhEOu9cgqzB3FaDlIi5IzmrcRr9bybgf
UA/nHvdIvNSxbVe+su1e4pbsECQKLbhzJFMZPG1utECIM5WVW2Ql1zKN3/MA3cCeaju4kZf67XwU
kJeuIc+F92U/9p6jWFjO+Gx/pNUuVNKgBQmzWWDg+i/Xs4sM0Bci0XGtdZLofH4MjnTDbZz2BHuk
Z9kQd+a+7tvSot3lcFdbkBZ2WMlTOeyqInHpWAsod4UGVTD90y0pRfZjX9ukp7ZFIxxgyHbol4HK
AtsqxcmKNYh4E0xNdAITcZBxpVl2Kob1RU330ZFe4hPzk4QKynS2syq+gUnFG+XA0Zyk9KbsFACn
1WGV2WFIuAxNgvTsP4aK94sb9vY7qHmfBU4ZfLDbb3EtnFlVuK+brvi7Tbq7/uxw3XB0HuZ/7Ogb
AVAy66sKihg2TIMkeG0sUDmuI/U2Hf2R8xxquVKCRKTs0sNze25NE3nxI7U1/+0Ea9PLJxldV6vj
t8wwuWnsM7SeYALw9Af/kujkUAOJRBvb5esB5MpjpzyJgM/orqp/RNavYp4GNCVeh7J+paDs8K7a
6z220hFWSSEg1sst+6VHXHFWhaOpmjaof7gdkYtxPLR0TJyixGFUiTPEoHA9gobnuSW72f4RDBoc
EYZ92/5zeia4miPYPlOWOaQWpEACYTKmuiYkvHmCixP+NRrusGlCCsYj1EE8AQX6EIhwl//+YDCW
nxiH0WkG6x+boaMID88uDVGLndc+1d4meEajsFIlyPJkTk/kWEi5qyZvogZ6YMAt4eGPdkkVxYQQ
49prZo6g08NyCgxjFaX1mkOv5KPnMaFntMX6Au33njIQuYYuv9+lxTsYDUdGoXzJBy6gsqkVfxie
p1sP2niJuYbTsAsBLDQEUZ6H6QtZNJ2U/R9t7/yPCxkDDj5eUgVT8O7tHE4z/NmsZl1Y91CeCYen
HU/+UWVmHAZMTmFpnG+gpMr4usOhD3AHeKEScwdDTfT0Y2dGIks9vOrp8Jm9fsWKDT9bMVmFmlQ4
VVuCZKI3Yf6W213alsezkezdBvvYPMKE88Q5DzwRZlMXVKXd9COnBBJoyxOqkI8D34hb4U/wwS6E
DGdROzasnrKWIp0ZLU62la1MTC/Wnj5ChpX0kl45WRa+Cs7IeXSlgppp/UXj15AU60ayYBpUsl1O
w34j1i7QNQ0jgo+ng4OIB8GEPe1YqdgtvBMviREiAXlDJsIgWA3wmecYb1WsCHrFz755jIcZTcNx
wH2WS7P1eT0zEpWkkGfM26a96GWn++qka70lZ39hYqq28JvxJDBD2RhGKmn1zjWcjb1dAGoSQmnb
9B8/PkUoaRNbEIyz/+nkjSJyKH57BfKsPK0XII3Z/w/PKKDfSleSQ18ux4XS6RLJBraALHaBZqgd
JM57umGAfp14IbQ/i/4oE2WzNqFQJbDu5zzcS1e+6qwqWMrU6GhjNhCbW6Vh7hy6XKUcmqbqYhsW
A6TfIiATud2kr4pZwoM9A7yzdowZ89eTbyJ/KMFxWnhrI/swY6xM9WX8f5ecvfEAZIdXgMwfCUFB
0xboexekHIVt4vkK4DVZseB8drVmOBtZWfmxN+r6TLJLdNgu3Gp5lLMD9cJCflPRXG9ns9mm7IO+
LtxRphs2Bi0UGjFmb+tc5Dsc/j2TwW+KbXyiZLpeUcETQ605iRq/xNyKdq2uC4WmV0Wx0qjSEa2c
sRxTLI0Ta+yw/TkC4FvSh6WSenSTu2VWwZbaI1sBcfc13YsHX7KJ9xeTwLXFlT4BprMBg9IdmngD
K9pBJhRbWHkjurr9WapyjRe4kGPgtgNyRtO79onQZJNiAB48RLAGhNfLMASRFeZDQ4CzgVg6ieIv
mOdK8JHiJKnE9CtVagm5kcp9ZqaHfBUHQRt1DwwFeoRRuICMbKiKcST7yo/mhmDyVJkFXZE2yLnv
oyRsDOsaYHwvXYFji7+xYKedEVRDeHp6AxB5GatRtL1VhAtd4UhsTKC6GksMkqZcohZTULkOlqs3
UqM3rQL0MdxRONcVFfAn6AZKzbcEfPrOr4Cu1O1ocTIcVWYSXebFU3RujcSxioeRrW/Ylw9O6CK6
ez4LzfWdb/VAseUlGjL9Bz9btzhmzhfHd6Dkv2cvv42eU0Q64cyc/8JXZ+tgEDW2ppgHzYSupnKz
UKigQ5rrvUQNwb4b3eSUJFyb/JfFb68KBo7Q8SaSGfxlmWaLjrffSqA+yX5txHPHjhDyemXzn60G
knE7wGUcm0RpXEC/zRnG+f2Qld2VnxL8pbWRiRXRg1IRe5p8tVNVCKM9eqXdPxhXzyK4qDbMDslc
TT3AJqmffBXDvV72yUEuW4p8KrCdnAgN5HuFobYqaDTAwZK3zrYd9e8kk9WYYR6V5m9UGttVE+PV
f0n96r0PjAOkhK2BcDjAuBCpoYpnjnf9wJ00U/1PV/Icc5d2zP/Md3sZ6R+pWqWfJym9DCOtFPMd
RQCz8bvdiqjW8jz6HoQDKxML2+Ea5VEqR92D+no4oCpezImWcY90nk1No/4+ufMkvd8l5CEXan0X
ssPxVve/g4sHLBBuQDOYucaqhW3PfRBF8iPoUg4Hf8wpFbdlkfvbRr7ESF8E/aSO4eTTpyOmRMZc
piTwGCLPBGIBFKU8XH69LEV6R8jmagqx/Ad00QQ5oWjf9nAFGm3/15OHkwZ5j3zYd0w5ZNcBb7Yy
RkQu6qmjumieCpNImd4gmSQ6lCUUI+Yq2JNsxbflXYPlzXByqObzNvNYGtVcDc3x6s5qCF+COhs1
SU/QqqjKud5tbMD+KgS+jeH+yUoDWJcyJkRYyzyVKXYx4uQt1FnTzoVuE8vXwDCrdLtv3r2W5dFs
Z9gmIAB531uMFHi+fJOdauPgr0xdHq2S8OfU7yIKyR/uHNo4hUheyKdLhqQl6s/P958hMapO6Qyj
ua2t7nw5ZlSvOGI6bnmMS3GeMBnOPqR1nLCDNC/ecbKOQotL2SL8AOkIfPba9HjrjfAaIoo/VrHj
PxQPbjxllPXoCPsT1jPUm8twnrYYMSEWEi0OCFXfh0Yzi1+p8CwqLCe87O3NpsmuHuu3rLuN+7Ab
l0I6EIb3KuGugWSiaUWQz1GPAGP5ismRniAXlTz+X+xznz/Lmv2mISCK/5NhvhDSHfFM/v3vSfw4
kPPw2/z+G0zrYWmU9c5MtKJ+ByfRwMJ79lA/UVy6yR690kdheEtWcNcOova24rGC2dv3DBsYm0Wy
RQgFI3+UOabJuzWGA+D/D8qso4FR1i9XatBc/p4V8FqWQrp0ZbvP29/wdPNk0N32MS4TIeqvrKfW
zFk65VCog25Y//UIeBQXlogOy7AflPLIBJLG1NUzJt4LHrobiPloYFieIAgTrh3vBBtYi9fjRzIK
Ho6MkyYSPrZijP2rqH6LSU7sKRHW7ooUmYmsBUYqoPLBslSA0lyn38wSUm6/FbpAv9gG1WAnkwLS
ISWqvfkZLm8A8HcTwzEekdU3iv+fCSdyZPcMXJK2c9hztD4lDwt3udIucAdWof72a5ymk7JiqDTq
z6g/rQ9JshGnv1HaIq0a026L/vksw7WsZ07lyPkxTCmJTE9wHSOyV19xPTt1nGUZwwSLbFN2AKb4
ocNtcpJipH/fPCNu4g9QMzqqOkOWvkZFvWXuT7yi7Qs9RmO+F+abomKbwt8ovICOUOiE15mkhtvA
MeoZSh3bjvokopG/y9ZC2HicH2ZWW28DnCyCrJjCUgt4G+Dy+VYsVxnkJTYxoFHy2nutX147yTC8
1JbrKY02aSIGhWss3te/uRUNWDY4DLQltDzpv7U1W2KmVnjZCZe7UIr4YMd9kpeD+ZiO9DajYJF2
xxYD1hiam7QQ5ow1hANPkok8ZTpXYZJPcYHRlLBQX8HQ5Wl628bxrXpVQ1iaW6OjFuRIqLN7ALEL
5p4pwHv473/c0GoOxNP2Nmhkuny4T0BQ92lR9CyaFtWc5/6lnBHA1/6AxOtJ2unhNdrCmopuQP36
GkXrKy9k4Z4EQBxnpALibhGf92VmJ/bPddy6zUG+OmnCLDTDtKruJySHVl3MhCbHnuOVjY4jB81g
VYieBr+GbhsSXWnSgZ+6cbpIFc1lqa/WBqjwz8fjLgmaVg1fuvzVb5wFIjCtbWLlhJuV7fksIs6w
FOz+jFOxR6nynObL7+qEXGJlAAbO09ITMBPNR2UcxYiSqplB9lwnQKFzytckT2DFgEr/LETHhjAD
T/8CFfjuWW+e8RLdp/olLZDO7nfWTODYoKeGLz5loEKZfmKJ9B7LGmxrEL5WsgsHu8VKzyb1HbN/
/a4I6YHhimd+43LTIGlJaVZR3TZ5dSxheah5UHD2cDP7jjLfNmsKdKJFmzk6+/x5rH2EMinY/ZqG
yXMVq6gbllb9f/6GEHT3B7aIA7lkdxK+eNGW2i+9DYxgvQnKjAXY4gbDwQ634/1zMEDpbmJ1vHrC
LALcgEZBo6de79gqVfQ1rh0C0uNrFj8JGtCk1RXWEfJjtIAkjrUuRp6Mh6jtSuDNTjHQhAPL0gPm
SJhAH6ZHbCYvGmge23ZQjEfV3zH/msGpaM/TCeZpwRmhHTbGNZqBjmfz99KlhGX74Rx5vHEzK0aV
dzHz6Onpt6QzDLs6hzLNoKdd5QLyIM9zDNBhppsT2OARDz1Skxqy62UfuJF3Uph4GSa9Qb1hmb/0
90SuQ1FWRQhJHxuqr3LiIpKCzfIpotfeqNhIQjHII0sBpOjpcWXCSLHcVkuLO6Hq5P1KUmW1QC2D
0TNHY5/SxG2T+MclTMFsr95YAdtlD0bHWdHVhLgGD/2xlxFIS6GpWRYA5L2KBZr0p/Tln6MsyeWC
Cncbp33ObSqx8tO9/mXS+qCC0KXKFgo7i26e3akq+pddEPMHEND7iQ0vjLu4et1Uyk3kBF8y2zO6
9nc5/69ifvJKNKYjkmewViLw2jImJNxdTxjWBeIvTlXuEeITpH4cu0bNImg4rwzMrRP1Mp2mivwu
cmC1Bmx5cGLULLX9ZXsdMim9cqDIiv4WNJG+SikukEpGgEZyCxPrEWf8D5P/FQU4NQoOKlIzDt2h
cUrFPScqI/63ylgkY1qxnroW1RDDytgV1NVTK6KUV75IMnnR9hg7l6DNL9w66sLHfTJZEXh+MsSm
WV8RDFomnfwS07sC9NsZYQHUvSNMMQk3MCzFIDsaArUsrsolKOmE0s9KEWAxcX4a3FFfn3j1nQj0
VJoK0R6/SU19gw4yomsbFnh53dpc587DPskBbRpgPXy4ghRpYFaBAUqNQTKjA+ulqVbezG9z/EIZ
5bmdeMSkas7/Nt6j2+1Fs/HSFSr6qCTekiuVRqNOaAo+AUZel7GGlmqd+4fts4X6FTpHBpy5SSxL
QS1Hrc/lb9nQAbQWaUfUgfNxC2EnCJumH49DZeaBLnON1Rq68+fRBV/ikZc+snUp+SN5PnABnJn+
VSoOPeCakH8JAGDwVj4J4Ye2wSqyGyf0L/8vxjxZANBzpFwH1brit/kCyMUl2UYIQmfqAdD9zw1m
5L1O1k1+a+UbCmbBCw3RS2ZQdEcHe7fXhIf7GUBYGPLfyFc2SagZHUNNyCm8QgeBHYn5mKeZq6ol
0hq/v4kz0+AmbKIcRS0zLkT0F7hI/nvBGOhrq/hTwFBvU1Gk5bI38BschtBkgI5XDaML0fkQ544S
BUDZcTdrauE5N8E4lk/RClm6lBrYlvZpAJGAzAyqvzgN2+UFzqU5kUYIribNZXIRvGv03TLJIuLD
fahjDI1L2VgrREhduEYuCi5gyBGKTg5VMnt2uNmdQGoJ3HOhUlItHXGGn13X5Q0Y6w/LZ2+0CA+F
uxtnu+0v5PeBUm8jx3qPvMyr8pdlw0MjpoVI06Zu8GE5hTVjhQt1dDXzaiV7FWujnKla2aaRq+Iy
j0xKvdgLXHhPqwqWKLHuf06i57m0df8R6UGSXwElckWyFZrXOE8bEGU6+ycUPLmeqP8yvj1o+z7a
sGMPfXr47NVpVSYfysi28pnvdC04E1YgnhA4fNehoTiyLhH23fn7n4XL3sEfn6HKhfUhOas3CfSa
IC8IGKDv+HWPwaFQZOvSas7jA+DLiMUPegEfMlzUMAsY90Fn8iKF/oihoH1ud+5Dc4Ylm8Dr7jkB
8QWQE4cMeFyTuMpD7M6hYdbn2V2BaAJy0q/cSaN+9InKztNF3202Jue9qsQ3kov8pNFJTC0iDcJq
QDYdGLJk0TLPI/e/HhvkzsPzi/moLVDniNWYbWgc7nH7byLg8bT+3ZIVsdJTuUgstSjJgIjZzxGx
BCFtCpOpjXjbEbSd/yqpyGnsZKAXKsbcad25tyr0yk8O3PdjuVtrfzn/P6XgtCF0tR5CXOtGPFEj
zJDzHwoKalAgmH5Z/bUl1fhA+FvlkZbDks1Q5qsSByvrBiOsKZ11MTwZsxI3E8c92uPWxy4N7gsD
JGya2q1l7u9LuJrCoR00g4/n95oHMkbUPkKdXPsoxCOPOmmQ1We0MrCuedbfFIZpk63X94g3VAXk
z00oFDu7PaEDUT+valjK98VZJyU7/uXyuJdygPJ8Kk3ir1hu92+tGHE7sGGzl8o77glQ6g2KfxAl
aTg8Pv559gpgEzjBK9GA92nF+/eH4WFhn1FUHnt9HxDcI4yLpuKTy3gLR8CXzjHRMb/SLIuSZDmW
88jpi+kdQTW5p0SsesSOL2pgpVh8DjbTyAqF3maZ3decu/glre6qOwBhpwNF3nhmbN61IeVrZsF+
MAsaDvhEchNTb475VF7eHuSKLZnw+b/W9T9+puDc8R2RwWsoZp/jHSSCF8Rk7tM2jEpfqpl1Jkx4
WDaU3HTUOG34Sr4q7mcPLMQ3nwggaRb84CmJLR83d3mPDZ73dEQKf9X2tf2VD8rGW6hsE1FcD+sd
u7ws5PtX8+dcG5PMn+4Bnkeu5gtHaz3AbS+EUkxCfAt45IbcJeTqmCwqe2NilInrwbKiXML2fOXU
gHgP6dHuGa+VsPewxqCsD8bhG56NGGfuvmh3lIW2jjI8HaVuZ8WlI7eKQdiPMumQ2qGjcJiRhaId
wWQQ8Ru7Qvs2Ofa0/ew62W1BVn//hqtI/IFwCFQcRUDzJjqlU8upgCukIOnvdbxpF26Nciuwv+xE
yt2WAMc9oq3rB8T9MJP7QEJketYHsAdg+JGhaQL9EmYUtWOg97ic19xsaUv/d56ufo/ECzhqmOof
AOlYnN631ZR7etXHtqTjI3mSwlpF6e4H8Acgj4pFOlzhDKxohq3bLyg3iS9AvTW0IAGAT4R6ROLF
xZMutv+9OC6cX2tXWJQ446dE76yOd6dgCGQnzMp6b+Vvcx2k9NbZE5AVHQqetthZycOPWF+wY05i
KtcTREk0ZZDZ2VjlnDIJpdD7R59jn6k95tLU0aXrPmgm+dU/rZUIY3B4EIuTjcrK7X0B4sDILJNM
0qzJ4TbYvVR7HIC63ASnHOSE839LH7PTUxwoop66X2INRvT+67daR200+O8ZkOu0fLkntg6UJUX9
6BqtyS8uRGJQCSrqqDxEx16y9sKMkdN/bDAvbGdB8j99b8pEsW1ecAhWQkc+HkGll3quMihOi0e8
f8boWom4psQVQ9GVKkqIa9rhZZF8U/3z1kyS/UbCMQNHACnfZNJgbBSoGGcj5PfHUVaju8V0dxrd
UeWwmZ5pLshdezlwiG9DB++++E6p8d3jigT7AQsIAV0HqOPEd6mbgsV3huySg5Vbys0htXfLYtIf
wo7AEFG+vLzl/6EttoJcQ4R//Izu+wCUjL1AGq6o29ygOW4dwD21upPUFM40tFe9t4AnWDdEDA/F
uNoF19LDOhH8TqVf4Gn4YGM3nYzvgHUs1I8+eG6svRR+XlIHvyCFEJp1Il4InBR9CLFWSNUQd96l
qnpXFE/vVEIcUHLMrJk6iMkt5h7SjwM5EohSc8qLTFWpNqCXvjHr2auzibE+ExSXxorKbd6di0n+
88oPeGnrZtx7N6yWqCwowdi+FRAtjvxdEFGkBm1Y7RvLLo6TwMndaPXMNAIBIXbka62j4Sx7Y1hk
Frs6WmBUkIkkh29FVf5z5BUkg4sfrli8BUYmANjHM7BfZNoB0CkTxymCve9Nz6175bMtDWDgfErC
1XrC9ChY28evHKeIPRIQoJFMbubhTqwKlVDVIkVG+RzFuc8qDhXkTOb7oSKcDohSE1jyx7omrtv0
wXSaeCosKMP8YTgzcCaQIh7GeVNo8PwJrqgcVpq1t6EUOX0A8fce7skySVrpDhyisM6N8tilZf0w
CmMOwGkRYyo3yxml8I2JZzzqlsKgRMbbXTojTLz42FtWmNNX9O7TqzHhP63kY2U7fmcN9WHb6CzE
AFaLgEK6nETyoaJXhJio/F/nLQE46GnHy8fgFx2ouJd/AtTUXEHUeAbSAzXqNLITA24oDZZu5pX0
ONQiHKLvmWrF7/YE3PJqRynRf38NCQtHdQF0u/0bxlE+84pOpksicSLfOJH7OsUOxDqiJAlWy4Cu
+KzudtrY7rIvoo4aIHmqrfopBLwYGxL3zgXK430hDgcj7sUkT5tlTxDCWHVQME2pRboJDSUI9rcq
K4RggmmUwG8PThpc+7qmz9r/VG/nHhX5+P3SFZCin/HrUUxyhQnjXbG/EgfEOsMyqL/FztxfyaFY
yyGjemlJBnUp6vR/OqVxNR96bj2bbz8l+pFiX4lr/wACPS16rPEm+OHJx5qTE+rpXxc+UkUQ22Co
QrkkbbG3gMIUcGPwYessN9exRqZNJ2ddr3qWFcZexqp6+GF9xqXCkCj94SAamPRQDYlRmVIL3dK/
DJ8eiOMgmmyHD1WwQmP2YJZfjavsR2zlu54yDJIes8UEmgEKzzObGn/1XBmiI49zZEScK1q3Jwuq
qzmF+HM/cjMVatPm7lq9Wdmr2cTuy77j3QEq5FVNAAveQnW+FH6rqG0pginwi9exUI9w8vALumsB
I948N/6chqFXfqeZ+7YlCd3E3lRPYOeZwewLFniXpHPE2oLA5/mbWxH8o5aV5xRJi4/0uN3bKME7
7aHQa6iJEE/QYCHxv9bBXdmO7IGC49jVbadqJ8ALmBFP6Qf90nWzQ21dSHaZeVaaOml9ivZTjh99
khRVoJf4XKF+acnEZ0cDgm7lSAsmzpZqGMiDtECia0ybjEz1VXLbe8Mag7HFv6PD7pim468hrUav
ya83XIsm3FxT+OEo9ToPe2hRYDYKG6qdFlmB9DzRVLCVkTSenPEWZYjCVF0y2RsO4GQlfZajd8JV
8HCZuzJ/006SUMDg/pvCNuuPdk4ECA+YsIm4NzS9jwei1oqADnvJfCpFY/tVtyTP14kfJeoFa4j1
rIbFf7ItNTmSPdecsIisBNvNwU/7weIO/SE0iduCYjuGtVlV48BF2AoK5Cj0ksyZZvTXNlj/LVhr
MJCXKtaKOXKnNQ8+YD0r8yh6OQ1bf7c1C3SnFqSceYSdDBSuEa7s1EaPE/snu2pJRAM0EoYEGoWb
xdGDVDOmEqXxx/a+MW2m43c/YM1/9BguaK2mwnkTmGK28+2BaxJYdOXrIMoN0TPV/NIblTd8Cs0N
nR8QdW9Oa7/HQIoxJNCVhPft2cXm2VIFWnbFnMrOREM9Y3ZpJCNQovrzDepxiEgmfDLKW2AW9Bqc
oW0lkN2tb+VzUwil6c+Tqt574RhbwaB9WW9okoiQZtElTK8xodaFNy58ZSQONc6bKf6wCgSS7OnD
EUGKyfnfNOSuEkkVT938ExaiTLbDV8kGLrffh2iRwwGg3V1js1LPfXdOw/2m5Yuk5U9YuSoaLm0p
zf4kWTK1JqXFpjjRV0Cq91+tguQP2X44SVtYi6m9ATVauizLryX5lYL3rfcnjWMWq848N9m8w1w6
GAwGl6Yf5zqbDR1Rm3WTpDViuVHfJhSz6jArHEYINEdq1jfbbhIXhd1zzmFOwzbdHrCpSJTyxWUQ
HxVx7xU3I+DdkfxT/bhRGmBrCPDRMBRXdimbz39q5yBzkH/w5vr69Cjl6D0SvOB47J/xpFiSLYJK
msMzu933lsZ4FTG9d9xbu1yXGjzNQVfQPu6oEYhctlRPT8hcXFOwjueYXCeGx690gb41s2MZVlik
KW0m8cHBcQ0fj6yNBZfFUDqHsHvwvHq5Bp/tBaQA/HnjBAOYuRt37UJj8gxtLP9WMq6B2EV4SWHE
OJHDw2wcSqZKEYc0CAmB+xee90+udSu5auOdrUaul+N6vKTAz+/QjqVHhVAiKf6F+Tgf9VxaA4/A
oai0mktev24LY57Sz55bVE2DAwGFThDamo1GAyxNXo7gXNNoEXNevm4JmvteLSm7zPBeI1f9NXwE
uAFvjTfFGPaBillWWP696P3H/1iJLDHMzeHquKSgoumzWkqJJbVHQnzjJCCC0dUvf+WbRVjLsnw+
DqS7uYhuzocLj9vmnyFgOzvPll/H1ZKihZCdYIa2HcpSYZsBZ/nZ+09XZm/s0aUNe/DNnV+gFZH9
x/Ba9xpEKq1dB0Cb2sK9RD44XrZEDN2HfY+InZA6RquMPHdFWmXo6zzFK8HcD6YhGayPaSM8hSCf
9Fs9qyePM1fxruUkA2nCMFIsL8d71IkU6+4yQcKTOAvApAhXvjh0WA2QI0nHInDXMPIJG3reDdOl
P9gWmnCL9r+yLjpk6doBUReA+E1g06KT3xchh1+DYoAqP1ZiYmTl8rfFD0QGrBqY1FJPSaHu/POE
23GoXaPr/nucZr2Oyg2XZ4x4m812M/k7K+mLV/m0r84XF876QgDmFaqORTR+jc46wcR0Nfqxrcwf
k3J3W618ARVqayfK3oosruDsjA+6L0kFJ04TSF1iK2JIH6Zxckg2QxlxsirAGzbZt80JRUJjoykI
tpjPONT2gXYtg3H4A6B8WF8gtweMwaeUcM/IHF8gOMkJGDRD7zEstvN8KDN6HCFsSurR5WADsBlk
pjCEpC8BZpuYDW3swIXUbVl0/Un2nF2Jl0RXtnAFr0KHHNrrGFPDxEkIZT+7jS4d7YGekscYj2ws
7UZlPwsdDgZ3TxXAV9BKedZOBWTuMcEdCufPWAKIKoR5vXzrvyMiYtNoeAOCY5Wvy33tpNve2ErD
tbgzzM34oS5HJNf1ouu4yekW2d0z+d9BxeU99DjlnHDOx6CmK/OWTSPf/0ifENX5S5EsCwaqc0cg
pZ6uIOsDvlxpZT7PRHaLyFW8NUhu4Bw5Q7rTQAHcC5vSUiKqBGwLZ4uCP2Pl1Q9S+NXfkroG7dhk
yFsuGuXs707u2FFoPc4mH+5SnnRe+qv8Y7WQFh/vjY4DgK3Jjw29uJy9y+/PYeMGmNut9ZhwdIae
Gfmjb0QsLv6KRMKVxAQaanK6rq5FBLO14SNGTb7lxgy29nsHWR7UFZOdUIstO7qDOPM8pQyRhaQ4
tWhOFOKbq5DHizA+nRdhun2ATEIFwHy4LXGRyT4NFlq8Dw6GUKLl0KJi9e4O6mCy82TRgqYBlcxg
wqgCyO7+imvqgMNn8U+nlkBdsyUaU0obOJ3b5Exz4yPiKxi43GrKok7Mi/pG6Y5q+Xp7Mv1eI+du
GnywyscsKbAB+tph/2SfeIa4DYjn1O6rBrZ8pae4u47vECNJlvWfsipLfze32DlgFsHQlqAEEymT
Est6P36STR5TnamUIbagNeq+6Ih/peqfGFcuzj+HE0ojY4ZQJmoiKv4RVpTqR4zAZGoFZMZeU75G
SN5oUOcoS+xKM9MjsLohYAXvQMcSx2LCve23jgrPCjnT23u5nU/Gd4MKbhm60LnavoNxZuXJw/CD
jzJHh1QWOUzBsX7dHC4lqHPVCT8Exe8uOPafqBD9vbvI3lSpr9bgdb61SHxRYHlZAgOBv7KfXopx
hRgRLPQnNtW7eqRPZEbbJZKfBiNbz76+3B1phXo/4VtqGwG7BLubgwsoyiCMtbnQMgckmNyCCt32
J4+zXxuVvpsG7TwWB8yl3QHqzrAF6cPhMVVIUiPnJ8HJ/EiPmpOw4d/8Teu/T3zUIAiroCRmDboR
gXs5hmVwFSxdPAk2tlUUy+CfoihNXC81JPqV/d6p8KmSJ+ZQnqxWDo5EfCZ43LfnS+kDUm1gENmz
RvjKwPZTuYBJMoq0Ye0sBEqCZV7MmLsofvcliLnhBCC/IQjdFtGMyIXQCua+cVhZuqZgAVZem87e
K1frJlDe1mtqPgreFsVhzXRVdMy6YsaXJeiYPhfXcOgAVqLqFQW4L+ySTKbgt0sCATZd4vFz5udM
1XmwmpbzSMG0jfr3w4beKHVYE83+82R0k0t0zfDWEhalI/oM0PPZdBvGquNN2+TqZpcX5zcuR7uj
AoaYrtgZryMbuxd2BsYGzkIO/FRsQj5sLRzO+8cAAcbnudKaU5Sd0azTdFODGhEIL8U7rO1DNlVy
DJ6ZZEgNkm99/JhK7wZ+oghumqmtCbdrdVusuUwLN+diBPr6I2P80qvY8uqfcCh0FWtn8pShtS+d
okbgf11pkXOLJsGcejVu6pw0+KrpIGu4gKXu9ncdGjKWqRYCRDI5a+KinM90Dxlu/3FRlFy56U6z
covEWPH7pK03bA3RrYEDfBDLLDqepBZa+nZKU2dOQ7ddqI0cvmsAlolenOlqhwWi5Y6xr3Z4BwJG
S/05LjJJuqmzwvuI+1MLif4CGKM4/audA/OcvQO8E+ZnCYTJm0eZz/YgkXZhD/EGMg/wxcqubR40
Smt5rskY4+JT8YdBY4ngLOiEfEH+Wl4ynaTLemwr0AAjQEn/nxNAN2OLrlqdg7uzvkiXZ4X7poIB
AGuqN4TxpMgqyPGjdYLcS++LuOWouT2bfSqvotO3VDb39S932gBMfYR+sI1xndHC5RWJHrx8/FNX
0RjiyMhK7UKps0ZaTu1LTIGu/fVq3I/5OzeHlEaCbFjwsn1IEP+XozcMs6TKGe8qYXRO8+BvtEe2
Riwlo6CWKsuOHVfu7lJ95gHz2GHvurNozq9QwsKAW9zCPuUN0BMKl9fyav+D3bItBzivnPSefe0n
QNHo9lYLSEUIHwOP9mvgu/pzg0FCGzoU3FLDmAKZYpZgF2D9ypCyuQ/3x1bJiG+AMg9p5iOvAQhc
UAK1wofrIaE/YVPFvCcWjK19lbWMuGk3dbrqEz48jEWpHVubyfIjNVM6x0kEDfGVpKG+i/KEJJQd
oGzDRTMpombsfzQPEOvb1UkBUx7fq9qmKx2GkVQeJNlfiRU5TZOw5CsOeCv3sTczHdJ+g3Ycv5fU
bCdr3N3KdyiwR30DbDV4ctE8Mg58qu44mIwmGfqZKFALzox+rpJRkBAd+Xop2rtA/aRQG403/qV/
ZTUG6+K4YVpMopD2m3sFCpDY2ElsVLBzhKvKZ1DrdWzZFX/P3TiOFvFzWkluNxWbADJoYiLp1W1W
58LPzS7HNwdncZHIIYDMQRp4FyruBxJb2bEJng6dpM1Jsv/aHcze/opNVW+Wy/U1sdcMN2HfZG1o
WGTMGiG/o4au/HwEtCZ3U/taIGGzYvvY9N3TxsmUMUDMz+gAfq0eAsSsNpSQJkHfc6VY9enzTFCe
URXFUaFEPnvhLDI3hMqCBLjz5kNVZMKq03lz/KIz6v/WuCqsHCb9YcLv8y7uNrR2olFq6whVVa+X
gcqq1FvA+8bKJQPSE0404TAg/HDIY/eDq9ziOJlhwcfQYHGjrYAxSf+nyvWzTqlJthkHdKzkTCZA
qOS2j28dtALPRsfaij9U36/Lz6HXTLbHHfz+PSFcqrj5F8AoPZ2PkuY6cDqLptE6vH23s6xzTV8+
yqjclmAyS6fcw9OZXwEexmnM84I2du2TSbBecQgwAudzSWB+5fObkyPanoKMyF7iPJGjLTbrNET6
BR7yQsc15R7XMaXD4WS07WXqiHx5PXZiGVOPYJN6pMfrxzc8asHIP+B0DcSdZEA6ZB93VfhgaD7t
U4huFEljHBhEGJFjN/tDhyAwV4nS/BfPxCcWwlR3E5qmVryL4maAbmN+jCdmPWp1Crcu3Su7YJ/C
/IN5wjYmT60yC0dce5/VxgZ00oliRXzhDllxTnECkVLmN29muEREgX6nRigV7vP+7XKHN9EWO3MH
05xT8LOd5LLGpN2p7vuYuwyXIqBokitByclbcNLvdJKJrGI/fquqHRSrUUlBBIHe61DPnJcFvraz
UGM+7w3L6QJggBtxcXC8AThsHcR21Y06Knp3kh+BDau3H6JNBLc2nLeLbLmZzqE7WSuDmqXTbUsc
naoCfxHZ68fLitEmnZhKvCBKwlCbgqr0E5NiCmPa/SXqXUwic+fN1jB1GCkKupqR9DIUttxjoTgY
Dv4hipgSFdU0ZgCRLTp9IO9swrpM4JWO3ryMIb//Rf2ZPX2/Nu4ROLtaojptnur4qMvnNebOEJIL
YG33KjcyLUAlXB8xSrKELOqUZY5dxm3ZknHraBHAZZcutUzqOoqsmNgyOc2hb95h+KXJF8EosjLa
ywM2PdfH1y0VW/6Id753y7ysICKhpRcX4lVyTWp1IRJjT1PKL4Ouwmt2bW8myDQHgjTM6ox8q5Jw
c0+SX2UbQA/kEiyPSp/jXF96O9Ggc2g2kS3p6h/9C6hEDC0tZfqxZUZwq67ZaZU7XNiKR+pSymY4
Clz2+t89bqPqOR3ZVjiPki1hKySpLnhBesWw3fRqs1+7i3SzwzFiYroGnAeqscDDtl3HaHH03pIV
CTWTIJK6xhRbGtN8Fo3He4AuCZkjdhN3ub/iOnLabTjgvtbexpH06x2V5hnZoXymaAFt+AUHkA3p
y3l6P8LQ24hJ45VkkBa+aToSGwUjx+e5biy+3Nq6dGQPW8wuHiSVNHGKtrITlrv8tP6mue6Ugcgr
Uy7nsp7NWR276aQwoH1uHO6ju+cnHP4qK+GoQ/c2TjrOAPH08StrP2YuZise6b0EGKYqAH0Nao/d
dHgbctCL2RE+KBkdklWKsJrprcwi5AaLgPBLsOeoMJRY8tUsbfKiZPTzedJPnoz2qjuc03AeqaqS
NK7SEo1mYWvumiNyhViUL9QdpumxEsFNUyK5PC0oikbK7vdPAg4XM4x6Oxg8m/vfmjQEGgojdda1
MVEF/psy6aJgCMsbUJh0Lj6wPJCPTbmllw6mmhxVDWi21km95WB/uQJ2XNk3oCckuOxVkPoeuKJj
9ixAOrDKz7sPBX/lJba/9fCeh4/9rDfpHpUIX8qQbYer1Hci/pq8A08QNGrhUXu4IeGVlm6q78NM
Y/2ypw7B8VZ193OFsEwpEwrRf7gseZa/ZPDIdWRqYzVIr0hbwX6jSSBz8NpR0AEg9E/DEzZK3Cd1
dELIlZYJiLY5o/2RQKpQFomtjcRmSOwASZLAVQExnItTqzsvHQ0hFZcryB60vYHSD9l14suxRTLC
IHKYOgAPKxW0JjtxAH9XUlxKNUiRp009C5FTsfLeGcDNSsk52FKjwiSpih0agvKg/MOZfZZ+fd7R
ox8i5QD1LpViAi+KAOsf9wdIHp8fkVUewKhKtap13XqoeTkcNzQs2kB6OVgE28V0tl9L3/i/qMjP
/xPNHtmVxZanFy2nvpC9rX7q6fJHlWyCN8d5A+XOgm8kvFgOylRHEyZKpGvihVsV9MQlpuSocvkV
h4yWkmf9X1K/VXkzNkgp++dcBPjHyeupRZZbTNwuG8KNnGwR6JjdpKqL+Gd8+RA8frSNZrI/jcHr
xyWDk3eGU2J5zLrp4jxA18NFzTVOm+Vi9/pD1PVHUa+EZeClE3IshUkjQMANjsAs+3PG4H1ZmT2S
wzEHAyMONU/rzNdjVG8bUTaohe9cuMSTLvagmkvsXWPcncRwHYZns/Tb5gS2lorlJlhOaG3t6e3P
OhSrhks3gr1Ns85zCNc5aTGznPkZt/Z0uzjZrBhqcHhTDI8HV7ieGVVP8tL30ANEmKKzyC2GV8QV
/EfLRLuoFu8cGfhJHFQUsXFAty23ZWI2sR2wMlf5okvIGrsy+kUK9c1eQ8bpiHsGMBSv6bLjglwi
9cHIDc5JIOjnBkjiL//y8lk+YFV0+6+vb2EIZqF3Mz77A7t2zwONXEKYQTb0ZuhzKkcHkQH0MGdE
0SbS+HYWdKxCRALSCWltmTIQLc9hz35M9VAWIVWkIr66pdno/Zjw5HXOaGFnZHKoQYMyS0OVP8UI
8oaSRxdc1TZDlVY8tIZb9872DcU2JGSW3F3DXVLFEI7etCmNXtQuldnFaCVDAWJvysfwWnrDsusn
aQqkTZvN1dkj3zTrvJarRkklN2y0CRyoWtGg4jYF8EHY2SGjFhkfF2uH4QE3HWqiX48jc2BEMWEQ
VNu5+g1XEQjuo2OtZGYedKCIhvKKM+ks2YfeD277sN7yhHJ4AfhUr4CeuL2Levyui2u16iFtzqLL
Tct2KVvaQIn0fpA1PkkjTSaIvnsWT+H/zN0f66C5STYsIDtYHZJo0d1UEVf5QdYgo2YjsgEtt4Qh
wGq0j/gaPMgMrcpe925F2dSdotgy8gfY6SX3JKG7SA+NzyQnM25D5X1C2oRaiZuv38fVSmWeWnLl
YTRMg8e0xIb5hK4hIpfEmkdymbPSIPJm6xZRi9oh+YV/M2aEAXlP+wKdFFU+AgYhPMke7CFMW6a+
bA4Ek4IB43QKMPIzRW571jFpF51xOyhX7ja5xAIJocqTmcG0KZ4tdluaPnK+xR9m3ZdtVjhrnuZi
mNr3OFGvmjekWg4bd91EKB42thZl8amnMOO5AM2jzuKQ9LglqaX/fAbjxgrDhmYRhaoVxePtmOdT
gBcYYzbherng14jwOvm8OhnWGLOtnmtUZwkGivel8jQzJqw5cd+058ZTeVY2Y+Ti7ZTL7xYsy9VD
ZSsGgldZadi8JvhYS3vZphcuVR79zjVbLBjo6moXwHgP3Wvdz7BDrh76mcGnZwNCb5VYEcin0NSk
iv2rsULZmS+ScBKjND1OZfT4SL0ryZwKFwLaD0FUXB7kU5x0JN/fsKVHh+N7+PWMwANK57jVuML2
fDZXE1hDuzchCyioztw1o7Ee/SAQdsDIom0+NzonL4OWC1cQYTshMSI5buPvHVpkt7I32c/0ZHqr
mxshteN/mx712jmWfOC2+6xL30q9GnHXma1PYI9ZIO1Whw4yVlMB83A9KKC4lCWbBZJafrLnjrKe
f35pPPWWNMMARM1Oi4E/93EZBaXfBW1yS7U01b5XDiZGpc5x3yAnakpWkgtvDaQNoViX6c/l/zdV
giQ1zAiAvqx2QPcRCZNq2OSzcKuHoRiSqXekZQwT0IYXkHmhzd5+g9hV5sXuCYcrMfkmu6TkfeAi
P+APVo7XN+QqPJrHdIvDtHrRldgP/WwY0YTuw+cI5fgOzhmf5d0JsUDrUIrAScRyj7UftEXzHIes
Fag5xVdYtoGqQRaL2SJSnLvzwxoo77wUS/Hx3+MSwst5T8RMFOWgaUCrG6Kji2KYiBnh5ZGgN9tT
pIYLWvjwjcVI7zKZGiBrDP1cQMGr5ivS7609trasAuS1anbVaWguBuHemA1Nf1o5xDeRd2NkFvup
SqbcuR94anPiUTlfBscXS3IOBzC5BurM38s0Z/VZmvu0Gl40Wf0Vm2nQmgbw0oVLio4o9XZWfRTm
wvtvTETWF7R+jrCl0Aea2tcQAvIwziIIjZXDXtWxehldscjpjuUWbYqZITCqBYux/uIhbKv5ACzM
e+Gmoid9YA80iy0GJqdyJcWgTwE50GdTcrbTAJTd/70SfJxT0yJPFtpggV1Va0dkIpMCjbTA3heA
jEuH0ZfjDjP+h/P5fHV2m8nnPV2kW5pVDjy1eKgK5B1Pe6Z5WOKpsYDDgppvgNLtgzN0mHvc3hvc
51eW9wmourLwwLR3cFHTVe240b8OoAOHREsNvq8kLJLPv6GvfJBKrhhbGWEz8AFGfBqA9HoPi/uT
rX9MshgEl6rtyoHsPMCKD7AhU23qVie8cWmtNEC2kCTHb3Ik2cwVBJq8KRefI3JRNHenxNmOmfFT
WKX5PoODro20wrfyHxSbUxHCz/s34ovh7BgcfwaoAPO9RiSzl4kH/IXDWOfCuVh70pSB95ZwDRB7
Jm+YojblbBNjq+bmqgBxAmYkCCxcA04qnMrYUyRALcGedOdzSYwkEHw3VdhmFfoxgopqJ6PqqMNf
1jaIOjqPoCVNhgB1ZQha2tx1Yh+JS6ut5r9/m/EEcsFKw/p2t83tN+LzvEs2ch0cn6GMw0GELGlC
inSr/FIPkDkw3DQbzZYOw1UxEyuQRpWepVzPWr8QJsp5cTTpTp1Czn/XixP6O+FxPT1FuJLVRF0r
QPlOxwHXUaMT95MVmoYd/RZpbnxwObzyJG+TjqPtv4ymqCW6mghGQH0R/vvP3740vc05loPTPYJO
lVMtwPr8xPWpNYffjs+gDslqHhG9gp6I3w574XDztiEqTf/zJ6l88uY/jVDZxlvLOSEKZSr5Kp2N
MIHoGAzKN00rtw8wXi7cI1cv14sGcy1pNI9r45ZJH8rPskBYWjGb7JZYTOUc3KB99BrK1YUAlu6m
ZV7D8B4RT0bJjxGVk4qzUVR26GSmPRf20VaNxDW0vUs2Rjk2F+Pi6yY/asVQy2Js2RAR32nxenSy
dapERXkfl21IwR1JtBHMnoCXrqU9eKC1D3FsVjD85OkwbvMiV7dD2YR6QGP7T1ycMKVbKyF+5sua
CNsvWoieRwmcNvWIld0tEf+wU1gxCt2/kJ6AyNcJ4Q21eMkMYVzD8ndOfpNT7WLkJBfkSTcLP+Ne
ZIyLH0XUPCZ+GRFk26cgmkDYpFbFRNT4AaeFOGPnDbogZKbJt76mc/5peW7xIjaBMJ5m/JrewRZF
Xu2Bx68B6t6KAfaSTjOr3QZOzqZPYloRqIMVxPiLXqbjmp2ML2xoFBrN2VV3URCJYMF8cve/X3sh
D4Pdfefqp6LmT4dXe+AhZrOJN7cH1aj19r0vuMi8zUA7NyRsPL10axR34rdzvlJXI/tCHj+bilVP
UvX7+Ct19W/O057jWy9FWk3UWohRLCIPvBmDOy7U5UIg9fuR+pa7fPfr4n6T8CXh9bwbgl1dMSDk
/rThGvvSAAMYrknZQomRGdGNiCNHBdzZyQBqp16XpXwpe3CV2zfF+6Name/jQf8kyziqidTqzfjm
SKaGoC8wtzvYKpGuZO5DDbWE8HBcI2VJOuhvbmpRkWyvBVcuQx9SGzkSMNc67u5W4dUgS3xd1dZc
8aioixfAkCU3fxKwx32bBH3N1/zdJ/6YEVlkKkAcFG8KcLIyQMq1rOC829Sz4hLz/XfJbiNn2ySP
p8iov+Ug9ae2ThS3+/Cpfy+FjyMISW1Rveunxjzq5INFzd8idxTpGRgyHKxgO8ptMawyZu/fyZwm
KYNwRCtTZ3E2GBU4/Svf/Gq/KW0YYcSBYhzEyrKYcPTG2YaeHdbm5tm2HnPS92SBS+u81DWKl++0
DitzAdqLFWUcyrGL5vQXuUNXIMrZ3EbIFxQ+WRvyBi3n01xTUe8TKeH3hkCKbVP6/ok/A9fl0QVl
qAoD2pwb1CllH9BvwOHigSeC4OPJn59Z8BND4qKEBncSFaqb5jSIQGSlaWSxYf8dY+0c5xp5cr0l
ert/RnRYrvm2Y+95ECMZhlxvi0dxJsp3ts0GM8q5n34e87x34yqKJgHiwLKG4dgnxbwOB1M8LpKd
Xq8FTt+6xd1FZNT48BCfrml9w71msCynQ09OR+henQeIQJ5sLnTmb+zkKR8G34TDKu6rBTz3wPfG
Ui4FlPuB1E1wBS7Uk6RC14VFTJ/Nf6U9vBb7GGHUF60GICStACzEoW4S2Vl3GR6Yttq5AUlDlHie
1oxuo+n4h+IH7MvQHmnYWmexbM9CUNsEXQ+AU5y4YxHPIbBVOgCzNwYc0LGlRNsXckQKLeQ2lP9q
w7VtbBYExRY6OMfVpSlmdbLTTDSmFbnpRFSDovaXsgEv/diohuLQUHv6wKG5kHojENsexGyvJvNF
8mDUsKh+CeR25ZFjNBbO6V5L1yh58KO8xKyPsdnODhH6BN1++gt1oYJHg5KUKwpYYklZWJn07OG2
pJ6HmGEna8nbT8KHkFPRN5OVFqyMwnnxPFudmFP7rJi3jM64yuJfRiF67+ziEwx4ID68EvufGS+Q
dDyGLMT8nj1IZAtSTmcKplFrPasVzCK1CLJO4XVr4zQDPpsW2nNFe9N2rRZDX29IWCbsTXXcLdwD
Crxm7Lyrnux6dJYui7AbNMAVDhOEDP7C6sZIyN3ZvnY2laEsxn/KZ5JT2z46kHKvOCoknN7DA7Sc
o8KbsGJnq1tIfuh7uqHzq6h8PMvYx9wLU5whGMFLk0jDWjfCYoAjRg7Qe9KhJrMk9ZVxNMkJ3zsJ
XEzZdJTmTAhy7mby2MlizCawc938xgJ49801+NfaZ9hhS0+dIIOV34jWZiYJ3pucLmwg25vE+koP
USVSP3IO3Unc3YBEvLXS2WcLFkUhfcr8ci1rlHZVuF/FXlOejhNlm+I8iB9gmj8lF2O9NBTSQiUK
HRlFXEUJEv4e28gMPUivw3b8ia9i+cqGTAP/Kykv7xt4y8r75wKEqU80HDt/bJ+LbZS4yedN+pc4
yDGRpxWjMPQMVpkdbnHpaGYn5NddW0+bVL94yCHOGdk92dE9TFD5pX88mptLSd1LpGMrnvedCOzD
JYAOcNqQBGQYqft0dW9Gy2djFCmGMsnXPaI+IFOoA/b3EX4CZOAG7/3wFCMaGTA6qRpqN77kiEJ6
SKtRrzdqgy32E99YObwNXM3aTupdZ4g5zBZQigQR0gUX7nhYBOgsGoH8rjRdpsDs+MSrbA36rqVZ
Jik5GO+Jtccm9LBysBNXS/JRpWab4YYuz+G29O9dQxrkeeP7mZrMK9sCFgDs5+e5pyLVCsH+Nd8k
jQL5lpheywGwu8AIjRm7LVR742ftvNWGyNs9SXMGmQx1c8ddt4Fcj2pGLRsZCN5Zn2UeZvU2iVJP
i/FOh4M9KNQloDCKUYCAxRT2AO8up42g+rXK9k2ji8oT/r8WYV9wfAWPjRGWuqA6omxpALIqIbAo
hGOwnDSgFgxlgwe3k5NKMffkvS0Ev4h6All70MswNp0yOjaZ8wbOT/+2BzKhle0mNquqqE4RPJkK
6ctYKh49i9kx9gSah6+wyxtfZqIBOEVbXAWttpI/VrJkuJDra5/W0p0Q/1vxMWaVqNu59v0Apc74
xtCgIvP1V+ReOp/qaJC5ynuevDyPUyWx+LS9TTJ0CP2/nymvzE/FiL61+ks7W+21lsM0RcrNAd7y
9f53vRYnSf6OR44Ko70fXtbIvwP4liqGaLnIRUyuu/g1Lkn++IJKgAZFoYzE7dKtmnIKA+J2I1q8
vcfqNi0DPAdn9X/kR733fjpIwJ+beq4KXlO60ui7kHIN4PrsQ0T+GeMx0b4yt70yFBdmtpK591MQ
jrTbgtPXnoHoLtVwh4ozZYE5HLbCei36QAPUY/aE5wQQqLMxuukUvFM3rJvRlKR8fb2Re6GJG7vl
dGx8bve6sT5n+JjcVN7Uhh9kWUyYXvRlZ6YVth3u4yxAbBFHXDSrEjsVw5v2O3Ii4MbooYQ7kf52
yRFLDTj0MnbZuGBzHlKHpf6/YcSTM0C/88MA0MSrGBFARTp75sOq2/t2LXnyC8rBrdeX+vZJO728
wuacrlsFd2Dz/2lezpgSK4ol1a0F+J+wWkTVLbWVJJIM5pBOGSc1uZES4bD3xgetx9mO6rf7TKEc
024cEzn0IOX1LyrB8OyD4JZ/e7iui4SYf1X34sPpKcWr5/Z5ZiEe1hGa9hGFbqazjzZnSjhSw0JQ
bzrPFMbG2bL/IXPdFUnyi6cSJJTQGGAC5Lk4QjPPqR2LfMrJI0eztv5RrfoeB0G96mql4nhmlHfQ
O7LL+7Zlv2iPW2ymmH10iKZuVnXed43iMbhM5psYVYyHWw88h4m5qdI2fsSqYamKZFjxYnTPQXTK
G3sS+2lBVT6p9V7LFIEdB8OrKKWyU3aMk+34mSUkLPnBih3mf7T5lAn75j5yGYMxI0xIlG8hmM9C
jdCEnBRPv8wt8jwQpoAC95DImTBGIbPeL0HxCYRWxsqLtCPeeHl2sgCXOI/qR5X9np1Otx5qFRgj
zO3hep1+Anj0d7RdwFc1jU1D+Fy8pM2gGNI1Axh3myPTz4/NmUGhtRrdBRER4GLbL08ZDeKhmlxy
HWi00gNXUGL+r+J7ZvrAASiHCI8A1SNf8lzw5VTRAGZLsMu2Neb1TDcBhiJss6ACYCmoxfVhGFK1
Ef5eI1lGWdol2ZCLG/XDeu1PGDFjvuce4WHpXjrX0Xiz/pxP4aDI7kAewpDUmEBgOHC/l+xZqUle
nls5nLPuCDAYRozHIZ3ANob7Hpu9W9pKUYlhXUanHG1326ut+gRuX3gdLIPZ6KhtQcrZn4NzR/HU
zkn+S15u4B9zdV4MJx6dQ2s/v7dT9k5zo1QIlWkrHYHJH/NYkp42BWjZ9vVp6MeeTBTYuQ80E9lQ
so5G4CBOkRHsa3tMP+vfQC8ZCW24/7Ml+b8Eyo5C4Tpk/0BWbYYh7mjJctL8lWqNYwqwld7nbr4s
DW+FobrOcHZNokIEHLUyPPg6IS0nmPHTmrvrjFCBBS3QRvTVjAAWCZE1hwaOl5XbFBuEoQq6nt9N
q9yQWZRfzEDn3ASHuvX2X7eqwHU2+LSaZ6KbIZ6Bm3RnPxBoqUaUC3S2SPOl3d15/hDQK9fX3NGP
fNtzfCNvjP0wDA535KrP5TaRVAKhH14Gw2jxLW7kF3HUzY82/WuO2900xUoLR3iS1jKisoNusJwD
16m8jto1ooSyXIodg79DfCC64PoEHd1DHDCxPl4pWJR+pPipWvMx/SWQ+YqY4U/6s2iIv2a+8Jpo
t/nX9xfg0gTtCTpu6ff+k41sjzHt++5K3/6Wieg71aJnBAOVci0tKe+Jy93fImPJZ8qQ/kYYKlAv
61VPe3+wjqTzWecvRKBov50HwWLHpoP4SoLnchiHaKzIKbgKugkrOIvC9V1q4qBEuJB+e3sboLml
kxbYXQPNBcz8OSWxSjjkbHHSub7/YahgKjdCR2hCW5baVkQkms+vBlO2UJatsrcPS+9DrKufMmdp
CyBEkI2Cvvhv39flMuprOcqUzx9ryZv1vJx2NyResMrKTX56rArrlOK1YdG6azsDG5x3kOh/t3B+
lb+8hww+EP7MHQkNNPSuKhoEUtKxZQcuwLmfVFfZkU34cBmUQPSaO+kFNp+Qtn3KdWmS6nfNJ7Cm
G3mshpFNwwFROd+sX2n7WQineLHtY2rYSfr/YJ1gUTmM+RJnttsoDfyhTyXVbhwxpmRfGqc8WW31
e/uB7+jTpHWs6nmbUq4WfAB23bs/7UulyYRncDjURLCMlfKteSyv9h1flroPhz+u/T0zA3EJdP/L
oqMi6+GO0t8m6pHe9awgnUDzpCuib+phedOoHnGvKvhl8w3f83FxCa48dPoBfVrZLXWINFWLpaf2
gCs00tLkA3MJo1c2UYgvlKoyEhSIjAYRHEsufoAontOWXkTtfWUrnqLY57DUREaXoIVOtcZyBg90
+ciDBVj/gIHLDHtD9jPDGOhncYv7HKwP1Q5HK6Qx1nfsQi15xkF0oBes4mhYS44NbaDl7H3EMF8P
sCoQeDa2pul3hTv7j2rPYvrpz7lh87Y6fVgk/ePLFIDdYxrymFxIJQLF28UOdoHRUD/YuInHWjD+
J0gy0m0vZhLAaHocVO51+fSBt0xSOfoR0FxsQTwg3fwBI/lWc6cA9DyKSVDrap2mVBhnWwy/oSnA
TIb4dF4kuYFZWoLU42+oXl647uVnliUoN0thW3WWwgSBJNsp3PqJJj4wYrO7sFriHN+M1FqcPZ0j
pLhUty+ZbuHm/KQRiN3u4KUOk4k4X/3WoTPnIy/gVP/NPig+qJvOb7wrzwJMa8RNPr/gtiJPc5G7
KHNtaA7xlZTfxMiKlMuUMeSYmdM5OQzjD+anZnzbYt7N2SA7az8sUrBK0e5F69dcMGvfOJIJRLTg
wSKUDFP8O01FBJ9JwVy//IxUZbHVC++y9d8EGvwYtbOXKLua/ksHqBL656EEXqd1ibkTJfdKEYDP
+05Efbx8LghlN5Y/uA252IDsR5oO/crUcx2TVMOZs+v5LJQJPt0tTAnaIPadD4wSnDgXnK0s5H1m
wCsyQr7TE8evzLheWnGwOM3Mcq0zu4oMcBXc/hiXHdCoDuNYv1Q1wf50QjqrfbCDaudMtcJInB62
r2rs8oDTfAC6b+DL2eQ7dPlj0IQr4GmX5m2gACYURIxnIk8x+ueoNqe5Z/3WOthS76fFx6db/F6G
9hCbgD621rzekfp1n3X85t/wa+PlqTcloMDA5+dpIBsUafcs5Han6IiFYM7O8IwUkp7epql4wfdu
Hldc1pziVXfJ16puy4z5+AkzK2r1qYUy5an8nzyZTV6RsQ8+ixeJBAtBOv9uFzWjCSr6Tx3aREVE
rfvYqYcZ1JJl6XOVnT/03TqXh8Tyqrvr/xHlN0/NnsQXIaCdYxroERukcQwlIG5oS31sBFbjYfa7
h6ZN5fKkRwrhShwicJjJ3LfAWQP+d6lbFIDwgN3LkYNKydUgIuuJYpDp9E8icAPIpv0Sjd1jU4qH
w27PU6I6CHAYBYEuWQyeYCX1nhIEWAe+ukzSiaARYW+bJrbKyoFQce50LY6E3pjsGF0MNMvhMPOH
hdVJbY5hI6/5JP64EiDXJtyDHDIncxnnEtSj+rixUxfm4Gam4/4NRpJ/tPJrZlEzbBMhvvGNA2SF
2zcp+C8TQHiOQ/chF6rP4z2LlLtGaG1BkSyX36l6Gg4Wc86QjfC4Xk1lzlj79hCqArh7keudPawU
BSfTleUdvPgHP9UgIQEhh6nBqwpqqu7aZ1Bt5pVUCTNhjVAMdihDJHPqE0TyKx0eMmNzF1lFhO10
ZsMlaWV2ljsK6ao4vwGIu2V2stFKVoITtI/ao+d14Id1HPBdAM+GDFRykqTizzCgiuAAuWEAjUUJ
Eikot92pGfE0Jijmp5J2FtlKwDymAUiqhwxU8+B46bVY52Q/E8z8HJ/+McbwZ3tePJxuahOlm/Ce
zwsva4+8TNgdybsk4eZhDwoBMl9rcUJA7CeQ4h3bp8cXpS2XdBxDBkAqsRgItTJTBvpA+Ryblequ
pYOgdcgJ1J3g09cSpdEjo0zlm1OmSQsB5hdbBu2cNDpJI47J+UHzaMFoKP4RJIKXx6kyZcjFXPGb
jiRtKSRqYFAi/4bFcbbknf558U9j5o3mcPRA93YRwRWjM5jsZylHMFco1EK6z/ma/ZFtXZ9IWr+n
AruRVAWZ8iWAPuMx4FVwa3evnYqs235L+PgZGPGW53pB6MmRaNRheocU33VbAl1go61q33yW49FB
IrKipnhVFZwjDeJhaAZRRAbrYxLo73O1Sos8ztN0f5gd4dKh6NgYBiq219YKVQZbSd+hMrlD0AiT
4IRVrcvPOXN5aBnVjx00J3Ap+oFFOKyU09SX7jj67BZmjj0NhutoC9G0lBgZssDTd1d6XMKqwOKi
yW75QOWiRe0+PSz60Uvi9UPtNYpU7sA0YAEMHFKakGuk+OObWMaQzWP+YBhdgFmNgWoHjDtL1Vp4
5DpRT/4O8bomMgKgtcNZ/J+iKaO4XeQQ55BPJZc/2bq+HHoFmqu2WYtqVGdxBRaF1dMiGqDG9Na4
OOzkWlHCf/mdaw4AG6gGCAxC//cNLyOfdhuVEM9GwIULFmHgjWRmWAp3267eZRnWAPdrDPQ6JMre
3F69H8wAxwXuav84cHC0BGxPSuK1eQj9jQ6x3G3VKX/ly3DNa8JBjLyVu+Mdc0ySmlpkg4FI0eBq
VGgsqUQ8WESvO/DtUcWdqASkeWGpmQiQH7tJYjEfHLi6NtKjTQwOs/dTBgeiYSITi6OXaETGR1wg
Igmi0h6td7+yUwlHhJ7N9ZYnrWuz6w7npaVIBGpC6BHfmouFY0dVnMSxrbkfPYfcKhaX9xSyeIYd
7DzI+1ZvBNYAfYXUcogAgRLoXeS16t5lr95/KO1oCxTDYERSx3PciaoWWWIP9IWa0sqfFGlbmQH8
b+UMx81Fyr769Bir3o4jBKxtw98gDM3Jm2okTV+nHPS6wnLbGicTDYN7+0D2Pwvej4OSTziiTeME
U/+a/UvKws0b/dGdduqaAvxA0LMnLHCfh8tMw36+ZQ0wA5UbtEklfCUPcGHT3KAhQTVImlO/Qnha
rwwzZo17wu0P10BZzKMSOhtCkmlhHFF3SmQI14jTqM8zB1S3yB5aBs/jSIUGYJty0EQfYGillmCH
9ClyVzXMsM3H+MjtSzaXsRLD8rrgXqwiLai9MpCjSA1IfPYtFtLiQnODp7/r3+7rZk7VL8oZc37m
SAePnJQs8LZLWK+h3scRmVahE3w2njzTsglQyfuWSR4Hoob3/REfFJvZLwhtaxX/NUaA84OuVcQV
onOb8W1eyt9GgrL1fRD5FNUZ8QqLWt0oa4/QGY4/MMX7ijH1egFiUQsJWTSopmZh6rr6JTcatp8r
P92bQkP60ZSE6Bd4kVQXuKyqI3pmWWdVgfRKHAktFgE8azvmQGJD5Y355NXG+eNXwVwlH3V33Ljg
4JGeYvkelXE3gCTy/Y1J3E3FKigG6odhWE2B/xXf0M6Qr2wkkXYNCSjoxbtm9VIbNiMBpxUr94V/
VWgXkNyyrLcnAeMY3iGkhQGqtNAiNuD/hAbfbWJAqHINlL6914r/m7p2B1gBAFDWvJIiVaWi1L2M
TcoY9qavZPQrrh7nCDONIb/SC/7uKvWeZYmfRbL0+ObU0Y9mCVMmGTB/tR0Q2lqqmLkugTTcQkVu
wWq8m/aFPM8TBCMiAs0zqIicqbsgXgETEDX+6vPpYelZdZMSyzntTAGYi1iDniQxj2sOxKqs9Ivv
tO0jZ+zCXLLm47MUpXxGWO424GwULhwnzXcPhuCNOmWMbA5BXw+CRuxczR0disXsGG2xFxwvYvJX
uDtG2/YvHxr+rPCwL3LigklcaOSVuLezAweMKEsbygbsxpih57T+bBR+FC4CQSLMz7BvcFZMx8S4
ECONqxG1FERjMsoU9F1LaNWJeK0e1xLuFLzYuzXGZngzA/NpNMldbx6YMZU1H7Uk0mLX1LfqyEas
5S3Fd2yZWXM0rlfo2Jpc9NIpGYrEIdMmuf/JsWaUvmmZszZpvYqHyaLHo1EumNKUOddchiFsbLnH
zDfoNj8J9lnK5mbkK3/l1ShlbtOmc7+jz7V0i12Im89CTyDZa+K7pbUwDie2fxox7l4ikXadw4FO
tLt00N9ojVQcs8Q6kJhx5zO4tQHq8oiWCHQlpx83RB97GaHPdxi38VGC6n3tYXl1VY4bSGzo7/md
JlMcl2TyyLIo0RoR05Np6czsR7B2mucCqvwIUDuCjt38rwp2Sj+tQypUUqezz+qGyb1zQWoxC3N3
3w8hQxAWQLtLcriWSvA+2oR7o3sJZSghEwJgtLWTQGD9jeeMf7tQxQT0OM0cA/xC1B+FnwtY8Hug
rdyxMMOJyYkmYSy1UxoMe/ALzUJ+HvIURT80UNx6zlgoilTnDM9eBk+UBBKRHh0DyDb5MY1jU+cG
iHggCwjf2vcDUG5wuAfKlLjJBvQS9tnamP+MYiimNrs84dFhia6cahSCSHVHrhWwbbr2jf9Yr30i
GByKeHJDu7fxgieSd5BilMMYBXVeDy2EZiGCuGX5jubwhc/0rZkzZO/Ol2EXAaahAgy+v8zkhoRp
EVqBNckQcxXZTo+qhpHk/voN6AVR7t86Fx2hrvyCVzDzU7rwkRxt3edyYm/T0IRZuCHzqPEWYrCr
MCQFl+ENFabYi8CG/gGsykToc+zZ2fqsqwjZUdq8lrYlUmQA2yf9AsAY4TSmOOAVGLa9cxPyYXDX
h487ZWxVxAv5f6sK0vE/MsuZ+zcYr5Sd3IY6zqdsG+eAKUzI/pD9TkOZFT8nue8gCl5p3ZmMFjof
7LI5Q3dGkOIU0bxOEpDZLNqufiwY6pgN9O22eYZSvXYzY+V+FX703cJHJoplFyllzEUqjOOM2nZA
90iqMJxatwBuXCNRl1Fo+r7WxwEemvnNIje0OHnxSoHeUj6+Ojjl3KQhbxERHLDxEIj/DRE1s6Ef
k74sj4Nmo4rWU41La1awNoHbfJnHrZtepvdUwwy/Jtsk787GMNlW2R5RiRmJwc6GzvMJsRibuP1Q
1ZfaGDNL9VjGmKp+czr2IkagsdHgqh/Mwc/mcGl5j3DPd10IPDSkQ9HlL+128Asu0BxZSeQW2bv8
P7e6fHKc123sVNvn7mU2QWJ5bjuwDBpUhQ4qig3GhiW9GhpKUg4TwFGVcH6p75oGcV85ioEH9ERN
fudX4spqWyKSPk13/uVN4OEWDZRK/u42U7JcxZtL7cYisI8ZtWLxKMsvESiCiUDQW7N/tjsRjsI4
a6mM+RVDcuMTMzPbaoxVyp+PFxcasyw5FcnLBYuIHDb25/pNjrhlCzqik2Q7z7gzRkTN98y3Pd4p
+u5HgGyod5TWWN0e+30SAfrGlNNPqd7Qju6m6LBf6olE570PLDzYqn65KS35eWrZ8HVeQm/PLYjw
FEUCJfGmKFI9wfvcpW5cGvtNBGYy0fevA8wkxwIsfiZpQLW0A3YzYYRfcMNn7MwDkLSvElD5OAv3
9wEYEu1i4yNuex0jPQdbIt0NjVOZNQ5Hl0CTozdZznNEBJjx16eBMn98eszHx+KG5bCYALYZM1TV
zkNFLj5Ovw+qL+BOCqOQvJTfRcYoFP9grp2aOluKgzKqDPmKiM5xW8ugsVctsIAyyNb3+4tgITAv
/JRp7Eo7X2XM8mKLIORzXpqeklG3jmo70yWLgonWwyj8mfRjYbzgqFbwhqaVpnub+l1aMULyDSVd
TA8ALuomd5+dd2pJxta8f3WgIaEfZ1gUmYb9zzyZqYxKWC8s35kpcP4rjmXhsELdCpQpkCFTLWSV
elp0aH9lrL9ENP81XMjrv7FHQ7z0QWgX8pZJOdPv0+qBqtqNrrYVmlcHsiRv977oWpU7pVzqE3VB
NWgBeuJSMtAivPDBn50XjoRpufbRB6vMTu+4+BO/qVVRmTDoc+6XchBNn2Zv7IQf7DDqEBHWo3kh
RwWgA1R4h1o4jUyB70gffw502pK0e/x8GLXJQ/C36a76mvfs7BSeG0AodD6+GvNNf4PG+knh6Hs8
ILn4rLe6e8ilPr81tcmnS231gW/I5cczwjAnCCts6Yfsu1JvcyCpt4P2O+J0COXRGbg34OfWaKZ+
oQSie+58GYedWa8DqMMNAdmAZ+YAgpXic/yJ/esQXZHUntOctOFXf5stZtI0XRm6JzydXzja97EV
WdHhjeBxbJixQR2PGQujTPNiKF8h1uHIhgEiv3ZlgYGmC64/0+PAymXn9MLrvwOP8x1ttelBBbmh
8LyPgFnNCbTFwhmPTq1A5rb/Q/jwoAIMzy1WBPem/z0jZvTrFbqmICtrqnoCKZ+4pWzWRZgF2Ga7
pHXAfAmhSBZ50SqowdVPVDRbScPfNd7/FwX8yuvZnwh3iSTm88rnkB+qHFbIr32EwgeZcqM+xhTy
13kZDusnmuPPaMwmlT6aK5ITTxizOpVsTgERhfXSg/5o6f9lowSTgp9Gqwjlnb/KdOqNRXCQZruZ
CONetdzD6jLS3DrdpAMrZ1BCuC2hpaI2iOr6C5VKIJhmus9uXIgng9NStTKtliEuwgEaNevaV0kW
4EqFBZB47VkSezvwmH6lrJbuWyVE6iE2oDhGbPI0I2FUjrLCOYyTDwUvigYlxlFhFUZ63WOVuKIY
8BTaiC9qEb65vjpk6aOaajwX/cduBfMwxhk71+S80+kkQe4bckbxHlb5az3s1oOjBX98F57ffBBA
6ltDly+TcOSYOvt6nUOjCEOOX/ckDVeIolAcD6BZQTiduQ6LVD1TuC2ryD2a/xzD7ZX+KYmVE7IK
pOebEBQ+1DSU1nw9RRw4LNIImb5P8O7XmzUKdVoh5TlkoBjVU4WuIFqe/L6LrDRMFzQaERswjPfp
MRW2LrW2CZ1p79+MPER/x1C9bqrGs+RqMsDKBHZXo56LAdFJQ4hxjobjiF4wsNnxocrb1iJTvXwh
zbv+6yn1o45ZX3QLs04bZsWoBFGQJr+cRX/WqbfsbvHzsjntHxMSJfUvQHQQSUBMS6Nmr9uYIxKA
6j+2MloQnCtEkh1YKysFMeuQx1i29jyXoNTnNF/gfumPe8nQIp9vO7agbmB3KowEqcn/q+1VDq0b
j2qpEg5SxLFRrjRKpDi1+fU7psC6OGcg7fCRBvicYHK9sn4zSjjBNYfKFgFoz3t25a8MbS01pGw1
Aj03/kgZA582V9t0l1rBUeRdW+aZT4CM5kFe3yPLwd/59xNXCPiBTU0Zy6jIW/jWjqUN+CAbq2Up
0cfhdz7VzqtWgP7G4oXfqKQ5Xg1wyrnv5V5OUZb/E+gfQBse8DjaDd56NVy72sHqYtrfriEpGAKG
VlflLgfySoUfTFKCLO5ZcBXghWsaGURniM/KfYgLi3Nn0qoHA3JNOqMTGJ57xR5JYDBkxrqJH0L+
SRtc9C9AuBUmPKGGCqNvulh+uV1vlQa34P5XYLXJc+yU5ChS+JTrou/upa9OsfH081ZPtf+khpiu
OQGMljXWUYTsI7HMQ98LWWDywxIIcltymYlEMKF4SXEzVDRFczLRL3Ucog6Vol1OzcLOUpcygH0b
fQeWsdXK5+s3j6y8Xi+eWJouY99HoH+PvZ3fco1xTK+udwOolMKa6jd3EFbC1tTKQZSDRFAWet2U
swDwDCyDNFS4B9xRd5UnzigB1WYtRVRESyIfGzJdIuu+mnQdyugeXUZyuC2gDxhAWDZ1rlKLxIwg
peffJ+yeZ/jVhlOPy9+vnBSGGjdIsnTNYG9kZQvDZ1QzulmcgqV9kHJ6AyX173371cDTdjkAUerS
sC/ckGjzDKtorHYJFBDoIYHkbK1nq8xSYTq7u6OVpW7BYvu1rtp5RCdgzLMm1boQCVO8qXLRu85Z
BuqoQ2pg3ZVbg9JSIRadG1J0mjYw4ha/JuZQGRJR+JpwkRqrWFYGJpaZhbGcJ/K/FzLmXjFhlU+h
lXwEieO6jHfLM6NTG6Bt0wQxDEZxpHkUDn4Q1PUXLdlnuln2z823kYMMKWIrn61iSjVLipHtPzWU
vQfSpFfwAfMZ5k3Gfh6auk1x5DgUqJm0CSq08YZysuCxVVsgIMICP43pjobqr/zA8NmN9vJ0oSa6
JD3MqmXVKNTEecfWpmJkz8VCjRnQSVV7Hffuidg0mbPXLIUHoqjbDeQT/PM2dl3HlKa4F4DaCLCE
w8d2vwPp1Zrc2jXD2B/BF6HEp3eipHq60E+W5V3TtmiUSyrCzVLzectANmE3RqQ0keG6F975Mjqk
+oAK5QiKdxjZK4qL0VFIZTOd6hlrg/92hH2y0jHWk/7xmdyGkgJEvQh9ZOAf8wKwfEHkXnmiOCGe
w0FOVTPJfU+GMWtxSh3ZQ1v1ssXrC8zzcFbaNhs5V84VgmTjV5EeNv6Yq5ri/+bjleQIXMhTf3CN
0NSALTQYwGq8ABpk1tppU8PzDnMH9USjYjEOV++YY2h7kMvKC2/f9NX/b9tDSXTx/AMVL54MxEjA
2yshQ/wHbK1Jyd//n7fzztmoYP8qgKP+KlbeiWmfiU/3D8UZFYC04FECzSK+KDfauqlpD3UllYs5
9AxyeKNRzgXS7SABYZdn2AtFxkZXIoCTyvkvird4lhWYMXuursFPg9Xcg3pwheKBrjUhl8Ehuxpg
wdkV2V4A9ZepGgYH8KEQjWQnT4CMiN4kmw8T88P0bnxSd1m0Jd3etgKlFJaBvqrYKwwU+U2nViBj
jsODgxgDsOJf/TbdTDjUHaUCBndKVqJaPIf/DbbMPgANZ4OiRkXuBXAVCaCmDa3BKPYQ3RXYD7Ul
hIU83pQ1IEfgcIemfvReGarBkxDA5qi0gy3jrzZg1ybC0r21nbgX1V+lUZSEIrsgTGTVpXzz2vND
vwGxjmoiMHtNIaivfKBCq4U4b82cXKrnNb17S6Rtyoi9fRI9qrdIzmbz+1QD30beh/9w7eXYOxEl
FBRP9dwEhkxk/Vsk5uPmBpfHwRO5WTzDAFtmJ3xvSQWQJhcCECxGez+CB1Qcajaspe6ZkR8mLx2o
G2WF4CV9KxU8/IjmXVXhlpuJzfn1MyitUzz7D6hybGMQz+FwlHDzO+sIj5kfJsQs+GGzMQAajzvv
bCy7v9tu++jNnBxcHchnujBsLZalC99DGhq+1wj9qMPK3ph4fZ6Opj82V//nn5b/bnT/XIj3BSpr
OqwE4UdoO+GBg7azeaOJs2INqjOqmzz8eAjjaeY2hg73TnTYEcBlqF2LAUfepVafkgvJX0XQhROO
2PxAzkjolyWIMSrcYwLV0fxxo4dxxmq2l3hjnFLo25kY0CEpYyPe3S4MB5hRBQN3YFtVvF4nHgtq
RmP7BchA7qWTsPdJFuKSwy3Cl3i7kXqkLEOcHkuwHd+6+vAhjvYlhRy/Ha1PNvCeCT5NUemjcZad
zWOC8tp0vLemETGhdLdrVbXRVbzAQX9FYlksPu6Nb0XipHWixEOJgHuxKIv0rLT+B98sTLA0MID0
EfGGODkG5Uuj1e9kwogJj3fTzkjorCI2eXWIBQWFvN2KWx24oob1FM9f8NAytx6x8pv+5PADleeT
YO21pkQYyqAXtPjGAcTjjkwyNknNM4CkQPdflL4WSYkM0aTU3n8skz1JE/rXqLNVTABB8R0F1yxz
/DgiuFSfToY4RIR+VzmNA1tjiXfGDOuTAfkBRyH0nKtK+Z27YpTGfIwvJSh+GwI/m8gBAQYwmhGe
8yDymACQlaoc5tODpDPpF0mOEPYnXx6iwE+tcG2JWldCSU+IWaPtkBQZ/tMYbX6brwk06r0g4UkJ
ZAzMOtC0hLsiZAQi/l/cpca0zfkH6DZHWu9UaKN6DO3fxc5mbu/gtNV3BlABbBzGyK4H4Cnv3l5y
/Dl5cfRNK+6OCem04e6lbP7iqlS5LwpGOjB0YenHorK7EXCyy3fWoKlsG3LkEdtrmvF3peyLeHUq
qId2BZNffpw8N3B4nbTwTVKyMJyHurxneypk5tesF0Vwwi7G5lmTsJt5KkG1Cl/rMaekKIXRX/Vl
IVWcx2RXH2SqndGU1byEfUYhPbTx5ItwXIzohXUgmBT329HHgqW/573c9lOXjG2IkkDsclEWFNbQ
88zy5djvl4zkMP+HcaVV643V/pCPAlt/3D7KqY0NCIKjCwHyvObtHoeraEMTE8jWgx8yiivjYCLP
7cKW/FZqi4M10/EXykWsB9HMh0eqPP6P8nJyvAOFP5bJh3a/+E69UGybfFnTMJLwms1rsf3YXP0Q
MhOu+eaL7mrJ6T9hDz8quax+RB/oMLVlth3tQFh/0UP+esNaV4//CLJOUbOvQx2g0eg35nlEUAVk
iARTMCWWBYG/1nTwxXvWgMlrxBTpd0488N9OHc+WtizxInqKqXnxKOcUQFzazyDXogZPRnSgFzOJ
kcQnUMo8yy7z6sg+XU1QW5ihPLiixTs7yXCh8ZKrw/2XT0CwG8e65CmYLU3Eik6dYRIjENh2wcpr
fvFdSi58YyAMrKUDqh0chqOt7eWqIhcgwajQT+QQu30vZjZXcGIsvc8Ti5F2IHc/SM7fgqd76P6d
/4Z2hJcXpLqZunccHBlL02pWcQAhxUaevQIS6ItmY2ER42LzHZ7LAyqqm7is+VxshOW33OLvm0ND
U8v8hSFVBswZQB8UcDROWJ7Q9gsU2N7JmlvZVHU8d9mDM+Iz2u1oOXHm7v9UK7SDHKOVcJx1veOZ
/6Byq1C3Xf+jKLRZWsUiZDDwgzAd4T8c2qjQHBTkGuxaEr80pBkoDyP/fPKOSKdQdDg7DHE5hzTR
vu+DI7M7R5/jZ4+Fh+0+pMXQ3FMeNAp6aKPzYyrSls5mdkVfYVAvglGb5M1znqcH2PZb1dCxGoIq
DePAon+0mMyaOCrxRBrHu8BQtLxVwPmyQM+nFxVi69wFLLyqXQoyszh/Xq0hgEH6GFEJRgPklMHq
L2tKMf+zMJ30J/zaiW9cXVy+UKPqGc/Qi35UUS7ykXyxT8fVHfuaWSRtnEdDKQb6Xw9h8/fKGoBs
ADgPP6riTkFpzvnM1T0k7IniXHUmD/8tXFfXjMB/Cb0ukWTsc7pXM/ARQtpzzJAnggMUxHU7Ejo5
lahqpLM9g9PamVmheDCCeRigdtuLvXLqons0uIqYytq5js33I6hpEH+WziW5T0uDdzAYaoIjViOj
VBq8rOUYwVTf/nDspU8wbxxO9puYmzC49FY7OaSaTRzO4sAV0kmFNcsyfv1bbHGK/KNuiqIxWWMf
Eedw7qr77Hjkt46s5gkMnQ9ixdiukuSiwZe+iXIyqjZDhytnxsZn1AW76Q25sxH4kZ+01ZiBsJbW
Hk72LAeUsabChkjk2X0XbCefJBZxijCj/PNQLTa4WCw5qyjHgpjm9dUHWWwt8vAZOWGxR++YrTYj
czQsVCSydv4i5WIwHJ+6UUtTNz6Dc8WTKsWW+hCktG/1ZBx7BlJp8xXKdA903memNXi2XezkjRp4
wKCZ0QdvrnpS8MKFyf2Rhg/bL2jCsfR0qApohnUSxaVRcsmQULfA403RkFnsVJptNSsGVExJFZxK
/7V1tr+MdscmzYE9eGRFubrh3CoslGDX1M5lVd+4uNo+614UfUrUsojyp3/UFEuw7Ac+0Q2FOXwD
Jyr9cLZLjP7aczKoAz0jGW8dreSW34NWwxiVb53TPszjMeLd0RLVZ3BdOrSbgNfzhIukNu3qENGr
fO2tr+ZiMVzgShCkm1GhdNf0rU80yWBH+/NMmpMPyGDlurivripPu7f/TLt+9Bgi5BL9KemtlwiM
Jq0Xomlv5XMzWP7OTrGpQCFkKxe12KJpl2XdJL7d+e3TsVdq2Q44mtMdVw09hP1/TboyjAcia8bn
Y4OfdFczHHphHIJ0TxzJnfe2nlzlSkxIch05Qsq5hg/HrvQFZdUlg1YRjNFGONFv1j8PRMVgUEWA
zTGrmTPI75NXPmQcxAbPq2eb+mz4VTQq/jgeJwHmmPZ+xtZ9OPY7s36fWQUi6IHGBjq0hKpypKGq
GPUtVtcezywBlfCGBNDdjpmGNJEX5urG8wl2SYtF0lvB4tSZAGf6yH/gECL4NJ5S+7pj1TjtuLRC
NrjcST5fy5xNKDuJMa1olj+ZB+Y+pbXnmawNBRk3wcHYYiWqHW4aIW54bjdXK7FKbjt8C35nQ/PJ
bK9o9Kdf5xbcM01PTnCSKMTT9OmQk1myArgSSISBd0Nc9hTJZjIOoAv8gZZTl4LXPcOtoR/RuZ3T
Thh7aU2/Oz1vybXb6CFIJ9sZRzyno/yYHemVJc/asy5YOAtYXZujXI9FBI45+wF0YfosU+ZZfOgG
xlclK0JdeG++d4NECmDgETi+XNvVyHc5blPAEfIHhC+92ouGjsNJchvND6Ol1t1xXyGjUX/NPq7Y
mhqLpxepmU6zIUq8puDmSxsDnbpgS/BdUQ9h1fZp1y6d4o05bqBkpICxJxjKV7O+qa1BVHpY/6gM
LMtUE3v3T5fpxnBq5umLCsCdhS6FBRs8o3PybGMXg9VNsetnSSaSYFr9VOAGh11ik28/3vQ8jK5Z
FpvIrH5QYUX/Ke//9EHnKwWrPEkYYKZEiSwqjpHNPMN/IGZvLoFrcTQVobaJVk56yjRabg/2uZ0+
kYUhZ7SQwIgpD9+y4zH9D+b/ou4rKnDIsPWjqibFitwOjI2hrhKKPSDP5wn50XWeWWW1Ac78tEOp
8/f/bswJCJ8hxUns6Gq/bRnmIvHwG2FbwJrbt9ZtpbmUYnV6pxRFF4I1rfIbG1TJpE6jfKWH4jqs
657acLGu9c6q+Ls3y1rDUoE8qtsVhxMlxx0CZYkM3vfLz3s0xl5fSixhrQiEn+YWRSPVU8W+3Bts
po0+ckmZZNda0oreD4kEMP7E8IWdqWsXtpHRc3GAOMcFKy3FYRprsEtQe6CBmGejqh/IR9gNGFwy
w9hjO6qzf0XfI5HhOCd2PaFJltHiqDtKDbNy0V7BstX5CKPMnO5SvvFrp55Ek4Y+9nKSSDzrxTWh
0ojPIQU0ELwO7ZtbY8iI9rpq6WQOaaCLWi69EVRYV7YvHI04QgYLH3utZqVs4rbRFOWz8RJrl+Xw
nnuhWwiwJHTnd8Afxy4Z0U/gRvSlrMe9ubImUEOcLRtmSFD6WY/GGKCC8ertISxUskYFRykrdYBI
u7tuR7SqWflPnz7rrmB2BRl0WOA8diSpbPg6c1sTEdiBY8UoSyQqfOkDFlE60sPi/4PTv2XLwunU
wnmPXUIu09fXnrbG+o9ZIf5QVmDZSNmSPndZwprfXxwrfBWHb2ex/iD0pv7ioAGdrnT8wMG67Azm
OYbm1BSS/kLv6a+5gu+oa7evkGtNETkFkoeJ/yLEOM69UzrHRX/BeDxrPu5vouFnn0T4eUSBHwnf
zMqtl7h3QiN67OgCVDc7n5YJlpw5l6Lt/2gn5GHNINYDPj5oqDTqpOYe0dAreNEKm8LW0ELxcmni
j12EK2R09UFWOpmxvFgPBvATHyRKxcE/Wnsn6jTI4J/fpl6TBnbimhDXbXRH1IRdngZ3k5k4WBGI
Nnqd5CSCT4GQPyJTxeUIyOr41gTu6hFQm9T3Z/Tus6RJZ5AE0HWWSLYqgE/Cw5U/cNsafgr8wFV4
0YLM3s9jnCmCXMh4JmH9QWcKKshzsmEi7wPe01h1hX6+HLASjjQhr7L5sE3AEUymBQhOjCRJq6wG
J8cspaJZLphLAAe+/2mbeaQjA7AXtxpUQIdV8eK47XRKTFQsXcIBDPuxqYpOaE1uayK9uG1TOIlF
k/JUiRE9SyEDXQednO8YyVL9s4QF6OXZVlBVCKpaArhnqHTpx04nJ+MI9YS6+EXXkhyIqjcbnYiP
MEyNzC/bH7I8F1TORlY8XSmc2K9TQwTua7PkzVNLDtTyOePR0j46S7Y6zMAorl5DL8+3fVgu0xfv
8pZrZvlFp68h5qlB/IpEvXP0l761b9bZHh+Wr2dxvMYcccSnzmm+9yV+nrpvpMVJ2BETtxIcWTs3
hoonGUo1B5bT/pgDZJB2UguUYjfb8TLfMjVCV8LTpgGjQHitRNz+Y7y7tjPk/QNu6bOX8Hn4t+OU
wUGF9L6tzT5u9gGxVn3HTtyFwskvGvt7PUpT6uNoLeGYVEq2EBEPDk7G7xnOH3drJIixPbs3jvra
F1rl8aPpMrl62UCiGHmhLC70Lof5UNE4XABXrFY6LN69YpI4JhwgGQoAR0zdFy85kLhOGFmJUMDe
/s6QOZgXu1v4mjUltFsR8O1ZZCOK/rVAgDDRyRwwwSOQK5JbS0wdMbNF619jxXxrKmddHaQL6Bfx
qDyFU0vr0rcjtOqJSRG6pHlKvPB/I1eEUFAvWmWzM2fc3h0opRjLvIPpIT09AwuGvMYQTAzgHZXq
rf7ivDq7skFr4tAjqbI3989YyaajWLqUTuMRUWi72s7RvRbD6/yqDPo9++RCAFzXjhtjPrwuK+YL
LpGr8fHjeQ12hFXHVEwSClHgq/Y6bcxNeLwI/PxS27W3U95uOzAF2gyz/HM5ds8N9nBox4T0cV8t
+d4c54B0lrsO30vz3VD0cgO3Iryw9uVhfgG4UrvxBCwd/lSs1+zS2CtQK9GcV4vJyEdWlAyqBfBr
OXdFiU+AQZB9m8TCQkvIfG9Ym6nTsWxZobC/IbPSLO8B9MtuPaa1fYdFj/zJD0CO13GeK5DwAi8y
Zu+XBPWC8wTNyUoNOWX3UqDu4pkJLB8qniTi2IBJmNU9NHxtFrV2DlYQJ9rh5WmkGL+SH0W1L0QL
i1dajXWkaRMz4DQ58+eBsN+a9aGhLCnItEfYEuhy+GAyeODIA+r8VX6wLflSoz7CC76r8nTwlVzn
LaC5X+03wRfgaF0c2H7exp85Ze+x91TrnM1CXI9hrfBPloxdDBlNVxYArJrXFmvEUdghatCwLitS
zJMlGLO6wx6nqBhyGIxoiyU51NvRl/9F3wGHfUygJFkvnDJCPycIVGNfyj1bvHtxsSW/5gYVMDx6
6jNmL7Z7I/07TNfv0FnktUluvaWSye7F0zrcWwyg49qIBiDrNxri2QN4323KBJP3Tlk/6YPrLpOB
v0544LzbjF5LZ5CkHmVJy+lLlD2wRSQYK8lkm0BkWg382u+zo2D15NUjMVRDqUGw/RkXNZqWib3X
hgbR6rqAL0+iu81y/nSlAgFuq9znNHY9BDNZ5fmtMa3phcX4K8ZoUwqlUxgSJQ+B9w37R4MdVCxM
6ngBIaVktfWsS2SNppGJp+M1MFKn0VS7/BmGEqZHmFIlXOZcPv/TgfIBx0GICp3L+pbczrXWzahR
S/Ta1vzzfS21ZEYifVx7jwqfPlF99oQvcplHUe1Ny9SaUfavQrrg2QqDYItpf5j7HMR4RyspUa0x
G6j+LuWWtjKtD83NxFsu20QVm6Xj2fo794D84FEVST7a15hqYGu5LwX4NqghCG9FvFKTOJs6B5eB
rlzwo3JgEyuFRQSYzT3dA5dTze4oiPWKbh6+dmo6yjLHcD7WfqZHoYxMHgx7aFLqdea30fZam2Oq
HalSYFSIQ5rCcj1zs/4bxTJ8oHUUdgy6090RL5tbK6ondUGeEhH2g41hsI+tcB/QwyUQeGCDD1gU
m5q8OoIw5nK6uIqCfknJesMT4x1+mLy2EUVgiS0FTZHWGViM4tVPyr9RJspQBiJalbv/UKjBR3qk
sjpCnijKrfM0soGEZrNeutj8HOl01ocIp/CNfE4pHqHzDDG+hfNOcP51cjbr5TTQxaKSrbBBs1Hv
NkJnRDwJQi79grcmjgin0ZZaWYID1uK+0ZM81XLnywd8h5MJiErWOlqnDU2zNH5CGMHeiaEmuTzf
1nWKRVfe5OkDzN3WLd/qu48WL7RJf2rHYWd9Z2ZfnBYpVWQke7qj53NByk2WnkT2x9dr8VvjwcuP
wXFLd2bKw4G7AXoanTon8w53MjJCI1kMFoEfx/hFAHF3fAlcGLx0kuDUNI3B8oDExMcmhRPFkeA2
hH49sTJAovwWKXeR4FK4hYbE+3DCe9fwuFeUC4bJpwPKkio62Ra0/Fi/ru6zMQx0fnogb3ZDXDRs
OlYdZBUg5vMMGiY/zgNikaZQXiyHvHjx+DZod9pnWZAkCZB6dTXfyJ3/m8KstaFx08Xo/MNoPaGT
E/x+dDyz5ra0HWAs2ArXuWL3Gb1A3BgU7J1YV6j2S5SQjE2umDKjmvMB8xfP0CXGK7zTtBTp/ocd
YT+tttllTwgCjJ8czGC1opiaDJlZVtmYogs0CI/9JB8a+n2os2+DngRuS80pExTwc0hFX/WevsOA
sErLhPqaOyTFj/YmYPkKv9AhDsEDbctglEzuy6DS5U3XEjtlbKqWTstu9Fps6gpC1kGuFc3LAvqd
XKB60OXNOLHAciNp70AqdiSUme9qbK6E7vdMeboV4Ddg3WIT1lHqZelcREUasTP+9Obl/TBAuYkb
bKF/2zS73bl5i8wTyImrVyXF0gKH2lEGWyKLpKdNpL8ATSFHTByy/4rNTS6RaeitnsQlEvA+CeW0
yUu9Rgqh3fWjprk6OnQn2id3U17gKOPt/rcnnadPf9NMNYrGEFun2DjvIFolqXWsW4TqFEmjESb+
X2axO2ymn92exZMo070OtaSIeD7/Ze0uSGhagP3dvsrF94LRJhoQmFLtQdpnZE45CS0VFQqICqVR
W5sM+Ptq1CnZei+GTTfHgA+Uk/COR3NPTUGES63zuHJKli9XCi0pEZG7xYPv/dj1m5fYbonFVY+M
0whdAkCy0JDS6d+A0c9muaXeckraGNZ4EXCJgsCulcRDJrLDUmm5Dno/cIT+L96N8i/n7lbSZDHH
0ZBTVRInwnTBA2OHG7z3lY5hoIgwhQ3Lf0pmo7nq6f3lEfXwSUbXzmnCtyJ8iSI6iqORdSgXqfNk
AHNrkOv55aaIxTp4dv7lauk9Xqe+JlQXAXGAywBDycKvUpHAnCmpJMIePtVw5JHonuhRnYo7tiMZ
8oAJ79S/lcwPsTxvT8lcJucTtxSgWWQqCbLC+YVtipUtslqAvNBWhDvhF/6ijEc6so7Kc2ARCMZk
uZ651cG0k7Ir1gLHQJA5q886AaIPYwnwKFnO5VwTwMFWE51oVODwIpGx+1zfxV7t1ucuji1uXzmS
STWlyty8w3zIG2r39VTDAzKVvY8jT9JybWF8dHbKJ3AseyJ3fvZlNE69BSrB+qDEI5zYibRxGFM/
Wdz7DmzJcnh291mQY6dzLscWXwVSJMHhq19KqYL82E2fgBgfiM2jsZw9nPCEYWVGkyxJbCazPc7n
zSrzajobi5ZcfYPWnchZx/cpfsxiYi5CX1GENiQ4s/eAoKZUNUr8kFW1h2sYSXLt6RIujHWbeuUD
7CPBJtXbz2VLDBtwsLvUPHpoLhmLRKElHQnwRHG3k08emppv0xo0GAyqcEaCtAlHX+3E2I02HSjJ
l8KwG1DtXsPJDIvP2i4ltlxMdHK+UbuAQ+EHzFm71ovLfk1T/H0grkPfQTPvFe6Dw9OlpcENOQQI
vhAnP+Zt4cTCJngyZDLJ7JBidgcy+fsbwocRthXbB12Dv4qA97sqdAI5vHmre5h/zlZAs2G0X12J
GLQJmFIlXuB4SbhrkfCOFM1/ai/l6akXdZpsmtV2F2LZAY/8MkbA97tNryB6glgOQC6eJ56OZdeH
vTgER6YI9T12EPWk4YGyusK1cPgX0fp/K+s+oDl5UJcchxWr/YYcODWhs5NGGE2jpJKQO9Khf0Ya
m3sG5QFgT3QfaNgNG0ByoYOWoyFt/5yrQ3yDA7RmBes9YiaDbvWxdyHs63xmQa/FcOEKeurzpr+v
lmRSAmQiKPR4Cq8GycezWirJ9vfkhQKQzUUfHv89sG9OHIStACO/Ger+8T98XoYLnVJovClU/gae
yCX3R2Tu5uoWRZ/1AIFHWFOSHpnBhzOKL+8+woo9G3oeo/xwEbYMHM+Xh9Rh17kXESkOz39zXdma
68WMVnrKxFONgG52LAZp6BAzyHuDAiDX8bGc3+Lztv2kKPr0dEy1YVuoELt/ePRGmZhEDg0gzIId
EU7JnMLAbqjov+XCD33du8iRnXin+VViLBnS+U/qAXhwOeF8Evb52OdeQBgliFX7FGt/1ncrtp+3
FXB6YNzNFe6cGkQjcX64jqQOt7qydemKOwwHJZeodRuaoPs2qdhE8ZXhF69QeHL4qSG2zVb1ruv4
oRiwqdiQ5KLfZz52KF5R2hdtDV9AaOp7T2Gr+tKfWpgSJsyw0fURpYWen5zx2jOs2TpLoaoXbxwK
HaJTI9cxZNyitc7XJSogUcbgZZs7f72WzjNfaP6kPRMqwFBAWxhbW0prSmQeIfXozh3WZepXt+CB
G9Awlwov15rsGA5SxYSij1UJBMsBYjW+dZMoo32+KEMe1v1lLW4viKtdLQYKqC4wEjaPemRKEy3W
zAK1hPNQduXkgfaMH+5DLxW/p8/w+vfrnzT8tZt4z6cDxRksRX8yMx6Y9KNzugX+5pxZ/JQytnG4
a34aoZOeYAHvER/faSRVfx24aOdHBpjBXadp+EPOIpqghZymwWyEq1/COM8Uq8BKlA7ro6BH7Dy/
3+Jxl5fRMuQJoIPWsBE65Z1v6F2qUE7lKqAZP+jiAUUV736Z6BBAWnk8eJ3KEvKPJy8PUm+cFAtG
c2zCEg2xlkmh19ZncMFNMQqkAKfGIjfyPjzyYINBVMUCqQjF+zT4+eJJS5fOywYgxY9vV0BGzhcW
IKvY+7Ik6RxWmhVK4I7kFXXLlfYjM/TqgPxdrCv93PrfMlqeeMK32YB6U6ctmIGPAlmJc2tIJ4VJ
DwbUs4ey3/zb3Ufws5j4YWNfR7Zgyn4UTfuU0q+ScesyfOxwfeZoVNoSGHmjIKOZEr3XhXOZMXgY
S4ozeIfk94e/2o1M7rmL1f1mvEFgHYB/ePu6DUMHWBJFMy9pzmww/Ph1NiEwtRR5s1MEerbgorcP
5wyAVA6fR3mAt2TZM0TQdNAFU0E5LQPc0gWm4MhrSkMFnQ7Rw7SuZzSrmOdJTFuRFLB5uATww8zM
JbScKK1cD8vwWNbS10ybonAMT879DsbyD0uSR4Vlj3J716e9eu5rEiEQWaqINevQXGlQPw++EJLP
r77/IOJwd3aY3uUaVzTI5bd/OhESt3EzE5olA6lGrRn9O8OC34kZGn4oxdbEVH2VmC9FFgy0HyRx
AFFNA1EnJ7mgdBlTPTKywUrUkUTVjEm9vuaY7AYUSsYHoA5vqALFTlWjdvjhGUkfP8HbQp8oCTAJ
web1W+7RGJcOT2uAbINcnFjKR8WOR4ZSK1vUBJW9V5dir1hddH61SSIlKI+m43meuHguZB3ukkrO
YzUtj4AlspP7JOLmlGjL2HZ5qiKZLjB8uj7fmoYtWprv56IMve6Ov+bf/IgjuFxotvh9p0J7Pyiu
M+e7OKoyM32lMdvirXS2StxSODQi31kzqavFBaLA4sfjVMTs+J5EwhF2vu1UGgpnyXZCMweIR+h5
JcEsQY6P9hm64crEgQvzyShvxJAu/5F4mSy2Vzs5GwJb9OoL7Ku1DbdGvayBdWA7vQvOlsJUuVJ0
0/I9sDAMeEw3qxvTJM/zhhuX90QReI/ESf19JOa6PGf2wd7HOXejUA1J426BUlEQxUXdV1jrJd9r
IAadD6aI/Xz8mnu3q8Uijow63uB+i7OWY5mGYXL0piXfFm4XROErXBtvnCkutTEUVKdWfXxQ3uxe
ah+JB/W9KCs01Wpwfyng1l3zxtE6U8/GS99t8nVzgAVESzR3qo7mKC7W9+qcSZ8vC0qio5qUcDvx
xCBK+nJjM2Zn5g+qNsYp1bfWG7KBDTPoHGcxwRLdLC46DfpvXPtE2HsnaBYJETCdvFZ1f+EaWiJF
OuY0IRGKldfs+HeVIpPc1TlbCfbQGcfDh7S8MzVIBhFdwFVSH8UEjAeoEKxK4jiZOjOiL1FMYoHl
lptOxW9Gf4+4+dkSkeI0OikhKkBfMr6/y6cD+rStFWNEf1q/uH5MdUHYe89L+gAUbE4Gy1xLTwf9
pI5j0EOdm3OVh5lk1PP1gw2r69+Uo7TSfFvWINR1I76cqfdWyvVwsdfUVu/0SwIUnIIOGA1guui9
fiDjmm8BUI+OEZFcv3pyvEIAJBWmcLwfgHbkjPIUBJEbw+jNEewyuISIqyUFe2P24o3DIjgoG/W+
AsaGdrDXAmlfi9vwjlDItkY5TZZEbZl4D/c3F0HiJv8eMKPsn0pAZiZMdtAC5G/HJNQYRpg+dUYg
v2FnE5WH5aLNrpNj++4FtLxbVaYqx5TeQAuXJfWHFD7G9TsBTjFum+mBoClIG7SW9mQt3g7ENvGJ
CVNL8jNZ6nj+yJPDLZpkklfjJZxqGvZShHhEz9XZ3p9Awk6HW4MQKJXJXFJpdJBvjMn63HLfhS+4
aIQNWMfBjmFQ9mMs2WN/NobfxRi8YnnOtDIh9zlH9FKyXMScpaehq81HWx8gHmzaYWS62k6K6slo
/EiEQ0WkfL3cLk6toagafkKp6U6H0/woaF6N3uCzYaR4/26ONKm0cJm7SgIuU4B7RfoFzfyv5Chl
ULhUMqgkGfRKR98oXp7vcW3fjRVhJJxgHPaXTGNUq4Xn6NT4yTD3V+wTwNfv9GnJOWKZmAaeiiAH
EKVTE1LwOgH32SWGqnGfsOCPeAtt7mrNKRYjJLLAbCCPeEoPXtgeg6/+3rZUQv/ouAyILsoTe7lN
OZv9fadn8vwo96YA4v4e5W/pTQdov+JTGijoE9Gf+/XDpbWhJgKM3kTeFbwjZV32L9s6rpVACmnK
GLU83kN0Uzgkpx5HgPYJWWAKXyk73S7GQVEzfjB+86IsMSm4oCuaD4y5XeLYSSrW+Ah9rQ5qVdhX
Vim5AffWnifqwSggDbncXoLd8dkbGNaZTG5iKtvWu7NC0yAJaq7cmaMwUM/4ecsoZeMxNhRuAiiQ
Lq+M7pDpncuy/MUtZtej17rs0MHlQUbzdsNX3n1+ELnpTl5Sj/txLDiTzsJvBM3/gdZtnOmguyy6
mO3parvpINA4KYSJ1IWHnIm1+YToB7BMJ6rWJo90JaImeWH6/jw/84Q6pCsGlSPuAJgca+4Bttr9
bW1a2S/lTiSwyya/4Wgh6TUP7RZRuhcVIWFlHQYo1fly6LKMjlnVnscklDGL/JGoC+AYtzD6BzDW
v3sMVNxCvEmo/yZS91LbjH99IpBYw9hUpvN9KqyP6bd3vTgeFYhogIQ0eqmZo0q+0LSltERrmDtV
LUFeKKp2woEqN8INWgwchAUgoERXmfVdEKFK/FlS1SIa0BviZNG5ZPUsxph4itc4rdqoqdH3tqYI
I1qZ3nwDrALFvE/6zYDdSfbsvqvhcjnU1c+1vgZbMLKr8Y6iZZNme3RkziiCsF3gbp9H+qMs+tIP
/i5VYN0W1lOEnIb5VZwIsWp8GaVTPvooDGhqm7O90Kpg6ezhuo+d2Tsv0SUeaT/ZdtrxcKwAvCqg
i5DYDcTr2/pIOqWYs9M4JxAEEmnbqPvKHhpzavxAJa2s1BwbpJXIPp5QHkNXc9MRkmE4Ayxu60ei
StZbfCl2XvwRmtvO6Mx7Li8+H0r7LoPhbC7Y7gCkwlltqu7n7vhAuuUqdS7wRv7WcIehQ7b5y4NT
AGwrLAG0pksPYDE7kFPO+S32ens+Q9MBhZdb+u94OCsyTsgzeoXi/xomITSON4grRPTL4ocIh4Sc
RbziIfTp0rx3T+4GdkCqEU9SEgFwfP8v4eVn5UiDMXk5mra96oYDEpQ/yuPqPiIy2OBjubJ0EzbH
jPji+9qFa8l1daN8kwsordnmliCg/w6Chnry+j1UnvApvpkK/JiOBIFcmZVnIG2nLH7FrheJyXZ/
kLsUHNPfui51/Valy+/e8nITYdY1EcRhOat9YYDrSYSTB/zxgFevOOEnzG+hkB3MvikAgpV0TSni
QYJ6BR7gH28Btr4wznM+LeTC+aGft/FXQ+K5EBkm1NSyoH5ZTzu4YjVHWT3oZ64oJOsSu8QivOZV
YCtSi1GMckY6TdBogCCJhUVJT0taF+0e/WMP/Hv3ry8pzMN/0Y8ZP8rowh0QCIpbaZb8sU9Yqv98
cBzGZVI/248yvhIwnzrT3qQtT/xJR7lpI1dmiQtNI6yN3HFtqa1QcinKXwaM16+LzjAlNLQuneho
OustLtbNDd8p0K+192Fk1AvuzQ0wy3s1ypfvhJ6+SmQF2IXNHCyCZox1ZzFDSnzF8mDXSiz1GGee
T+YfUGTRypBMs/7UIAoW1Gq8Fuar/HZT3lqbQCZuzMs8yhGu2LUAJnYt0XSiR/Aau2EsVsmmF/pX
aM0wLcO8aEpoPHEPKSC64KjQbP9Ag/chYt63B2wHQwj4Ptvay44Ko7+tyuEr0eZ65ahDiZSRyZUg
13M+rQ7f6w9djO8DPNCZmpVgibPJ3NpBHr4nDBw2pMji+MMoijq1ahy+njBV33UMb78nsKEjLc4w
te8Yw78a7ZtsrL7GfxlKtmk/UBArlrxdG24Ylrt9I8oWI6pMeGSMfgr8XaUh+jUlvy8StLQ9nj/0
a2Ci9eNGCXxvMrBGcU6vJHnRd5LftxdrBRofoQLDVlQ2ZvqxwZ36zI1EQTmvqTU/P0HZveumyvuW
lbboTMrLBk79Waf706+vgIK+nR+Xvh73gsn2sjzfLowzgV88O7aRNEHB6UOnzwNvSnTQr0JETe/o
SkBWLuX8RtstrYwo/5mL0dM6IdkF/5lywRVLjRoItf9c13g7oO2Hk+qJfzjlc5Faj9jjc4aHVNx4
K2Fw8R53WxTBJlRzD0wzBfa1/ZCT8vwqCDnV1QIW2T4rZUB8vTIU5LbrDCY337gmqrpmjTJe4may
jGupC5D+/s/UA0SLTNSLFrGHB9ZiHS/LtFF8judUi/o2LWMHtV2hiLfQggCAISY6uOmTckvobsum
FxY8vxlkBtVZ4IfP0XyObmEVaLJpj8zeeqrHoJfJEhtCJR96Ezm8K9B0j7ejb6s/Xzwic2/BpIev
TGVqnwlnPseFdsuz92/ziaMCtyRkRZsqQssUVS+P1T7AOIm030kRZUTVMonzqNCxeRN5HquavUi6
keQeAz8N+FodY87cCnT9E2LbaEjuQr1Qh/5mwLrEXoYhx/BelUrq9L1lMpfxRut7amgvvFOqBQIJ
obl4FvD1jQ1pHmxfH/CRSH2kvcrpL8DpnNWh1Up//VKup1S9eFyYRHyPQpYTTYac7dINjuqYXfo9
sk4S7keM9aXyjY45LSDABlZhnkXkjrdVq8vh52VhZ2e5zNfAc/1wHin5OnsSOXtEhVKzEeIyCyfN
Wp44rbniCgDKLAE/vD+JgDYuOsEZ+zn+6Nht1B9cpWGmhSSoxEFVEDgS0Uhc+9ZG1GBvFqMMFanP
7i15A3B79ylMVOVpgzT44ZbfgnSSpTweogeGxNO/BKsWJo0bOBDvCOqP7hzLpHrcSN7wNND4wwKp
HwArhnFyrd6qr/0H+Its3Zp08gBKEa1LoJ7iVmT3WClHGxbPPaoyR8DAVcILFkHOf68cXQbyOLeP
vItRs+hlj+8UsE2rnj/w3NwXGt6rZMLespm828xk307AuRFe+TWmxQBcp0hNRFFxSzSwUh9B0HbC
X2KmA26vZMNYxw6f21ZAqa7OdtRIbmxl3HQ8NNorD6DI7qnD0pmP/cq4YrbDqI05f2/DxQnUUD1I
uj20n6DDTvf/X11vx/xn/ka6ohOyoNEbTcBdY+L/iR99sUnrcmWP/MVsy1uX2AhnM9w/xJnDyf4N
hbfkLKgeomcNynlT2dEg2r0v94zAIrMRSsZUfYSvjgNKpxvjNYhH4/Qbyt++WjRLL+L9XpP99PEx
d+FTfOHk9k2BGdjY9/KQd4ca5hm1tpscCF4lV5pthoxJjDrY34O8kD285HjrTCoFaZEA7yqTfuau
l5KhgGOi3C9mBbSNsYv5hpHvKyWQ+vXKD3fH2KYRZfATEYQT5U6inPUxt0Q7tpCH3KbA4ZI9GNS3
VnYboRUgy2YumTd8gDkHEp7xy9fWHwulVWpwY/GxAElUhjNGOQzOILXZ4OukSDxxpgv1116EsnZd
CNo+bpIPt9pkD2KNiH3Aa86c4Pe6I+Ngf2+UahyUEXJn8DLkTIoRpZcluwPvg3EvgD6Xm8WwLdRz
W7UZ4FqrydcU6AYPUkRwEtFk85eQNutMtzWotpyAoje56VTksaODqR8LNe8DfCqZkCqS7WUuJAIb
FoErXZqceTrBWyHmZgBFJ8huFPorEfROsNZINIlvcLtGC+5KYUHh6KEgl25siJ3dmG9kjCNgvgMP
JhBb5jiHUXwdGL8ZEB2SsTARC9Cw4Nkk37+RmbNuYddqtKWbCLNbobM70+1avoTMiMdXmdpziIYn
Vmc455nOunAanK8YDqwkwtMfVut3mBdYY1ndVFFuY953/pnjFO0UiqdV6P+HGm0rTV4jGLY+TrJw
ohVXk2CldJWtEfhk+rKc/wZHgL1KL3RmfXNDWJb9TFss3r6EGGaCpqPmuogSiI5D2m+9xCdFKzpD
UNMK3pRloiNjGIcMsKbThdmXQx+6TRDeyzPaAElCRwcMN7akfjMOluAtP6IDJxY4KgXrA1KRronL
w1KJCz6NY4IHkDrBrBAsPnEUAIqNfpRzKdoSkeT8APu8tnurBXLl1vf1ql16/fCKTLWf/YUR2PHB
oUAnBXVUNbAc5NskK4N8iJa3LTW8JW3C5lErwYhMDKTy3zatc2vSQRz5GYv96dfO/ovrY9jcjvo8
hgL2C1lxdZ4kfOKmKceiBx7yHkNuxTIbwaaOL+0Mg4wlLrP8k6iu+4pm2gilynyJsWxEVWfGQr1D
LykQTh6AIrrM20Cyjw3p1/kxNj4tlnVYoAVk2bEQ3AD8CJJ4Mb0F7eIWfbbVP1wccNlZLqCSW4Lj
+Ki5427TSl19Pq4nfHCmgOEXTO4xiJkXxq4vOMwr0ygWRT5vlflWUpXn6k7/pre4hVwNdncHATJ9
awsuiwDZVN7ZkBpFtPtY6suiv0rJYYhZTI/mX8AQT6cD7d1skAzDyaxQejT4Kti5CPtywszjcy0/
ka1jEZeWqLryMYlNNDi/mDwLpQvkOxB3lFgqIXCxFzYo8orPgFwjyNuZkRX6R2ivKCcEMhag6Pjd
CMCzwK8616LV+/kXzXty7Sx2gVJQc0d6lv9F5RNA5esI1M/0rCNeF6TnGCyZHUZH1CAe/2mmShL9
eRO+WDI3DFFrVvVLIhg6sG+wCW0SAyLiuijvgTrInoAGiRyE4WCA1R4XtKbtOCAomKPBWBMZpc9r
bBGSqYn5ANSkEszRQmX+nHvFao20pnVwoFrWcBFyuszfzl8UfVUsR7+jGSCnrIx5nN30ssk6Zg/6
OB0RaA1jgbf4Sm9OZDTV5HDY8UKDgdoIE0QbWw+Wbc4oH59jDRosYgPnwZSewIHtPU2EEZvFz1Qi
hXtnvylbu82B2dEJXfvT1tprSNMcpib9IP/zL3DuIX6WoHSWar/jiKi4XoUTjcVggiAZyJ6iaeQq
CJ/k3QfAb1wowcKKu6vr9lnWvBJrgf7DHwUpBv3WL+ZGRqQAnEhl3ZgjST5D6qwCvWsQAWdIp4zp
L5r3dFuRAjw3ZhIhR0h92OOO1Ez5hBVHlMES9ffr4W+FX151qswTwOddnT2iIAzBedrnB2kxMyot
k0YPhIL7qJZUvO+Zx7T8M+7YlXgiV2sA6k75JgZaAB4pyBaQaHes7C+xYpzwj2bjA8Nqr+qqVqoJ
Gf1aMlAqwJgUa6GpMhczNLsk1wHApEdIvxIzqjQScFac8fZlYCfkB6Mh2OxSjGEwq+kcPg81wyV4
wXz9x9j7WZxvNOhXvHqhIZbjPjX5T96sZ8PBLPlUdpEppfV2yal8LSd81n6mLWdYT7+Av412tN1u
+FqJ2RrdIc4UQ2XAHwRNeGcfPHeez1ja6gutS98aMk2bFeGIMnO7PgeXoHKoitnTwTwLwfWW0PtX
FmnLw4FunolJFPx6SOK4VhjKiG8Zki5N8Lm1/wVCcXtX6IMCwRS0TK3xB2P8h7l1zJUdiEudfeFZ
DBCCJF5XeGUIrNnV8FpzcGZN2Kio+aYfNhKPtj4Df16HOh0IY1Yzs4AvokUykM9+VAIOHQ9il+iQ
o9+NZWSeAeQA4J/26sx7Qrx7b+sePNH34Z3ZKnJywbf8R8K32ltUYIT4FK0YvS1rs60AU7pbMA+F
fov3EyCG6MYuZ3W+10g9mUk/hLH1ja07y6CJ0ld2+q0BbWl2bT2bISFPWJye1nlZHnQDEPAa/3L1
l//QAmN0mIiJE40czsBquRn7QtdBgk8a9KJGY6EHf3oFb8DMaPCTmJSrA6irCY/keRRcitqB7x6m
KRaSGbJ2rnD3iKmMHTlp4ZgI0UExlLtLvldIqYptiOFfFogl3XBI3aVf3s8i36KyMLh47gowN842
PWZrBWEJ7W5/CyrZ97NZXTQ0UJgcayjuHCMU5IJpERDw7C/QuOwgXBVmoQocpc9mrk3+GcwRlNZ1
R80xgl5v+XBnp917a7mR0dgI7g9T7/24AuHCN1gUZpqFvJ7+Vx0tkMLwqzG68vFGWtamBQIFCG+C
CmVGTsAP0XnDHWz4humyrC5/3nuK9iWrHQdMtjcEjZZn/PY+rHtVKregCDLj6sTtyLiuFlnkWWmN
hYcY/IZIyDm4Oi5QNvzOCkGdwj/3kspn/QFvUIBq8hnHN7ktzwICyvpOvSV0RQ2LnGb9fj358gqu
9i8aKlqllAqpofme14HLMUNu4vZexSbEinrs6aUYin2hQCY/U3+X4DkiVYWRKMd9qaZAUBQXgd6O
gPwWF13cV53bvPZGG0Dx6HUq626OUSRoL3jG6PSCr03d6SQ1Tom0bk08R2LvWJJyU7KXCA/t5VX0
h2dgcxXpSyV+LsW8EW2qs9VVPWVcw6pQnyZX3h0DKOlVU0E1nVWpGofU2gXs3Np3ulVXqvt3J/hC
iJRJJe7ESJ30q9U1Utt1hNQpQWFQxMvD5vbU7v+HoJfxcQlMgbq3n1Br+lRGNO8gF2MD6/Si8yTM
xNnb98rmXx2DcKHPuoFfpXWtSvvYEX9Znt08u93ILaRK/4jinqexTT4T35bvYwnEx6lrJTOp5efb
fjqB+H3BRAOqw3libMxzsWHLwljlKJUF7p2q0noPKY2AwBo0UV1x7+f7RDasJEW/pPjwnG3It5ak
RHwFCohAoqWWr9MGDi+T6OwXSmCT0MRp4f0Uy6Y12LIu9CE1RPkuy5eVpVvJisj4qYmsJ45LGaIh
+8Zc9aM9qJVNg2e+HRqzAX0EsE2vYQsQdPhjvSBAeMvDfXAYHfZN4GZ5njlOQkmpDMHjCGd36mhI
dE69bL/xAJLzRFiBnEZyN8qx2TkcmorBHnb6ftpqmb9jRJgmFX+2tZ9sl4LG+s05nM6V0Ixeqb+l
vPqQ2Fbfp5vUrOwZhzp+S9ZvPiJfldyxjkQGrTO9mCHQxCcmkdQfVSnodvcOL9Mq8Qmon3ePou7O
XmHrBLMz8gWQ6EXHxfpt5OJzltQVCHZERBq+Ns51Q4wAdbEhGe0+nf17xl3OkvcPBtbGkqKKg8VO
Y5kYnwjQzEbd3Hv48KuYueNfCi3S35ouYlcWRxYUuoAfGe0nzRAENVWc3411G9vBxzjFI/ZD6glx
VD4NIvysYhY0V4Y53F7/MxMJDx0xHlVjppEFwUPH4vVVBjqYl7iKgwcZKYSuWQTOy/fKHa5RBwAo
uYMgvS3YoIXwL0WKZrQ+kkWuUcebVgOHUmTGy2ebl88zE+t4eYZyGADSprYIztc/psmuPZGoJZAN
4ktHfM74Zfkr3aQ/0qO5cqcaLWa+TZ07gIEhF12B8tMghonlWhQ5XAY96PIvCDT14TyV/gf5ywCM
3O68c2t09UrkOYugC1KIFKXoV7dPN82eYyd/cLRMr4diOPQJj+OkyS8CzERu9go/DgKhTvImifTr
vuFCubVSa1cW0BR/ZDi64id+kUD236dFzYun3Mqe5gVrVyNr2Hn31bX3LExM/MQ06HsLmOGaQ/nd
geZ8AKWx0vpVTdgXGFzTHURMQptUtn4/XUusoZw2oVS7CRGgGRz16tsRwrgslcxqvE4X/56EayuP
oz20ztjxOjqiQLUxZTuFUv2uB+HjzV0cEqCBV1GdkmQ3v2d7yHnffiWeF5ghMFlUE5liOUzP5tve
HJyz+gPE9WglmdphJ22ga5S+tM68T3xsvT8QZdTrUyauvg6tGX6W4htNgoC77FGCBvFN3GO6pCtO
LdWPKqr4WqiMA3pFmz2G6A2RgVcqHPlQwvLhS2LIdmSBIZQz1O/XojUuvZ0Ym/IK6g0T67Am5B2y
aHdlOknj5Qz39RYexVtF3lHhHJ1mvWWl7XDbOzrR2rJtI+ljSX1K8D9DQpoDJE+0YR4VmFAm/+jr
3NfcZPrZj/kBOVSOm/S0ZSgcZ4GfxJ8DZZ2+vQrmDA2AL0AlPsSc81kn5gtVmynwp8lhQatJYAvd
2XQz/FbeKbGAWI0ImM/IvG2P/DZzUbufCx/Qh4ursjQ7GMS1mwQ6BfXqQWB9dJDiE76a2z7zgX/X
g17q/FILphMEi2O91BFtYrMVnPZ6YD+3ZT01/oUnC2PR7MxVBD9GHm4c8p02MS4ulIfUwWa+gzFT
sBw/vPp5arfC0xPdNRMxzMTT8FYAuuq6O+B3A7EIOugvMbxAkGSZWZloxaaKtBbWks3TTcp7IqWx
anrLqL+43YPooxZ5jXx0V1dgXvE41fPVCr+FT+1KQbHmuoGGPN3iD9xvrCcI6MljwVFA9bnCjQmG
kt8X4Vh0nQdCkCAZrULlTGW5Jw9PfSNPwclCNuO6+873M5/CnSrLEB0x92mtAU/G/G3POXDD+Z7s
GV+OlJgSLzhHl1hA34rD+8RK84OHg3A1LKXWPqc2Xo5aaCK3symE5p6+f2x1BAqqvGH0bUrfE2kg
LC9xXUkR3VY2nuaKIIQqaGv65ofTFvfBofBcSeXDon4TqshZIxmwFZz0E7kjm/vJEBUKasHDd1zO
12ovrLM1pu9hiJTCKzbTEg3SCeZLcVIR4/4rKkfBV9LnwMr/Ft4YqBq8nC6VBtcFLXogXzqFAZCZ
ammeI+2lrUyer1nH6g1OyIAXTJ0pRsvJ8S9jCPNYL5Q35FI60xERbwk1DBdgVc66rRGIZVtjBbcO
UJwi5xsvoBCyWP6mAMcCFB5SrUbBDEUjZySl2/YOxlM8f3/n4L++C6/jxYTq+VJejDz5UYppkhdW
j5jfDr4fhDW+8Bq4eGDxV7jWA0vbATohBVMtXwszvqeG1HhVly5Boox1gYAp5O3Vn2YJRabzECHH
F/DDVhJ09q1V5UA6m3XO8q6TaMLV097UJtQvXUs32kXt21tkLRf3zrBqWgg0zPx6jQ6M4HQVvPBL
iWk5EY/u/lcq7rKOOQIN18zO8p6lIi8PDe3nN0FNHkjPzcKXb35zkXPQq9rIQ1AIDF6JYuz5jwVn
K+SbRjnaA+bCiQJo8s0Ta+SeO+tsuMnbmqh3vzvE1euGMmlvqZ5c+174javeRp2Z3u581SzxtZr3
wuMnpxBhY9mtpD6yYzDnzO28Jw1aB/RAtcduXfnGTpkPy1/Kqw6OFQIEN++pR9Y+va3UvOT521rh
JMt5UZRBpSG672tfqeqLfrQvpjFBPOrctpQHEOsLQh86LVtg1+XPZ/JFABkgNtRVIZ0A621A5cta
r0VvJ/04/BtNv0OeNg8WvJguDoWJ5axLZosX9Qs/Z3bLGHt8H26YvqvAnkrm3OmhlXmh6uRQJSSt
JRe9yMrAPYHaCSgCEgu9MNG3ZY1Br0md5DrfDn75t+lWXdnNZwDkrHTLHe25kU00bbyAwqy1vwIH
6EX36MtQ+11Z5dUn9WGmpEQw/Avi1ZWTBMaFSyuKq1U4zIltdx1Q5Fv+uEKoqEVSCXIn4EXo7mNH
XXRWtkGHofNF5Do7OLyYYJclSDGaXciyoBqc76btbqYuMT/jNsSKvpjQ5PPE7FS2QNwEehCk65t5
+NIhUJz2wW9m8rQBOa7L1B/lbeSKq6qb2RvM0+w2KwGDL5+zHG3QHsTWMRbKuRDLEQ/RZ46WS2zF
4pzBi2DhI9ijp2uXXMDYfAXFWXt32uPGkKlKTZc7GJ9qgM0AurhCWR0oVggOuQDEDtp6dr+rE+pC
MSFCxckmcniP66G7eYF5UxjMZQVHAGQeUHBbOaveVpiBP5RzAX+v0Nr5kcW3CE6I/qj9ot24PXe8
YqS9gsuxiCP87NI6+ztQmtCH86ghz1fZM8auZu9hW1UQwAwvKXkxMRFPzNdEuVk1T6iYHTvzad62
XxZUCxzjQGC81xjGoS5J25avfykwK63WdGx5h6PtHH9zJvUNrjmr9pYNXDx7Peahq9Y1H08tQWMz
F5RZi4YKBfV648M8fgXXyWhLNeG5dgeg2Ou/uzpy7r+pA72A5lzfmhzOxfOtgQioJivwXwy5qB9y
ESv79tkwO9FE4/pkmezuGFiJbyvwlwyRXI4UT0mHsINDjZrqNhO9ZimYlrz5CtDY8hf1aQRzPOVx
joQynQIM57SxXaXn0H//NEFLZsHsH01po+feuWgqC/7AT24eOXfKHtRWHhO5bVPfCXuCcYeNkzNG
IWBAl5xeeALtC/K8EhiuOch57af0JmTfRI72dc3AknI7amfwdvQ7b0/rIflgExuqjcJnsecyN16P
i2Uer5zHZ2JN4J+bCKCaAZIIsJDSy8zikvBzV4cOfBC2ZAY46KsrxydY28F7YNDdc5r66mxz3Gpc
Ya1YktFbiqdhMYHvqfhizR/l/qdGYvR89NWrNLtnEmA24vXXU0l+xdHEYJAFUZlax/2tldBwazM1
P+EfynWKndOnmTcHruTjO4TJormMXhxSg60zWGms7hpafmEkv8M++d6xxTx6lWChHCanHKZoGw7K
UA/1kv/uL3ei0YhS1rZoijDOH3tW382u/oKKbMBWsX4vQxl8ZBOJwxofmRcEhTu1LeeGCKO4wMDF
/nWYF9A4kmHGIH8y+QxvX4pp+dQ+YPKd35vtRASIRsZyF/xuRyce4IZr39b9jesCV/kynXZy7IQY
c0rZAzhSfZwUG4yB705fXbryNYX2vGtvCBi+lImSR47J+SuumOzv3nl7hg/8TeMZvZ2hMv5EtsVe
bj8HvWZ4lq6Cwu3EuGptdFhFtDejJklvbAe1tsxFtODW8ggCPBMhOxiMaA8tggjMr2NwvlGFQFW+
ZcMu6l8uUKkYBdc9RzQSm7SgxjNGp7jbQVfIkeqaMql+8LKq+lLLkawE4928CxP7Acgy+U5GugtV
ac4AnNO7Eq/XaOwDwjWQ7mXqqeEulc6hWYROj9qmxD43tsBd9zgOfnV2s1BSgKOJlaGQL0H681TA
JCiMMQEUUbl59CgGAxaRrCLTOd03aMNcAHPxzDchYoFJliCmo/1QfzXvJWCNY2aZrIqUAGjqc58e
LyAN3Ssdw8FDvAy4s/2+Y3A7YVcUznzVil/L6xKKOjVXFvLW/S6u7Ii9J6JehlEL61EDOr+Hhn3k
aagw6CRgAHD7pK3XIBtnNGSNFliUFYBv9TmrebnM/SKQWg7nxWvJpRUkEUhynOGiWipjESrIO0h3
bsP7T+WSque0SznYK88J4wlX2Wqh+ECIvlBD84sD94mePPCXWyTcHXWFtZFWYu3t6HjQJ4Lnw/f8
ej9UH++iF6wrQQts+eQ3R4wahKG+rHBgz+ICz1zSe0/g/vTazb3qKFgfacumT1onrBR7e9HVCvbf
4asQeIF0O43Y+9nIafzuwb7seXBk7bNx43dSQzNWlz7ksAJ8JUZn22+3cj+59c+BS4mt8pg2gICg
NAhELM80n7gSlQmWKLHoSz0jwx7qV4P4+u5lqg/baHeW+JAtFXYJMGW0UmxWficZhQmGNE+ttJWU
pRJZiV69KkgVt4JZslwGVXZIGQ9J1Q+PBWbwGZu89sncwaicsJMIgKKM+Vlarvy+hqAW0KPBTo4/
NViju27zaBe+GYBPT+llyub04afeOp3L4OKv3r09g8GJrNjoh5ATRoV89Kh/Wn2WS3EG9CG73AGN
N9qSPqOMgTarR/pAEkikuJWJtrIi1X6Z8mMiKdxT7rsqxXV2/A+wXg1p1xfmsMtmK3WOxexKra4h
tUruddm3FYlnjhItZd8BlibweLIrVtc2F6tmajDHlZfSnrwJ+HDSU57juhTzBOzSUtPAqoIG7y9P
q58VgPNf9XgYPY6kh5AYuO97d5zHAni7gjwsmS0cveLcOSCflNvYjvywGERyp/h2IGnm6wI21V/Z
SGzzG9qSf9jzsWcEt9jHx/n/rzlith3wME8++mkL/0KQPYZknJ94KA9vWsDtLR5zoOhrjJolUfRu
rGzZ1A5pG4OEzNmzM6NsDeP4eeurbxbDF5j3wQZVsfKSLuxreCLgxdvMY/taWQusRWKfnSj3Z9QE
3rn46np2lU/Og8AzHcFn53y63aR8SPMVMkghR4+o2ULKTd2WmGJpYBkgD8ELAOIszs6+KJ/rfEQh
+xD1QiKhv3utPXTS0aSj0VsqXdCpdxjDOoGhzajg3wMApONfqrgjSn4D2KjMd38YjIMxH+zUGPCT
nqX4jXRuJY3D4C5rMpZbVRS7SAJzZIrdVsQ+7U3yKuOB5a7aJOa5ugXZLA+5snNq/Arzs+RNd0sN
moBPVin/9LE2rbrZL2s12gJ+M2kKIlX39nKJ7t3HJtm/qP5IseBCEysLNgfNFUm5CnDEYmdVqRKb
jOziJLsUWOL4+nr7YGEDrSlUnx535PBQNW/+b/R9xFtz3/2qv45V8Mmub+UYDLqFvVqZMo7TnGPP
OhYxPYMIp4jB67A3xK5MheILKKRKYsNpYRbiSHyNi3Ki/v0hEoqdY6CFZc/qGqi9u8e7xvOWapSL
ZkbWXiMujGnHCiwlXwvNRH+I5PaarnKuMIArGmMbsVi0v2xZ7wk+2vh3biGsBqjm8d/CorEdfSyQ
QDL+eTaGoXUE7cUqdSHr4WufSqd/e+OrEgEEZI5AWFwOwq/VXKclBR+E+0aITqXOB1y5MDo3aqnO
rWXseIa+rKA5TDTr8CVn9Cf7c5br18IIkRx2OxM2ZSeCVk5lSmQhS93KEqkEU0rt6gLCQUqUTVHY
3bbDZLeVpZMWnscBYVshxdHL0zf4ntVPU1J5iXp9lx2H8zDWKzneh4WQpO4iwaXh13KCcL3si8gy
zkt3cI66IGqciqSji2MuISh9fEVulFHOodZvhU8/gtbPpsX8k/rMJlSl0ezxr2rQrwWGQ1u5ob6i
O02VFMQn5SuMylwtTCQd73TSwvWzOPpIH+kdbmO7oNOlirMyE3TELT41FRFrUPXfvVPvfMbomWJQ
/b69bHffODwAkNyGj0JiFhfbN7pvph8bLJbW6icO2Gkr7Bj9X6XVy85kNd8kxYd9OdVjwWsiGViX
PHJFuXTP4Rv1ihrHc9Trj+u8C+Oun8BH76uMb9AAQ2xC6LdcyBohRjoJT6VvFGKXu8VnqbNETMxA
VqUjSurnY9HYErnydLh6tN0wJzda29zXNtMMHn7GVh1k2GmQ0hxhPSvHQU64YVTgBIOtHDiPbJaj
fMif/mY4NMZunOLJZxlZsXO+k8PkhxxSLBzrMIYMvibJY86jmbKv9tE/QUtxy97u4gGSMyj6K6zr
/FLPO53hfKWBn4Xa9nnXUVDDyeVmTIksFnnbJZbB2SZMsUq29WzChAhVB8FZIR5PnSZbZbNjnk9Y
MVR170IdtRq9z1E0xJqEssHpk1VJRCEoBd3oVyuor3bdclQrLTcSv1bSuBZVPkno7m1d3bXiWVHS
ymDTrdO3RKD6bW8wj3ahXkVQzUCfkcCTScxSQmoMhUM024rLLKmkp/8gzTtMQtWcZyYJ9yNGd2pJ
dpU6UHZSvncfO2tZm9Q3tEVOf1uWRnjJbJh2BnX9CnW5LuzEfKfEgopvE2MHX0B8FOeo2x5/s1r3
RYJqWg5kAm2AviYrdxVlVZComi+K5mkVLoA9oIq6k9mvz6w/iDN2w05AB7J7Txt+ApY+CY0Se+sV
SMUBPG/btyHBdNd/+N32OytM0ps+3unNJpYD4KKkWkTS7QUuzMTit8zpa4sLLkgfAxQT25oW+JOc
NwneaqA3jkbt8j39dIjqOV4BQAgN5KTKobJz9LrwtGLkn5joRWMmHcELH9oWmC3PepP40ofZxm5m
BwVHkMIfaqj3WMP9gxfk4AY/Npv+Y5FWUfAkqMz1m/1fzoV202erb3rr9dn2L//0HGuoQsANud1e
HX4TWj2exRaBV1YeEk3EkNHg6OTbTjRMqKzuw3qpQ6qnSelW6357CeQhQUq6MF6wAVtmvn4ZDvAG
Lv2ZuxSkb9jN6ahy+cqVRn+eVvq2M1w3iAABeEXQz8GIMyf85KtNg5naPP6p6JUNnuswZFx30roo
7+bfdjGavS1h4rVo2oDgHf2fnZ/0t759Q37sLpKoOP0y+N2VHpY+yHZHRV6F6AxgIdLl827njTW/
U18viDAVOxPxpPaBeo01LQja5hNwMK8NKJOC1EXA9aoQUOUk0nYQwP8pnEk09bhKkXgkBfhmYpik
u7KqG6N739i5YTx5NSCKyMOsR7RW8ffszJ21E/89M66Lxa3T6SD91QDoubhElHeDSLHwOBUTcDNp
t0RTLMkvrILf3QiCfWoaCtvJm3c94Bj8B9veMF0UMAn4UQ2WWYqQqAnx2VFVz5+KoNn8ghRTvcO6
OF7ZVwpYhL8wn06hWhBRvjam8/rIMv558iJcvGVKjlsPZ6A4TDsjBjuyGQyNx/MnOLPONsRZnZtd
Q2DCHC+o2VsD3qc94o6DPHHJtuvBPS/wZgOE+ySN/yojqi5NmjRRsCC+Q9SzKMu9XUg4J81yt4PC
4Z7pd+HHm7oOVq4uXM8DIKm+imMSzqoK3kteNHraI9a1Hy8iuVcWNPqCSB5rNXzvrwJgmzOkJ6+M
1SUxI6cYrDe0AZdINsGHX0/GPMOoyvKFmPSd/tqusdyynK/wudZWYzN/oQSKEA+GRxvofq9OaTSS
3hc/F73qboxA5I/wG5VjvD8UBuuq4HM1CWAS/4ou/42jub6WPwVgavX4kkMewvP9GyCRtwYpYGOG
CF7OvY67PmVC3sJRena+AJtNEY/JIZoihz1jtHeOHbnNisWATZmMGMwS2YwH0A4Wqj6C4pZQCzLA
XHctcYFCapjS9iW2Jjl/2tLDfdn9dH4VGtjb1B04MO+8Q5F4Ys1wm7PbM+JKVx/vHRSScqTJ78+5
6YLj8kHthWKqx3hmyXWKNrztpaddPXLXpRo/sPecKzSS1HoafnOrdrgFneKDm0tViiNnC+pEn5RU
W7RpsQjHE43h0TtmzbEI/rIRUs2lLFkZDMUmWirA2UuYyDNwZXKYGlRvZcCvtkQzDQW4QcRm/2N8
3dhAk1beodMRsUkZQk14JP9nUry80R6xnkLSvX9DBLv7iXlPTHZCm7wPivCXjaXXLRBErosN463z
RpKNTXGrESvdVAKJKqhnqwtBfyJEpp+TLdVs2PKYaX4lV7lRb3K/nSMqYLybQn9Buf2dkrDbOFAz
SvPVKDAm+QWltqjDXPm348GP3WUrScUClsoOEW3FPWi673bOnalNgooaLRCSCLuo3GXst8taNvBe
EmgoQ7/UF2np55om78V/1Chw10dCmDGEOFTjaNMqKZ0KXMJ42rZJIgwdhhX6SPR0KsbTCRMeel5l
QwoV3jdRXzi5k1+ny6SGga2ItjEz9nF1NcuNyvueGjufw77NOz81RbV6DBAj/x3oVB5CT/Hq8foN
XpC5Fu24hKOjDCoirMEEoBd18UusIg7zCRDTX44RNx9SN8dhJg8/tH41M9/Q6S9XEo8NkQ476QlH
bTs+kGkU+VRBcx+wdvC1XWYWEqdtRK+Z7sdkPEIm9bjz/SiBKbiKKSnrVwXEGcKAEl5KB7UQsPtZ
p5M9HUq0H1a/9kzktyJJ5HaHq6vTlnxbuczg0HYDNgMt0bKouO2QuiQBm/OF1zeCPm3rZ8ajfLKW
hK/cZXVM+3SjL4bE8ywwKpAh1AL3lS0g5mHh+FTa/2fnbl81O5fFahCg6Kyketps4UGwt0GpFmki
6/7Fwvq0vBHRn06KOyDjH68CfzagEavz5BiHq2Z8FfrnK3bMvvTCJTqSWb6IZTaCxZPaKrdIrim+
CY/CQxqsh8E4QssQSNwN2DbEmAsVzuJf2P7PmHiIo4kvx1oKKlEa5Af+6AIBsAHVonygLEccUHMV
TH3h+2/SKaEM8A4uyN4xOuNkPuPyRXqdc9DWabCAEm3S5CzK6mhV24+P0WrYuZpmxcx3F5cj+0Xo
mhh+VY8gfwaf5Dlni+hneClFOwMF2ia7jJJvhUmo1l57jompBkVXH/3lCfYBHG91kETU7sztXTN+
oGNVkdiygz9qEPb8rZNxOpltZJpIWzWJp7TWFTLq7S8nt7Mfm9lYUnzrRuhGx+zp/1Kj4DolI84b
WpY8vUtaqy5OjsRH1vl9rmUr71l2e0PzkQTaH9u7ISLUBkz5/y5DrVUJ3EzgL/nf9Vdcdx0yFQvv
VSrZ+Z7NZa8taOH2gc8QtRhSpIPxoEFdZKI7CGP9Vspxozg56ML8sZaqM+bYdecYUCqyCkqePFZI
J5fsb7T6H2ZFaVNvHM/bgFgBh29hYRN45PZuFUS/F+jhqCfclCJzypD0f82glSTRthBq+wRmNfzE
IDh+DLuKrWP2J+g93bjUmY65s51WoPN+Sn99bvktRk+4GhXkdONFJTLONxjacHC39VGKKjTcyyBH
D5Fpaky9YYw6eQvw2QGuChHZFb9h5OXvZg1s87UCEY8dop3UinpJe1/hqOQvyCGnOnOqndL5T+uS
V5YX9l2pgv2PXVSSPFxaZZL6j7hgRuA/JQKEKaufvVh/mJVLR9qMWTiOLuf4ZDvetWuYxV7PKwo4
GoIhLJ1L0Tg83dycJp6hAHsh72JJhoaOFIKHy5gOlvn6Ndp7p3G4TelKE0ydSdCYVLCWyxplzO0D
NzwvDd1UrzmVQLhpb00ZFyp5HmDlj4Rvus8ROM9VxBkWC63TAV9C0I4g3ipHjdaN+mock3Gp3b8x
6S3wRdJF0Z6oI4JwCE4W2bbJTkpncLpQkdcWKdR5fKgXJbJn6dK7rrjoBELpX+oldnvfqM/XvoJx
hvHVu8H6Koh46dkELIrerlBmlmogIbx+usFHsym6n8zdE19/GKGdsOCswt6Qn8n7upx6kPp1OeKa
qeJI4BwDg6Hun9trYa3QxYcz+PFBvvvk0NhC69fr1W3K6wqSVUr5H39QjpM6VMW0D+BbpWEUt9RX
E2eR3m18Hp2aD8MrAKLFKsIxTXKRHUmex5Vj7+jqXpDnjPxmgs53vjSkbcKlmdH5LeVKgrBe9v72
b8bN2yV/B6pZWirWZN6X/KI4hXW2LMplzBKtR/4NJhkXF0gjHJcsml368+26JMxs8aIk/pKo47dD
+2/xD+gN/4EligeAQzD4yNiwGF69Vqu4Os4NeqhAFRxnSWAwqJGe8Scc7KoGzKxUVISm3lwD+YDt
QSAHIibMu1s8ccoyMimL2TbKCiXtq2XsyjQZwwL7DuF2w9yiQH79wMm8i6WcqjhLhg2CQYdqI8p8
26swlonNMThfgzecRBG7tEay1t5N4vwFUlzTvTAr3sIIJzDUQx9WzaQNGiMGIB/Q0rSIHKJ65n0C
zQYKw7fuCFByTTnvcB6Jl6/+hINU0KWvLAh7Wr3MkzPOzw9RPbNdTGWoewCb9sQJtIvjEPQg4IGn
D6WMxLFPRAOe/ysqfKbmY2bDRJIK12anEx1YOP5w4Yzn29N+TDnbaUf8FOaKCB9FomGm1Aux+phJ
Uv8gwGNOYot8yInYbJ5VTmz1VXaA2MFAVMOAbmvIxs1fgxvUVUFjD0xc3DpVEQjxXkVo4BBLZOtL
omVCOsNV7+F4CAhjLJogtCxHs3tX8DR5P9nPPylgN/WUT51KzAFzZmVbb/Mm/vt4pRqCgCuhimBP
vaAnCEvU7Tw211VajbIFwQCua1joLv5rGE6qiWYKPVyc2uVUcwP3vctVMZUpWMAjZVN4qocgBSzn
hozCvak9GmUvc7TBLshETKAbI96ltF7TmxeisPeNb+2vtG/KGA6Z4sKlTAJyDkRZjrAB3Wln54Yj
1WPNVI2PhWhbA0IMF0CJqFI9sDuLKrOpPG+fE3Kqo92zM0yLItWXqTpG/4HD18ATE7Qa8it03Y1k
yhjEVnLgdPgG1BoqA/HD3RJGEi/jvkTaqWL/sgzOQV6lRFsaqJ01fiK2zE4gdpmTAJ5bHppOrDsT
bfJnzapnftPF+gmkXaSdK4UoGVn2I5nda9ekZRhYrqvAGhAmiz+GnwRCPVWQquQLBpQi3qoiNBTU
XKCMFE0+lOz4wBkJXrWAq0cV5Np2drq+XaYzF2w9zJiEdcYkS2mLIAVO1kSexXyNJYnDqgYjkyUA
7f1anT3q1uFOvabQo4cHvex1k9ddBT8S/PzNgEwBMzRNQT/6QuDxIT1PMx+3CaDN9nkTOo1RL9mw
pJLz5pt2CuYo65yaOD+L5mPZMOCuuDHwBLr/FTmHJuGbDXFiKvMcXMDZ7OT2OYI2xl1AG3zTMZsK
Vvvam/iYzZyc8m7Z2u2oa1jSCiJyGYEaGKQQVeSZijgkyn+pRHWSADWNKzc9aWrKIKTMB9t9a5i9
tL0LCXs1nZuUrPRdHHZuyPkTfo8hh8hSV0kfKaqFXFJdkNndJimBKADyaLk5mCYZSTNaq8XN0xyG
mwyDUfZqr5EhLdWOwKcs8MssA4lf//onf39qJVObZ+21KPfXEvzHLVYDwXPrabFRMP6ym0KoGPKA
STwq3JBQbWFEgUNNmqVAo84FFzydLpGpJmr6okywfkjt4RqwAIrLcJE1IQPM0fOF4rw4MnJlnPbC
AmCs2NbEbpi2Lmu9/mDlvkI7sCBE5EUOEBF2UD23BbiQgZS2l55dwQnC0CHnHMM6F+Jgmr4bny+A
2h8Sw6eBKeIyjmizcPXoAQqnuzjoZrtRaSqrj8RTG1plVBtIuLzrJnd337tPf9JfLxASAPN+N0SE
AXPh01vOn05PWyp3YjQfJuyOV0De53Yg9J3BlTrsuR3YyzRajMo8JrpgMH2yddPVj67NiZBs3MTM
6SqoMYDKqFQtC4Uem595Sij+Pl4S1YI3WedwR9/w9NS/OmSPhLRCl6XlyCATSARZKoJhIRUaap4p
bK5AjwXGIsT8kNY2HAGuadanlbSgz9ZBxlfEBzNESJGxSvQUCqBSP9gkGMC65NvVzSFyz6Xs+0QA
WIRaOXvSWmF6DCo9jXKJE4ALKfkJM8pKwqWG42wBmbcjWQGSWXSCSRwNeH1uK0YTMwa6AsR6lYPF
GDf2R91kyocfNSfjq+TlalPYIkaStzG6rgWAfGsxf+yAShHh+YwYVRNDrf9r8NJGE7cx/XbYpIoy
ySaK6AjdwBRktZ3ushk9Us1297e+sK5qcEN/m7r99sIsdzjURaKq8CBXYtMy4P1wjb/7CXC/TF1O
bkvNNqiONuzzQIX0C9hQGrOa4hZJ125ibNzsKV45jpvm4FOFvVH5Pdn+Yj5kRRZDAdjMiqlhLy4A
H6QZt17OC9mgmzVlGvSIRwonVXkOS4lolQbvTMNdsefORAdih0pbQluZdf1/dLR5tJr25+93/iEp
ZhjeKAURc2VZ/qH0exfZVyzDIyZMdk0mZQR0WJVmBUwsh6H3Rg0EGXTYVUdfSz0HtmHn58u4tE7R
N0vB+RMXsc7Ubx6j62y6wTg0xrg0uOv8WxZgMToSj0/wytDy7SiyaY08L5e2qnVrpJZpHFI/eY5H
OtUloJW+4FJ7gyoK7oYaZ1M2wDISEOpCb9Eu+vF7SLZCp3Lp5Bz/cISqSaVpkq/vnOB3aZolZvj2
sP/Zx3RHjff3W3Ia5BG779PJC6RFXLij4Q+TuFedQgZnd4ptkoR1wle6Mz1hsXtP6lKwKOC93P0C
j7VWECgJNbQkVOXZnh1K7OB7oJ5xaZv+6vAWf8QdlKD286r8tXJIxSGgD/jHDQeZKAMWKA4Xrp23
LihmfTKCS/NAdmL6tLRZo+44LQS4IH3i76nBvzAeE6TdQBojguaLggUZY+k/XM3/MeFhe9cec0tG
xfQhe1WBawHW4xDsoOWsSKrl543kgn4hBeWmIaOHUpm1JoOEMKgm9sMPi64T+PDbFsZvOr7DXJFs
AWei/h1fAIuKAspelbiHUSm8/RgXcTVlvBXaXTe6XeSexsYc9Yf8nWpryWs9rRWZCEamuJ54hgU7
ygaeGBeelcMX8ILxy/YDo/yeW122rTZ1cBu17drz9787H7JyMDKIbxMhySowgQ97H4RFQDl4QHzW
DScVrSs4lWck+AEuykvIXlwVhTK3Zj7zlEgmoeJMMIUQwMk85xo3o7QXIPi6VQLrXl+zpTylD71U
oAAMWLezaaV8qJMZj+oa1Kmf1QEIvERYq5NZu1vVJlQGIl0iUODgkusePjr88YYiA2vlNFeEku2Z
z5oBoRn8Jq2QSH+VP49nixQ0+hewQ/jdouiiuRMBiiN8WM+ncIKmwzBfXRyrIY/4aXtvMXAOx0uB
wbdaHUgZ9qgmbVRxpJppzS/O/b8nwYeXOZ+6dU1NcrQJri4aZjImOcWEF1Qil0jADcTvORlM/33b
3M8wlm/t0oGtNE5S+RVHQRJHINf5v6JxU0l+maOAsG+3bTA1XSupdsQiZGZ8uIeipgKU7CwB5x4j
ZqTKSdJVGDCfttrEc0yXBMMEqzqdvZ83tJ2GkFTGn+E2QNTiz9vY4VavGe6DOhqYQfz65Jl6HiPm
OsJYq+cfvTfRGwmPhuM2PdBq75cT56lfGXoZEiTMiyaXNCUlILRxKYyhBXyoW02autNXS1iCZVrQ
F9lof9+dV7G0l1ujahcDki2BaVLoUz2nK+FZbq8rSLiU8eQKbO+2ytFmX2IiwSaOHtH8wIdcwT/j
qeoVWYHyFYoVQ1CAriUMd4k6rVNXYcIqVfHthvDEClmJDppSEvZXQyhvvQWY4wWW2mVG/4IY/Xbk
GUAVzJIb5IsbNfoNeS0Py2fjEtQHR2/vGW1O6d6jEkBO90Vtg2SHSx97XaYiI8mXsfXRkomVwsVm
cHUkyrOnarl2DNZZrQ/ZN4SFem5iR312DZ78ltsln3j0JjWLo1KoWIXIIXCVI4iFh9PAPXSCT+ka
SyT+akzvkhDr3r0gISqsLvKxk+oXG8D76o1Mn2P5IlOi4tMOn8Dvo4hNgvhjGsIlQKV57C0mpet4
CG4FjE7Ka2MVUn6clLK+Ro4EbXtyi5Yajo/2lBqCO3u0XqBd8nMXRRl3I6cnPD5pFxRjUshEQcIy
ezGwZTn23+S3MDPP2T9uuh51Z6ALSDnTaGbnQfudU/AflDx6+GVeffjcNUbS4jsFVaWdDYJ7tvn2
y9JeTYs5IGBMMwDzClqpV+fUF8IWVoU4zb3Dxy7ZDLRq/7oVMXZxbFcrlVoWBQ2mMKfBGNNFnKBz
s1nxoCcQ3+31kR2BXlucQDAJynplUZ6NihCHvTCebytPXc33gDhTMpLPoM8dmJSMbupklhtlY2Ls
Ry26Mt53hz5Rn9F/ofk83wul9t3k4hA8IIyO6afm0gFC29MNYFTiE4qLn7snzNhK4MOdz4YSdwgz
ffrnrMQmOHuM8ADbSQRp93U8bBdPfIrRqhRU1Vebj3b+5vjzh3y5X3+BuKF3D8eSmrw71yTO4nVI
nXRShB+7hpKXh2c30Iv2uZ/i1MqxfpUphyU1FtgilRWOcVT5vxDUPzpGH0TgaX1theC71/ahKzBg
4hZ4RiS9fR6T95Yjk7rpGA08bre+cZPecTb8SCyC5o0X1iSZ0/rzXhuTANLf4FW/gFdAxCsFGD8T
WBSKrwo0IF1UFZqGlwQ7DyV0yaLFbAPJY3Pjuu09sWi71uxoP1sadYecNbUMp+2za8sN06WpTU+o
HI9Mj44Y4Y7ru9Fw8HhLS8tCCwt5xFPNY5SOwcWNHNvdljrVme8tJfaQAbZxG+aRacscWLWfc9wm
1Y4lbsKLG8rSqHgL9XRnJRd6hMFKlBqB0XzuCSBGIwcGrKvXcTRaFYDL+JZ43/7lpFGfhNXbnrdl
LwNSQZKwNTPO4L0v+HVm1g3qeiMUX6ZN+A+9WS19wEr2s+vQgkdQdlFM/kBz8xsz0zzN5oeBh3VL
R+F1yN+gdGI4GgFwHtnQpfvvs3MThgUDgmDxin34+fipI0Us/cvxMQzuI+tYc6uQln9duCN85GY0
i+yHKlfh2/8HDYcHm3NLJ+04SwuzXJGSfq0c43TIsJESKl+RT1Fh/dDDNXOUUH4IZjGxEvVsPkOB
cgGG2V70B3sht6qoY64EeJ+SSR+3r+e+MaHOhmDyadjFtIbrJNKKX/w8VcRC8YMPQQjIeq5pFIUz
YQHXpVWQNJsGZUHxE2/enqUVMnrI2qNeLgf6rNmlPWKppwjoOjKCJgvAEkdQe7uaeKGyQNdeoCHy
5d4qivzXZoZX192g3hbu6/Wka7U+QnKdkpKmDaU08AJagBsgf36SKwMXH9mRunqFpVFkyW1aXjRq
8o+t8d09uxPwESrNqEQZjb3ff5kf+X/2EQQGTTxBj46vYnE7gakhyukYNzcbArcq7t5iEZX9Arij
CEwUHznmADtbBHMoF5rR0V6GCxBOxmCiSTAelC0SRGdhBg0Z6d+m+cVBC/ZTQiTyP3KX+wVnB208
ZXS6+oD4I36NBzs3tKTJ4KU6AIm27NGIMeY2yeNRcJ86DUHOil19xISCogDYjRRfLMwC0KwCjK6i
qU+PAfNaAuTmlHFsMsobCyAceoHmlV7IJW4ALFwg5jzxu647dAa8mQGVePHmVIstsluixdTGztnG
sOAZTZAM1X3wEdDkAs0dNe07Vu/ABPJsIhsQkciR5ZEHE2Q/XhLG8iUXC/Spn5bejlAH6+akCOTG
svfAEoA4pqLJGWKwryECsax9vYX8gRrcpNWRbqSB+jsjXIjb1BN/mY8uZGpwk1ij1lPNgRMODilU
jazIJru0HDzfadHcmy6vbA5CE3HXKNmnUneB+CIQC7H9RQVPossWzYPe5Q1DOeZILu1izQjyrOhh
7YWvBG23y3jt9j8wh+evMwxJfWCEjbojvFaHHLs2sY11qDXm2ADqVZcuKNR/AOQoVo63oRRUgAwZ
GyICwJXROa3jUtq9Yca+ZvBpDidIqWY5aN7ZTW3u5XkviUNL/rKbCSXvzmH0nsYiQCrjnr5lgB6A
zPBUNj1BWHYE3IYspLozIc4qXn2q7/p6OBtbmMRXusQOzuBxetXpQpiJfe6kADxj4N986+aQqeUb
a2mtDE0s74It6LyemRPkFfJshL9WRNnJcIpahczxWNCeESItbXod9AYYvNNPo+2jHefbzDR0R49d
i2z/C4wxogoDmDArSOnk7TALD6mXhq7rhgBzdDKHwRnsgKPF6vOkcnJU3XB9O88RIs+5Dq6efuCS
b5Lvlxd+B0sW2NPxDQwusLK7dIMa1hbJwnxkgVqVdWbPdK2UjgSgw8ETVlIOWhncl/oA2T+Iv8Rj
T1r+DdKPD5xTLqIFaqpN4C02k7j2E2FUtxEw/Pi0XyfLBRzH1otVE/DdI3vbbH/q1ShXGxxVkF8R
lH13Dby8S3e0g0AzOkmjkimOe1/3HPsEEr/YPxP/qDTuOO+DnxsGGFr3c22TTwJPMFAOTf4Yp9xH
rsMlvxOwsG7oBSyVbuskOX8O9wNXb5/9eaBCex56FBVpS2liMZnOkey39D76fQR2mSmopQqXWmIt
3nEz+9A/fcb/Rq2whuStsSYB3xiAP98JhJFGoay+8XvLA4A+088FOjsXwe2woLuqo95kpsFzIEE7
g7k3j39nI0U1pdUZwNhDWfVq35U2tRHXfjN7SpJBLaFPb353FSiZdK3JLnb4q69aCCNwXl4q0pmD
fpbo0O+L41CgWnAccD2OTAOz+tmX7bwwACmZLQcP+DWFvNPXhydigDhPfG9huKQhQW1mrx3+od5M
/KW9n8soR/5JdcU0i5YGnB7eiiLueCDGG5+ItHL7NS+6ji9Zwnci1NVeykk1eh70ybtnPUf7Yt/d
ndQoRfSP6hxvZA4WA4LqXqzDRCVnkmtsqRPM5shLEyBbxZJnihWYPEymhIFtmAUQGxJgrmqFwZtE
sF9AmZlkVzEnObIKVjnys4FQapxgyy+0a/Zv1GvV22M3Wc4wXcjZE/zY8RqHOy5LW8UbuZGsJT2A
tl6dHpYa2+FxBx8EUdaJmPiA1zSW8zfAcnql55FQz7YHv3rHr8LZV0tRVBhK+Z9KTroN7qxakNaP
+WLhvv6fKZLGL1fG4EyeFaCRx7Wh1LU7qxdChBlj7DwiH9QArvaE61UP+uhDCFzuI8bbyZwjUq9F
xhPZqcS+g15xNNWryeBS/54FerpyL0wcp2K7rBhNTrcdjA0CmOZ3AegXKXZEFgrB3zcLEuoVpMoc
/U8nJWKQk7aOnDCrA/crKB2GHG+jsE/CTp+qSvD1EvGQwk3xULwe/nSoSygTMGYMlB26DFdPSWRB
uRHYMCur+2cJwIWvkiMb6V52VEReutb9xTrt6MLhqNQugAzCDbmph8Wy10cQUdvDtoNND3fG4TJf
fzpyOUeSSZPCj4wDkHeIb/+qjAxKgXbSicsK5SfBY1xTwloxYcMbXS2T7mL7BEm5pf+Q2WmKY8VT
DFi5aCeq5zvrQryfnPbwpUED5LKKBSiNr8NDHb1CcE9FJkr2keIvZ05LYGZc7wujYDrlXEgNncsA
82mdpjQItzUF/2JDauYJeR6IEwVbgQGeXq0M3nCPOSm+TKbdy8fc3nr9yNWD/BWf5jwNdWJD28/w
VIrkQX87XOvwCT4S80n8NQkDPILath9X8FELfqtinPt/ER9SK1u+I18e0CVIFrHHat7vzZPcNQfI
J1jsJOZWZM+zoSseUEArcBpOMyICKwhwYbqjNJoHQnGo2/kCm7pm0mkpXHA2jAfadY/fgkioDZDS
zmAImhE50+HmjdWMYcP9rKOROSy4WeG9UsA3x6VFVBpVi76mF7hYpO1X9Y+F8DPIrckU4c1/CqWP
4LK9y3uEpI5GeDhWuICpmfyVlAb0kZgq81htBB1/Jrma34mWBSmqnajRyOZ9RHrFgEHWSL7kxfEx
aaweqveIrxHg40t4jUgs95vZp+9Kk03+H7wv25jkMUV2/9pY9+Q2k7ljV0T1kvt1I97nmw8yYbuv
KGVO/Ncd5NHpDMxswjk0EuQK9nZjI3XZYWPFgRmJZ0/Osduu1KwkkonuVV1Qh1X2onHyC+9UJH0C
48MF2JViU65v6BDw1UKzlgEsaVbY7zG+ZBIfTHREmkaGPJ1YshOus2nO3wlf1osVY5PeDBnu+8ng
1vLXszYWYKbZnbfsvmcXEXF02ofx9tjGLVFK5Yi+3KcEGFUDu55Shtgpqo+P6e6oqa47KklTgPkj
Zh05tLV2uK8eHl5ZCzmd1ANLktlh7PGb6g6Y+7dQr24MlkOTaNYQGv22qn9Go81e1jL4TWdM8wT9
xSH2Fn8uZhVUf0ACnI7IsaNRRKhnLNEsKv0olTr5+Ra2md7JuKgGu29murycVhqgwhAMVay4fj3N
hWYZTc2MAAjdoCNEtCIUGhYiYasRkSsZBFgcEL611mhBKQNQLmk9uRHfDhxDha0v1WJzihJYovBe
yBim244MPZ3a8MPGtEwoEUSRz4qT+bibuT4Ww6S+kjjvd3wOn7hDSMyPDjpX9G9wiMZpfLb7I74f
fzRkTpBm66FtvxOsAHbCFx0/hT3gHXU4rRrepMtRClzaFrdHbuouHUJt4pTci6x93YJlScPbEQP+
eaEpTcTiR6hZfIgd6GxO8tC6axM6fXuHi/Q3qGr3KQvIqw/260tvDibCCkLW4VSvl1oJ6bT4rvJo
MfLVazz/RaS7HxtJgP0XuW5bipWqS7uP/poQrFs1clKDIWsKUpzEThj87fkVXVW3aqxZwjL1LS+X
ROpcDXuiD6zMwZkY6rGrKf0HJwcVbeZZTRGp0voWw8AsVt6CaIouh7wIP3mKMvF4T6TzxDy+WqUQ
JBPQRmdyk7Krc06m9AEiTSaAmfQirU/CUgE8MAzDcP2TFkCkJZUqJw+s2KyflyVvtI64A1TtQxQD
1OvV6HuqFRWA2uOxbYjiu8DUxsq7LIS5hszoYutERSHtELjG5FQRFyp/PwMd7TjMx6DivBr9vFrt
hYHyGhpMefI/iDq1ixpPkIhGU8S0P8LgJ8uqj9B4mqGKuaMMz7W/v7XLcFj4Yw4/k9n0oCt7gC0h
feXQJXhxYGNpRPCgNtY/EU+7z1q7WxaFV4xYhVoxLcXT/+XLvnMKqKM+JaOGSfAFJU7BWfvK4l0Z
TuPFoeW9bW/bP+/p8v3Zt3EGuyF+An2OiD78sKhNznu/dQ0AIbICf9XjpsIl7XWaj2jy9hxrpviA
zmfcrOPwpg9F8tg04a15N5XRyUyWDqyqermdqQvfyFXaQ2gjT3HpdKJknEDcfPYHC4VY5tWrq4B6
rRLULKA44l7NocLdFH9CCLkt1d2XmkkzKrTxO7oS+41K+NWMcSKbEQeUpfmIeaJ+VAxO0f5EPAmv
n9YnWFvM7iF7wrECNNRivHLyEuSupfX2EKf7Bhy7IgVHt6sU+5fA/PeHLD576wh4ZiBdE3mQXVJt
8P3iwBcO4oTiXX+OAlpnvrg8JY/Uhx3cFSOAYaopM356e0qIadUcKQ9jKN8Jfd0GfngKswe1dXiL
T/rjG3/x6UhAss4iqP/gOYS2EjPjm9m0ijMpcYCJYAwGb/ZyZP5K9cCEAUo3vk6G6kQa+2yHDP+Y
S9GcV2G1xgV2XIPqLyCnxJqKt34T4f/kw/wrSQHt24Tajwlkg4piZq6COSxfVTgK9s5J6Z4aJnSs
b4wPNN3mjgaeQkQNIbFB9zIvHEkV5qXq7qjQB0IoHNC5cGbsXcW8kocyGaFFLxrPLVfGMXVgYe7A
qHthT8wls5uYkM6tuAkOFW8XcBc8nXFOCFTQeUizxrU4lg8/cm+ef9LuDvgSsQZKQ8o184wQK9VF
A1f1azKkaUtFspBdq9oLnkkzfe1lLuu0jBQoLcDhguLA2YMRVf3aK2YS02izNY2yoJRux3kF3akg
olHGwBh1a1q8fXTX7UGCsN/dVg8qZpSdhYSLMqzCMQgvO34exULM0NW0HiLDMQsnHhUdLroBOO+K
H84WPN34B2EiOg609X4AOHXtL/hAJQZWd29utqMDVNCf1mN9sPQLvHVptWPaqzoBbIp1vs1NCrcO
T2ol6BDEdbeXuA/QFhEajGcLdgRYhdA/KJPMU0gutPmaEHcefcpHQvPxvCFCw9ViAgQ5jIWrIS2L
6TR4fjpSbQz6dMYbIvmotSfszIP5ED3V1HKwQsmlA6jXldJlXhI8ZNKiZX/1h1QcJ+oiMw9UHyQ/
ceezOMEOzDf6gtYozFjKY97o12WPcLhUAwZd8+705mG0CPMLPA59RO5r2yPLXnpCEeX43RJBupcq
Vvne0ZIVyjGYuntsSV4QxwmXJc++CoqxOhZxBhBKyxwJcPvir/BPp0NnwFQMRD3+8Rsyy8mcxsLP
MC1n60ptotalP0/J1ehjK9hb9EwZ7zJtHyrN5gDE1a7gIL1vZUGm3YwV7oAJCYMTCG863251hcgs
oGpFuqXHi+cTJAxm06a7w3HW0TffDqsWNZyqpwBbaT780WOTeZq5sn4CS+1ni4SnGPqm5wGqtIZW
w/38M+G4j2xC4SedmM96c+yshDHvc1w86AFwJCImUeyLD7XHd4rm2tEMK/dAM3CAHPewasA5r0wJ
sPnsGBqbk89GrtephaM5aSPDRH4CZ3Z2DLxqx5HBUCrsI3u0X8YcFYtWtXeaYeBqKJvLQma8jCyo
8n04iFDHbhXrrUMyUm4TClr0O6DrHL5AYtf2/A68XWWf0cGtMaEMpcB5TnUEuFlxtSWrnmtC1B15
Q8dCbjGGxCugecxb3FYqIaGqPE02KwE1M40uq0Wwn4pGZ8qVlnOAmpQR15f/vydMquNXVutz9FTm
PFIj6LOQRIFW2YleD3E8P97oq87A/ttQnOP27a2SVKqeP+GDiUWiCHvkd06EzlXyTTICdx61XXJx
gFHGLiGAgM2khI24EbLxbPk/U4N/k7IRr/+WwJY6s3KGvXySy6lpTeLPy50V9dmzADTraiDBcUnZ
wHSh/ch/Zv9sq0gPh0ug7VZu77nnV6+sy2cKUsQP0GWNNxvjodaC+Lry+UdmzVrfTGlBLoKmX24x
xzArhg3Y7ufr1Hiw/QzLFfCrAq5Z30kPNWcINKhFsEfdHK3P7iKkh8rbxpUa1mSaA5gROnqmmvD3
WjpRE5fTCZ4K4valVIzI49glpfxwfk16krRkzp++fZoO3cYYqCZU9BHeLdNQvtixl1G83Uoz0xFC
29pgweLRMNgsJ7jSSV3UAGQ0BIFe3wnV1W1QsiGXEUdQHklB2ikdZuiSqJjClwtekxVqneynqwSM
MEXwVrjGiH5CQ41nm/b8vo95tmpp+XXlV045O6JjiJRqO2heN70tRWqDwny8UjF1denHcgqarrN8
1A/BJw1nXjIkJeu0xiq2pYUtt+3hKnCbpz6yw7Hswm9O0PwBtVEOBGTahsAxHKFTL4b/ZIj7CLJT
W7/JrBlf1dCsdOotSNyUq5rLlE3vAIXZ3PWU1O4SvfJDxpYI0ggOebn4AFUFP11YR7KN5QOG0VOG
ndSMCqPyJjPkIKYS5tZ2BAoQqvS78Ac0EDLaI3eyLoL/nS9cX84P4pLVIPMCHmhkQ/CWj+RvwtVW
L8rTyLe3jM+lxOUFkqSNOkAT4uxz1EVFTlAgERGmwTw4P7dHCW+paeTNHdeDHTM+HG935bk6DP7k
jKgHT+wD7ogWUKNTHbOZyKcCofPM4sfoWxEcjUl3Usti1opa/uCz+cKGh0VH9keSi3CFoaJvIRFP
GdiMS22ADBD4+1v45g4Jyk44zxYVEp8NfpRDlcfLhpG5Ag49ZkrSyHWX4rxds5COUg91aIOUubdt
5mnmmutCT2wBBObo8Ls5LSQnmsAhU49PTniBjoFQ1FezRN/W9pdi7kMpl4xaJ+HKKJhxFj9AWMC/
5xoK9Z5eUN/QhjAjB9ZEacy0Cx9g3oIoADzB9zNwface+hHjpyAVVFLMHpkUUO+IGYDPAr5Z8WdD
6cRylmC2fc4bbOhwlbQqDt3uvHpRL48X2SrjnvSO/MPSoO2MzTNsKQN/nVneZVfdwUEUbNXYKOnh
aRIKkhb9qoYJDvLBZ91xK/1vuxWlIR3dNQdoGaJ5x2w8kiFU9ESVBjhsua7eC+vt1hTVxyMK+Pqz
1TgGoUgj3fC2k78fGlA6DwvbHKWX97tckOccBhSxYkSBdk2oLek5+We04uKjVK21FtYGH/V56LAr
k2mOEkxe5HhF/TUWqBupZ+d5A1eTHvxZO7azzOooMivHNojDLJiJQdmflM7dmsErQhsZwqLwC2hq
5gPFVo8fywfvXGW8DUq2KGxxEgYZEW39MgESMzGe5+oykLPn/Y5M6qqB5l/TmX1M27R/Le3oyMIq
2/BY9HL/z3J+Vb5im5ClspviQ5eXRfR7HKVjkB88JvPQuuJovcHwGhzWkXTmgiL+HiAZQEkdgVFE
ng5xKG0tEAUkhv1Uxiv2eJunCVdmawJSB+4EII+0xV84iH9nmZyj9e7m25arVNVzcNlCF39rFmcN
t/nwOrGI3c3Izz0xPzn/MHb91Sts1ghrsBdkNUAkuxUXodFox/U9z/a6Hl5S4nKQ+BbYYshKyQ/q
dHQitsRxCR/a07FYJ3h9lV2fPjb2Zs6s/ZLsFRcD7ZLZtRMoyZeAq1H4AjSKQiZtNc351mwU/UMC
6MC+BdnUx+B564y9/v3xwNQ3Vy6FODCoUYpnowpBlNKaaSX7JZrMnGyF5BIQLw+y6zm2aa18gdBi
XQTjRCFIt5y7uIPPDHcSbH5MfgfNoh+RDDVEQVPzJwRqYvwsrh8U3jfMjJZjZtztP8s2+LTnV/Oo
9WSa2b6obYukhoz1SKVxFYBTcDnexyv2mOx6bH/2n8HEwsZdysZr6oeD4lyBerABXhPXugS3OEIk
eCvM8SNrgenl0qPUqFeDmlBapnT3WreX2uieDHbO1Seg4ALP9/itCyHVgFkaJrTvfu92NfxuaGDU
/ZovCdqgQQYBAQRRGVyZoR17UaNS3AXontQlGJ94WuK4eNe6cQQqP4fq3+WVjMKhENasijMOhgMX
GS/CJPf6v+8hpARLWVtholdVgqbgG3XrtqPf4Zq1XAnVOaJYOx5YkOiqS1Ozabr1FeVAHKDPsNHx
aQLS+RRPCidZvOjd1hvea+uXxv1KU3dpOK+6KLOCIkcXRMD9okBXpVPWlmjsADdLioIaITcGPYGk
mkYTbOVQF0RnK01bc57UR+wmvT8/Oz6iE7mmvvL3RnGW3+jSVStILvpLTsReridMTGoQ08wL5kT8
EGMtkjRCE6xvyyxUzGf9/wF08mmvdpqrcCYJXWKL/irLmZi5GA8OrCTkVUwiwSrSTIhtlu1JHj65
xPAX8nClFCDucJFC73XGdvk7IR9Ci2DBhT02u5kRuNh7T6X14yEX5/Z09ObVe+defoxGmnzvyM0S
JyhXTN4KV8yyMU3CxEtM+as6VY9U97vT1KuxRAzzi4NzpcRnCOylhJtW4+iVCZKrd91J8DXvdP6+
sHlwADCvoWCt471Lp41QQwK3r7EuR/QaF8InXiM6ZDVb35w839xEYmDXx3tVXqcO3vfiiwHU1iA8
LgqzOrGLgaAzZLgTOv7XETtjV1J/1qVFWZuUjOQ9vzUgPRXsV/qmDVJ5DXb5GTiabfi02Rjc7wvf
Y03xy0niOUSQwmhT6q6YnO7HoNK33kcEQNBOlqq03HABqtye5m2pS2u0wjsot0UXujB5b17C01NC
7dCWF/ZTHPXIfIR9WhApMWdwdSXyPLPeAJqFJKiytkHQ3y+NZwaVf05/5fsxMuG9El7IkBfOeT9G
V6xtUWrGzwSxZpfnyJ3ES3uQOn+MzDRgPrbSnpzCSVQ8PGNTBxzoqR7LsqpyMza3wknBubaBffBZ
ukAHfvHW8pSZRsrkx09i+1PZTv3A8kcSxj0z8mPlyS5CvzadWW/JXaMiQXB5pRFYA9W2Mcm3uQBR
gfKEgdLDh509OQUxwhCcyXXUkvRGPu5nUboIph/3D909pFaiu1D4hHnBE/1AWHP3fpAzR1a09bKi
dINfRENrG2UYwRsizwbM6DqOWL5J7T2m4XXvYvfUcvMsoSGUqWKT/6TSh35LXsdFl3d6qpgQxGYD
n/DaDHOMJjb9MunNrKPYDFhsZdwuoGVAn1+euJoQ2HSE6dRx9+gF7x9x74HCuWOhz28oOTmwvv44
BQMWVIzXdTlVZLFemW63sCE94YgdJVd7A0K8BxlpadmyFvZ3iUYDWf0JNkKCYVHJET3gAU/BRqSg
06kCT7yFGVwr9jldXpfFFEukpeZmDydOqFx+tG/SKF8jWgncQgQWUd+Yi3jC+KsewYFFIRKmcgmq
dWNJhGdvDXquR9X03v1FHU8mGYU5OjrdxhTjewyKrLbN18WY/q0eyRTsx3N3mc7gJd4YVWZZe9o0
mPlIVpTk2gSA5H8JcJe1K+O7Bi0/551+zOE6tacGQDT/ZvyB24F7m5eNhQc8NGBkNDuGm7Fv5GKg
ssaz9ego6sRovfth+tg3qxf4QdhBzdoRbG3BWSGkUgRni87UmIb3brsfQkcT1qr9f7EZqqerzqym
K3uoEihrJRBc7+8LIsaH/yuAqDx5U8R4cwBtrMR5OxdR5g2ykFAVPv4zmcdMCXJzmYdE2TL8ZbUo
XEr+DeOujqTiQh5bBd66mrAjVeYHHcCDXQhnu+o25rfI+VvjZXO1l9zwW7M8AQrzjZE871NhHI0z
Jz9igGRDNRce+JEnmU+KeA0B5PlSDIWnUrjIrTwo/Wm3Y/Tio7rWFXmfMu58nyiHkOZlpgFZVQ4A
5i15YH1fEsLzb3pVXd8NGXaw60jRL/ip/z7DLn62dlwiiO+4ddX+2ReTUuQhY10qsxwZJ7oeJ41d
SwrMeYurHDnPeKAScYKpgebPmzO8TGcwnwrrpGmtOKdwRxgtFnb4Ls7P1rpVrxYo5N1G+xw9wVgc
oeqZNg9sLXKbr+mO+JN1y+MET+1XNrn+kuvIpa6U67WEEOeRa6pUXxJmjI4ByhNqFOF0XTQ4+2NO
gt6ESTVu7OulFILdmJ5Kt7aTRmnBaVWDzvvPN3SQ+cu9r6yFQpYVL+oCxRndeESbqFSg7EsYuzzL
6mT9ONZXbE6JcBtyDWfpb7bYWY4QlkgF5nlk32AnbGPT1hX+8iaqw6nzVOdTHDMXBgFlnC+cBJjM
Hc6SPtZvXLVqRTuxNuOc0W+tinML1rAIaz0pkjyS/2L2vBR/xej9fcVYP7b8SacsG4VLwndCZfjl
HuKQvYzUudkiXKU2V40o7Upu27elGkABd+1GF60o8obVs2rDIAF32JUZ/SAGaKln/E9Xf3QCHhKv
c9bQoSJi6T+poMhfqryk9h29tD39wq3V6Qox23sgD78ZTNcb2KGp9dWnboN2MTYFffaqoB/sRtDt
AhX7MTmuFSRzIHu5O7BLTCSCqqXw9eg0DWE4pWVi/6oAGP9hoOeulIzFnENKkUqGeuIa/Z7Pd3V8
EazGJOhQu54/q5JwT5adKxY9gXJmvyjxqaZOdGjxhH76Ts5tT19aZ8yMbcXfgOotEer0YV72zp+u
O/YEunDmya6aACs6nhESDfs8PsNxOkm0HfS/SZ+P41PYumSN/t08EaSllZPfkzN2g5Y9Lder2g/3
SoqCv9/ltOM6AvEmz5MBfRkvuCFE971v3nLxtet9o2Db6JNSnMOxrT54n1o2aQNgPZBwljNrkF47
L48Ax5CXFWiH2GRFVX+vLTmpaVWeX5CpW90Vmkik+p9oHsK1QJCq2SyDOg60lK3vH91LoMk1Q+bq
91tFVjLD7XRwJ+pEDRyCPT6tpkyK11sWM/B9qkJGslCmkQyRY7O1ZZav5OXoFNj94TJbC+Vt8jSa
/BQu71m9ZU4Ebal12B3/bhKCvnTlI1Bufy1QQFn6QjmZKOYW6QsKA8RjzjvmM5+VbHeM761aSHCE
bxtpHZPFRwLBpnLLOCdTayl6phqN2zAC4eAy4+NJN74wn3y07PExtz6PDqipSeKAO4N3O6nwsZwQ
TX18LscCSjcatqpTE1jj9dZIOFRVlA3hPWmCU9NUWf1SJZMbT8ksbHL+P5BZtcWQxZgyDMxEHCct
ojYR6AyQSxvXFzzWUr1duShgzbZWgp9Ytzks3kvu8mnB9kyE+HUIZcVhguEjlPorniVC+ufhK38a
7BvO/Kp9uJS1JE1C/5MfVwBIdaODtgqRvjcOD7SHTBKUYygb9cC9mVp+sTrvbpZg5CNN6+O6zrzP
YdfgwpW1KiOl2q6vaXlOJ7zpptibyM4fqLDJaTN+OEsPZTCBr/GtygtsrrgsJOoBrRyB+ilI9psM
itZ7PQw9ksjWybVBDabmkUJGWP0iv7qDVk3GboMe2XoW1+jEdHuTubZ8Yitq0Rh2TuVsxUA4/y3D
TOp0GOb1CePxiGVrEBIaOgGkI4LY4fHsLewoMHN/Ohbg9ODTUrfTRHLb9JwoE+Mt1CJ32cKgC5UH
LsefMPRkJ3RtgXazzutKwj4TCucPWSNnZJ1StHgCvVdhfb7h+nA5JunKlnKcXPXcZqPIY/LnMkJD
isPLUV6+q+ohfnZgWhxm4twAvwoIw1Zi4WJ9BIgg1X1Jdd5toYH8akywyxXi3ThyXPlSh1DEoCfV
iw3uW3tWAYs7FlOwQkW+9c0/EnedwC56bGljmJx6sl4x6NRGAy4uyF8el58GAv9Lv7QmJIbxnrsq
9eNuGM7pjoxQZ3u6O/YzikPglyBV7+eGqSABDH2ECN8ltny3E0r+Rhhxohir1qI6Qr0xMUgIzkE7
wOEqx9v+eFEPr1XJ4RHgvpM0mcY5H/ROJYQh5i0U46m7ghKyebE7qNKR6HjR7EQ/Wq/D1FwN2byc
ZCAs6jqybZFUH9J+kUaRFw4xCzUQ+73+NuSxP8ECDGHkWNNGK2TDYQUPuTtqE1eKNp4rCDhbHPJp
NGI7EuajjkHAy4zThRlUv7l066GFyAMNHpOuubkC2szdIH26Zu4tl8XrP8oZ6mRb7kWjd/LQoT+h
7yfqq9CCBb1dbvRtBJovYka9D9gxu2YJlTSGg0mfZo7z973uOQVuYoMdm/Q3SqzTmNkLRuiQXoUb
WzGLxUvM9ymfPPlp/yCEiUMwBEigyrvPedpSSzVqmbwlboVGBQGKVYCFaLDmoUEjDe71q+mryZHX
/7GYY3SFHl/bhaX+scZ/A97/97YrGib5ed44wd8AK9ZK+TRdyocZXOrQd/82FGmc2/qKW5n6Cb7D
+v+yAWmnJ0jYOY2jCUWkLOu6m5lkJK8HR9a79C7aAzD3hC4bt0tO0wY3QFAW3daplN66IH2EXAhR
L2ZtZLd4zjS5JnC9pZL01Hqxz5GeSJutWOGhKRzoZVICUGHL7iq6XUv1+WJQ+8B1rUgYlzN9/w20
/RMtwfl4UFgoMoJ1oFtrfMLjALe6QuI9Ko3eKAtttFFfSnMVkaRM3rimpEOlCqmZ+C+kbpD4+LzC
0tCHCZjXZZXTk5VBLoLD/G5MWXnMDHtMVciJhu9726JkeimjlYlPcOOGrkJSoYBG+/BrbMGb2x/K
ssBiir8N/E93T8AMLuD+j/bLM4Xo5FVlqDUatJ6cWgyACNhnSU35UhR2Hs7Gh6PBijmEOPJ5fvAC
vwwE+JAmt/5jt75ycPV0H0H0PYAtlyfHNX2d/Lplni2BUqD2CVTVH8V9vcmA5ulf5PAZ/HRFNQHQ
JLnp764dcoHvv/glTWWZI3JYbs3K56aCJiZJglxMeLX0MzaSA9HkzwgojDc4kTRMSvU3mZ3//Exg
r+ZyDAAcHH+RxGO3rcA6Fx/riv9bvaZfEyE6ngHRTGlgvSssNY3pRvthi9cnGvTWoBk0bTNIC/Pi
UXTjpOLCFYMufuXWWPdqGM707s3+wMklK3MKvFpsunnbkTDBFOlvcA43zWqC9bap97+mCB5ou7du
oBNzESxr6sQkrr83lPhJkD83DMVqtCpHFxMWrChpkD5jT0Eps5+QHLGJypvkTSMHzTjPI8PwmP7/
aRNA7KnzbXBtvZqcknyQkOU2Gj7zeTCLSQXM6Ti1+A3n7n9TBHrcnL4uqBHeh8QkayXZXYspZaim
gfxTYaZhK4wfGcakyDpMe4eaOylW9NY5TgxJixytmWwDZfYthCe6iN9KHPCY10W9ovVbXyFZzNJf
rYS3wQtELNtOBDPAAvC42QTXvmyU/7IiaZlnRlann3vDT2NheGD9wPHzsFVZo0GVR0gQYEp/WFZ8
+jXvjRVkm+IEByZ7C+XESlTRUlxpAeOJFNVG+bQ+PzNwuEPen5gcLw6rYZ12sFkr27NAEJVgJj/i
fm2Ikm762kRJorFWd5S9WqRU/Mx8t2QgzcgkTMyXHhplFtMGjtBzMAaN6/gHfSepr6JNBFbcmgql
rxXHooynsE7iLRsWS6TuYwT3cjDatc8WE1O/TnKskV+grb6+NQSqohpz8LVpgQ81yoK36qbTkNuM
4RIq93uGbimV6v1AgjJjjDqgPFKpoC0zOM9dnKtwQwo2RlyR+WG8O/QBJ81yVzOR3Gl1m8t9rbZO
jdc2kylCUD7oIDlRt4dj2oCGydjiK7gkVaSFb9fdjyrDWxxkkuW6DzfTmHz47+bDx8l18vFm5GZS
GYe7YFNRAPN4hgJohuQ8qSo9KmrCIA8Fn5VFUKErvLG1AyPaj6UxHQtGd5Smz1P5xIk4IVi53RJE
JTMLbOvib9FUgOwIQpXDTUaDfO0nIGTrqj/TXUlRXmzwtlQVigNZD7HmsakzPgUPWuhjJFCkVZSx
02eed9+z5Pl+KH2V7nl7iwNd3zgl4yxwvxwkGh4ZLf4jXBhjz7cI8pcOvVsqpc28LiHtVv3tXboL
dIF7vCnsPlC2Mzy0MhEZ1cZSlh3u5tXTSP3uPnfHs161e00DZ6uRZMxOfH3+GpDvrSemuCu2xop0
YBcK2LhhxVZv+ZyCTXopeJyFcKLe1qWZ+10jxH9uIiXpKy9K5qNkPdkPpzuuTJrlNjrHwRDEu9b3
L1KA9Kobzg8rhKqgYNpU9gBTyPCTdOAn/81mP3HhrD4tYbu93wbgz7JDD+2Xroydez89jFT3JXWG
lZ6XgKfdZ+0zHl8yA1XRxRySXP5D0rduNvLT6RyOdpzRR3j+M13m3422F1Ixzg3mtaNbBDh5Egw8
1LT6TA33uHVdkJrVAHvPRljNov+Ny5Jxg/rkZbnr1mERvuXQWXhGjJo4KZcbubPD0Q0kqGp+4ga1
Zm2ZyV4qS8ChogVLSObxnY+yeecS/JBR3a0Id3+16FycSScRqxm4d63MC5ZhFxaGCNDbzh+rISKu
wXatai2IOSWM0cSaQ1Upr2ywdh0oGwu6WqbEA/UADTmsJZF7gwW0qXH9GNfhSTfbJPBdNWFI7bc9
FP46vNNdRwQjAZT9fZEp5HYV9dBaVBpsMQXtP6rqf4gamFIcf9RZFU6pktiaMVyAyXG/ob6euWGA
r+Ol5Xyblb5W+35nVD3FiCMLGg6oaiX2CZ4/rctg3hzsZXmjj3Q5njHw1e2vLe8xtCXEMk0RQcMK
wNn9wztvZZcCIouSifrqGUkjZkg+nMotSM8qIE7flUsgFYUil5g8FSSASrDOpQPLx82FEJdyAXwy
/MTLXelS2lDD4gk5Kl3hstRNtSYZwgTPbhbVmiywEY19fSUyFfHGU/O9eaJl+4F5Sa1FeHxoPF7R
wbevztmFvt0pAFVAIgxCRFHwl1ZW1Cvz0yziTZ4H0TBP2ua/VUuH+aBKs/s5fQ009rr77ImcyO+p
7sTRrGChiaZwbCq1rSIAYRqmuqPYec3c28YgWJy5Y3TkEKHcm7ybuXnnJcNo0dJMLKVJPpPI1/1Q
YBTX7xPRGBprTHJBS3SijPSfHag5Ux71nobmDxxY99BfhP7eQNHxYVMY2QwU3rMaiui0lknfTqNP
Vi/ZhWRpFdgrryqXFbvN3DV+wLHm3dBw0hZ3MdR+z8gt2TulArOgqyZXEjxZJ4BZsivkd8P2jQfI
oIAnRx34LWM3daTWKgfY4/4O8F/dZkzE/AeJ0s+0+uLJiF8kFsQ1wFUDpJSvWeXqFR4yIaOsyNTU
8QC0aW7OF340I4/XW2bbwTwfsbZaGcOiRYvdXsY1ErkB4IMfNubB8/YjWrKOUW7C4CFCnkENsjJl
e/S03NX1tDu+31k1weT6Jnw9g3nrxeRPWVJ9xKlBFDl6QUwkyOaU8RQ/qmlqlrrzovZRnS72FYTZ
XnIqGtTBs2kAUHX+gTK1U/0IISbVY+CTcsvVWIUmfP2VMnlUng19cWVuw/GQeK9wNrinW+MF4XUn
LkCpr395yoJzWsLlzmUeaVdvVY0uwK5YgcRc4pycDGhbsa0xrBpTbFaKIdw7v48RGgZGPlUnIB0l
g25cAzCMWd+pABCxlRPYzm/a71q1owALu1z83iogssWShK54KN8HhOBxorzfEAH6JJ/BaQW9hL5q
V+ucXa8aIOmggyqy9y3MFDQ9tDbEu/Hx7VjHiFOgdMksG1JT0LFrhWGZHZ3etdTdz8h7wCW34fV1
Ppx7JERchvxhSZlSrDlgHy/+r8BuEMR0gOH3BLRAiG7RaDPt9PaKLlqhexl2kkKXgVWICwIK9DTM
wuDQOQf/SqX86vdXPxMb+8/XDWmOk4+S7U0DnWwpbyPys0T+36ZrTrES4DwfguWPcv0hg/slH+Bc
LXSPmstjFVhSH46RBsUqk36GS/wixkXo3kbwfxSzucwhrDQHmPMRRa8QNBN7ge1vy/ipbtkvHSqx
S6Sh/BIUWgIF3Q5Q6U04O0QNp3kVq1VlmE8i0rINMWrZqshN9lRI0e5vFohSsXmD0V92ytiGoomO
kza1tVb3lhSuQ4bkw3ZHYOB6ay6VDDiYzrzFFUIMlMDxdvZ4JByuOWZ0/eCu+FhBLpF4hSPhuTft
dIZrBVycC0Ot4Dyz/SLE/IXk0nO/CnldEUj0zpZBECbR09PiV4+ktl+lClXoT30uG1LOBqpMg6kC
4nZb0jTwy/oYHqyDsWI4qk/fV9EaSmky0JkL2kM33ZlkDE6t5ybPfGmEPmwKqwazXUHHlmVUcxXt
j9Z+C3jCTuiyIdpSv38IMiTc6Mby0XGlTkkRfWNCxwlRPECKhp93PGrBRgWKJ+lwPumH/RATWnEw
K+GT32N1iN/jaKgfeRlC8VMIrGYM3wYwG0p3gz0sS7JtbHyolFpQhx+XtqcoCQ1sBtP9NqAcchMn
zquDB1Gouxw9SI82skH7/FEn0CzJT0G76VwWpcdIHbxozIT2bi6YmCLFykw8E5NEayHaIpNMWj2I
7j7VwDGjD36ZGtBQi/59ep+Hi+E3sKQ2XbKAdaNvXA1ZLQHIJjdjJ7CvuirpP9545BFoUZK/p756
OD6rG0niISpMnjHZOVqyWqL+emR9sTtiKofAo4+Qy0WdmD3u81A0UxTyXawAxFKjQxE+29uwT3ty
+o+z8wZNeHjTx5ZGKQdpjutZImD7szTMN/Sr/GlpaCtEG4IVUbpraEB4vXYtChCc/MHKzNhAuqws
D/co9BYkbbouQn28CqQ8eW+F/KBVglmyxLoHpuZe7wRxpDdHwdLVl1Hctt4kRyjAd6tOTYz6OTSR
5Zcj/V2ZRRC6bqqg6b18elNCBfjTM6+A8COFVIcE895G579GXRV/zr4NnFdJGUqN6DBCcbibaaV9
eZrJHTMaYCxe1751iniUCAqiTGBhq3T7hSJvL+WCft3R4mCY+VprLk85700OxKoY3vng2maPfLVY
gxJDvMNCh5M1FRi1F6sD56+XSPApmXmsQ6rIywaXn2xVu35xjuMLqJGx3Oy7UJ+mOgYThJJVgGlm
NTVmOxJvu2mn8j+ea8a86nz4Hy1brntyMLxevw3/pE3gvDZcEYDVzU9yT5/OI1ahPhd24T7/tiBN
2AdQLQc9hulcOwW3QojjQp2JFesc7R4nD2yKSqWHoiZOxmgdGlPAC1U+MkHPtCtwiBibaG4mBFWK
c0aWOMMbRTwY6oWC2hiSk5KghVRdZbcDIrsASGTWK/UzUD0xppHLzfCITspND0EXs8ZtdLwrgvA8
pPOC0VDsDdn3n/G+EpmBySe6DS0aFmlYV5cYIkR0fjTBZWUCZIPwgsuPMMBHpu5nlSgrzdkZU0/H
NyI6HhzJLaSwrZGWTtRkgswZmbLfeKvbaUPqEzu1z72AjOaeBaEn6zgwUoIEW9XSdVPCrERpJWhG
yWXVUbQres3/r8dIycHqXgNwrP67b7Ip/BeG79/NfLZYba43ZR/JZskaC8JCnI1+c2DZPT4YicLz
9Ulm27yrxIJSz0f7vPooKuKMMAhbIIEhnl3wuC7D3BNcGxwStcWEodSsKJRbsMZ7Zh67/B862yfY
MAaYZ7l45dJ6bzguyaSVJ81dtzHHYR/1P4qcb7BcplB/ToEXtxlUWygjjwPbEH+6FdaaOs8JGsDc
HO9qh6GGc80YbSEtgdlEwlN1LY07dNmmKwTNbWR06g4YzmxyM1W19kaes7lfzB2a8Uxix7hg2qAX
zhigBU8wWrp93BZZma+/12yqzpAHOvIA2igdrJXWgwREjgTc1M4qLdiHR1mwr7ZkiBUGVYS/XEnV
9LqjYmsc2KOXduL3m7+8EdanwcEh+MOSFW8gX30Iyd/IdJcqw2y8IDbqb4BKxlr/P5iFuJ7ECr94
u0AvCrIW9xZn69Yz73yViPn2jqU+WP5RB++zbPKN5Iu7zQ0+7lG2mKof6KIQQ0JLARXaJBb095Wd
ldp+Fh12v8bhnON0SRM/l883pGPcm14t8xOlx5VP1h6ln3Z5af2HqpmfFaDQkLbaRxETY519BqFl
Nf4nyp+lqUMOrpQi5A/N8aOZXZ76VjFA0Lrb0t6ViwW1W3iKYsnxs3DHQor87VVI/H95zupEDcvK
Bm2TsnImc20Q/VTjt1F5KWMd3ruQMLakCtm+WwVgd1Lr4m2nC1DOCN3Cv2UDiEUJe//SrDCLw10H
7Hfks75mnsamE9okSbS2a1/J6VfYzQlY/TFt85QCdji8J23+ARiP5/zQaF+YfjT08BxVTZKRwBIg
/ionnd5z7qs7lHXxweTSi8gdhoeiFoyoM9r+IaH37uCfqqXPUJQrhzWcY0CeRylKO4haDBF6yFKc
WdPfJoiJhsrTd3CuNxcGP+m1QoAhe0Wk0dNiRhg/NWEuzurtqY3zYIbaX0ZZnaYtcDIyMPlBFj8F
d7R/MWCvuEJZlRe0XrjXz7cVnojS3PJCmKgqAqMFHhpoLNj5iGBhlmQYk1PSLdkJ0MA7lXKrfhNN
Y+buzx4zjjUsf0NqgBJfPMqvf8JaHPB6ql+TMFgQw2P7ixIFcSPT86aIO77ZY9tcQar7K4a1xSuM
1XR9ZRr1kn9rKL7qFaZpWa30lmLVZczI7sMOVfQYugWEP4Ks5DnPXD/0iKfUg/wl7a9osF4OEjX4
hVMFZeuaNB1niy0l1fgNdHvbzrxly+qWWQ9dQxfsJAZF4AUSYdoZFvde+ZYkPKYOxwFmwalCSTFl
/CDJAlf7eRXEcXpl8ole7B0s0p++qeMPu5l31hbUxGc/IqzFqNzm3NZ0qSQp45Pya9WBmqi9pC+b
2UcqWU8cWKim3Ault3Mt6qA3GFdeNX9Z8C1XrvpgvICh6MCK3jnaXbi069sVbpHEA1LQMCS9uBZB
y4WnV8jRB9WGaJy4or0mScz/iWGhsY2+o5T3vAJyRU5GldaTy2hqVr80qhvTo54riIw3oL0xmkxj
HYW+W9bedwplWBKuOcgL/1CQ60Aj/ih28ooK4lL2PGb5f8o51R3rqbL2MbkuszCwbFSwaQJNWK+q
WnXWcP6haqdV6xwhgGJxfdZzj6/Mrg23ECN2FUyQaqcZ6nGKWCI7fwXT/vBzlP+4X0bktcaWEoj3
oKxreYSQBbV7TS1k88t8KUaAgLn+Xz0Mc2yVvssqoTO3oaQNU0S/eGN1yoM5t5ECbXCmogsYccvz
3H5HeHPlTlpPgb+rP40eVLTkF5bg/aFkidzTACq+GmVw4Nb72RtPtOeK+r2bVWe2z7tKB0du9VwR
KXla6Nm9QjingqjJPRDicH6riLf5w9Me4rILfuDJAK31EwZ5+iAXR/lLV9eyN0QUOx8Tzp9oZHnp
Thr71XxgzeVDomCvJ/QTuR7PO2ZVO9aUl1I8HUYJCrWF7AHEKFUwEvpv6U1+ByZ+9n64u8SGH9Ri
V1HXWW7f7moG7DAMi5AS/t5PFcsgGAJFENngSrp4donsHuGv9oGEuESAPaAX2wNGJH5BuHQnN3fY
Uf1zw0PLOJywJhX1wCJU9G1xCmeKU9PtY5RmfOwCDTNn9L4uZa++rg0fbjG+ia65uZQN7CLtxsqO
0a7vlRfiNe3gOCwWmb8rJYYT7HHgFIHq1k4OPSkEqicvyzIcN8uRGt8KZyWD7iTgxZWx0AScnCh4
NK9+OGZqQTfZCywrHUwG8AvJNcoTkE4aoWOUUb9NUy+i1KwQR0/zjLoNag9iXcIzEBA4LQqaN0UG
AkKagHnKdi7uWqg9uBugK/TkAhXwfoOpuyCI4kvW8AXolxWgfsCJzqDBBSNcqHhcQ8sEwGrjMmmR
urOnwdMb0TdmQRFpP61WvvAhsnoM5vcIrxyHYUzCHhmPQ2Vs3LR+n8B9LlJcXmAFraJ8rpK8IKQt
zUHUywVHb7f8g6YwSR2B1iLH/FKje7nqFFLTMuR7Wsd2TYwF8TEEwOgWLSKVaumaBhIQ9dhbvUD4
/2Y/7JCTZWuFjezHAaaDXTRGcBiyEdbHwzb3upN8ZIF55zPfG7qPg3mAhC6kxWAGWpao4GibhBmu
ccb3Wh7G2YoHsHMYzEX0p9gpT6UCuleiT565TROIH+cWvsHyXE9lymS0yMLx81RHxwY2xLKXPlOz
N1pPYkdfwbxAmL17GCYgRj1Bz/9rZgFA4itrxdjp+u3oLkzP8RIPAOtaPgaVj6vccyiK1K8IuWkI
zEpZ5iw8ki/Y5QawbZ249+oW/nx/s72RWtGir0A27Ck5YYywMetDnwBo9e0SKujBymO+HLyYsSWl
G6HEA6JFYtJy/jxiSmmPN0sOat2STd2OmCjKdFYzpp2FuCAIjSZbJ9I8a0BNHrzNFuRvC+y9BMuj
e59kinmzrnkcIMM0cig9o6E/QhUfSoBFS1KRhvKrRPDW3glBHY8BMNc7g7rx8CkgcXM0P7kukm3g
/+W7C/rB1qsSdhIt82i/JqPHliXlDRB7raNfxLN6mwLuL0cjrZ66s+Tn43LKPcmIWM/9Z9XEeyTk
LnXKUmcuoPGXxAxIbr4fMfuqokkXAnxN96q3xkDDNSA6J+kXq9WCkqqBZAyL71FDlYGkBzWZIN9b
PgmWyAHeQt1wXTfOxZqC8A00hevUtLcj9hFb2UlcT6bZwzqYMeQ/cXZpUIFuw+biIglSLIkzi7FO
V96dgT5AgR+zdwU3273/RyDnqPYEp0PIa+3kN/iHiXJFES3+Sk1D/ZbPcPRcwWPBPHW6tLBlIdJ2
zOFJjInCiCfA6J1A6tZED3P2ZYH67huUIVT38KFxMw3kgiVGFhi0ekhLOrYoLOfIzntPNfYwI4O6
W94+cMJCtPwUCye96mmhUvDS4DYGrCfk51l9JToUZTlkxcqNplDmdz4xv5z926O0DEd2utIaAAeK
YwVPCr67fuINP2h3Zp7z///4+BXfJxlR9Y4RMo+kVMl2i30gjq4kFUqVCRgs/i0qpesH2OxsTEmg
2ilHPKh4d0EoejI/optKTXOKFtDswyfnH6XRuZH/SFONCN5PMMxPONDjClfuu4NnspN5L5tAAMRA
ZuhjU107jiTwzChNI07n/N9udMKIwWeUcCIqNcIBKyK7rs3SCwPyBWB8l9iDyXOi8awU191KkS17
UlygNcWP6oBIFHLzp5mNZN5iTho/OucIuRW7V7qXocr1ud/n53ELK7R4qs2/eQoj0g8ijkmTO0oA
EsGr4yiX5Ng+CAkVAZBF7HtnGGxX2+/31nHcsp53vQ+RvlpvINVIv/mvPFEvpwbVgKP/cXzNCovA
OzW1rbew4n3VdFJ+epcxy1pmy5Ydrc50p9UFHz+uZ1rQsPEVMm4cFDFVcSjTCpf8oiT0GH4lC1v7
dIWESMnP47BtCksTvA0Xv305tlzSwyx5JAakipdIhUWdsy3NEIfL9yhm6pjD+uSkWq90+vXHFoSX
iKlAMdWMI1/6X3YBdIryvvMPce11Y2f7Q0yAqYJKGCO0MWMsgMIDyxMWh14U4KaxMr2CFv3eKFmw
NcWB3ld8Bo4uUoG/lnR1pFOoiPSFcFZ8JlkY6+w32t/qGITzJH5OOLZk9fH+FGIrU9zt93CclXqc
a+73FMtpUD7hetmF7GLlF18ioiUY94GCaghf8QdplyabPd7NjrmUd0xE+uklWgXtZY9pebn9gH32
LObpFGanpCu82bYYjJzpPX37cfShz4NEfPWP14/EgaJ4t+QWdocdWL/GqchH6Y89PgnBQYUjSIPI
cBY3KLUtcYNGxg905y7DdnksPbLwVj4KuPg7MzkthQeWtUmB2noRRt6/js546WVjG4QGybELN5ND
xwSyUhV2/L9liMbEXKPmXXVj+aDGxsjAoXWAwMS2hwe91t3VGDWyzLoyU5PUS43zI3vNYyMzYneS
XQzKy1njrEkbhUxXI6A1aIo2CH/WALxUnfuyuQ7zkWZA4Fj0ZODle2n2Xb/nsUkOjz3SIOym+krq
GtD4NAHrvZQ/aVIu8J+I+JSjhGqddtHTZygREXIDFzt3BC/yPx9aDhX8p1vJnhJhXMfepBCWYxbm
9sxJgRXUuFONq0RDfNbU4IliCHRzuDdTZhuP+MflQqfgbCZXofAHW22foflDDMKoQNwgnUnk4Oxu
5x7DpWx0okL17Uex0wFqtYZV3cJaG+N4x5Cud08OqndMpcGrmUztI4675Y18Z2K1yaNVX+2wMJvd
jPsPsLbNlJ5WdzXuIaoWzF4BHsJjbpqLqg6Pwb63ZzB4uXppGVWbAEliZIfGwc4lKiFSUSLOyaL5
k9t95s4uNkA6BPjPVaBsALuRTCV9an6Hyc59qEqkuQNYYdz8SSUbI3b4Brid/PNV32xXYHpj7Xs8
7lDr0g4mbD0hOY6OHuDDnb+zRI1sACiaG1YT1kkYX4PzL12sEgxNnwe9qln+LQ59cSAPOIIi6UMk
lhy4+ZNjG/+De9wtYDeKR3z1wZFmaMQUS5Q1qc8MNm+/1jMQfqd4VP8Mtn3KUpQZjzv7AYOcyWT+
BHEK0RJImG2Zm4MeIIJvOUTtA3ZgfEmLx2WqAsceve6uAzatZ7mMkG5cULYukkJZ1g1VyLeTmdyj
MjVp4ygTmznpbSKy60lyxR/Z6qjW2Hh4s3IofaXrdXnpDw1GVflfmBpbNz8qorhQgoHPSk4xDYpZ
40DUITcp8iHzYLEh3x9NZDeTVCQ0W8CLdSLB31hYvBhmp+FuAL8ZhZe95opjOX+R262to0Ow5Skt
BdXlc4uwLfnIH44qXnGo2/MMHx06OoiRBKwbHPis/tKiHDVzQBnnttc36QhRaoQSY1knI6zG3fXo
JaNgCtDcj2Kw+KmPsnraSvQb3WVJxpV/EyBt/UwV/TJE1N97d3jVQXqRwGTRuZY/zEfrjtatbeG8
bSDQPwAQmH0pWJRwPIT7ZHPq9toZRBqXM43McrgekkjDmwYGeQy8f3nY1Nsmawg+TJawYa8EQ4em
X2nTrccRN7LHeIGSFzc4nywv02vJPo9CmZ/QBuSz1x441cQOMY6fEGatPq6sTwXrnkRzzuWMM8Mn
OBti4FXL+dXcd3Gh3PzVrK8oh4DL5zStSCrSAkCw9Qy/1NeoU9sofB/YNrq+XeruQ8KLPuPwQXZM
0BvJsKLpuTgRFby6W2cLcTu+XL0mZVFTLrcu7JnsvzuA7EsZQ2WmFCF4qkNgCEDQoKWF9d7/bm8D
EyQnZxP3G/ZawLI+yOIBs4H8WB7LmZ3IqoB8JhQd1MewKHLk+GRTVbIGgOuYF7oNeuG9K8ZxC8hb
aZwc7r3czgUQFBFeQ46PlId5IoUTquUEebXt9N+cE3NxiyAwuMHFJ7OOzaQroHiLmhZOf6ZEwy2f
kXzeaBnJ8zWjhzRXrXajajqOafx+wI/0HXFQd50VMOnszFORLq0/eNJ6ROnXMzD7jl8Y+eVFth7U
9lQWaVsQ6/+YNGgR60iJ2pWOr5Eo+sgpxWkzYAm8WVaRasLIhnJr3ssh0Y/M176lnhWPXPe1Z/vt
/chbOwGp//1HmaREgtH9PoroZUpU+sAK55mGwyI5OXWVbJVTleB48UPG+QMErwP9kv+B0+kzJt7M
Jrs7pF/xN8hrVC7dX9Dh3ICHNmyjyBU3URCDd8Mv+gnnPLy8Vj1KK0WRnPQ3oeL/CLPSX9o/51bB
oB3AU9+2DXT57m5++ow2KCNE7pjb65YCDwH9Byey4lVW9n4wHY3jDtsVeTI8Us3Uh/e0ClqpmOfN
A5/2KM/ehI+LkH3fTOVl1FbLIgj1tpZf5fdQv/LRx26a9G066z4kU4CmggIucJLiAiIp75JdYgP/
HKkGIW6FJKPhQZ3Mj0K71DlVRujA8Sj+lJ8G686HL2wZ9pzM0LVyqpXh7wCoZ6Uh68d0IorJCvu1
iBGsnM0xTEJ/5aasB+FnJSV4T9TVDaDZ3Jrl66ECQcXDGgs4m16yE9Un8S5WWPrtDZjlSimWKTgJ
RbcyFlYI9lIK12HVFcxy4foIdnvNu4ZiZyRM+u/c+lwx4sduZCx9vF9Y8fQajK1nei8/w2t+T5yh
Es1N4WKe70V6HXJSIWmYHHSXpM1RMGo6HFYtGsAvOJjbDtySPRU8aoA6YU91NQ1fHEUb3/uY8Nuw
FCehEurS+qKs6vLC2vjJ1sA2VHOWaGy5sPsIpT5NpAPz3ntzqhlnd6vvZztfmeNKygME47IiBMiP
mYgHjhnqgd7gP9HUexndCYWie6RtH3SOpA4uc0Ao6d96swnTb64XNvpJN9H4LyWTj+d3ASo+qvtX
Nbzc1DfR5NA0l8SHj2Z7cT5ZoZHnCy5ii/ooTiZ2S8KmeIACm5kUZ8IApJFgo3wmyyARxbFGIQ8c
YnXcBoWNFyn4+0h1c9oqf//HiXDmwQIkGWK3N0tYPafh8C/oaVrR9uBv/IZvX9GdwC6hdNYY3sUR
AWeZcOsWAOsVlLtxrUWFLYq60StORVnIqAjOeHEG+NeVUqyXqZJeNoI160AiukyzqtqLiQhYysCi
blCNqu0aQK4l+frDbePDXcw3chj5Xc6zDuifrOfxW7MafPLSysaM8LKHDir2CHFcCB0BNIu7trVR
q4ZXF+qgrJFCsZYfYD3ZqfaoKZ3QAyOwqoDp1A2351H2h22C5dOtKTiGQ31YwxoxnRIpSL7ZqRvC
vXQWzkiIvh4WW2Wv1mC9h3lAhkV2BYH0pH6NYFPrwi13Be/UFhgdNzk/lTqdxEfTdX9K5X5eJXs1
32JbxmwmMDAaw9kJ0nP5gm/OM7svpHPY5PEtVxriKzYfje1FS0y4MmsNWq6nLkPdF23FYs/rlJLV
9EcQif4uYyktMzwtOm9qjpjM7DoqMFi53O5Vpg/mFQMNvD9DQzkC7hxfYbEmwGu/qL/3F5besE4J
2rAL4B9zf2GTM8AFefIA+HA4KosWZ+ZYIW0TI9xZk/5qKhogsmGO6UuiPbTZfAqnWMQpVSiEeLoA
qC+C/H3gi33VgSurH6wzD3qyouqMW01EB0YinMayEhstedc6X6k1AhiTZOObJPpxRGVkHEjvGpdC
+BAe1dOWBnz16MN+0BKhrL5nNcrePcnlUvlGH0+duE6km6HYe9wEvvqNt5QRgmqMQ0L9bZC5DQbV
Gp8XeTIq/eGnihHTHUi9UQjwDg+7NjlrruC3wiwqbWhuf47yTFHWqIdV+a7dCjBXBBgbg3+2miPE
/QbQfXO0S/bY0YMuCG10oaxxgK2Cw4fLvkzBYHCzgfVXdRFIbOPpPAV3Opp7eyfGUQgOZILF4LP5
6jNnl588caG1CB1kN3BcQKqT94tpb91vQeAhiyKAWa+tP9Q9vDBAXXFDjmfSm0HkArJ0vzPkdQm4
Acv6Jy+Vy/xgNbnG97/aYZj8CnhnZC1jowUUG+vRA4qr9UihH0t+R241705XXWwE0H1++vIv24vj
kcgYsFGLoe/py677kT8WKbeWG5XcXvookXVosC/cBMRIchMWx8G6TvDDeEvZA+yndB3DqEC5Hohi
+puIgaqDQa2FAl8R37Lp5TU9Zzp9B+bcMoUdoPbWA6VtV2KaZHmP/NeMAFBXzO1gJ/xxLD2tC5pd
YAgAbkXpES+yH1T7ovFa/MTkB8Z0t2m/2DxKNhat78d7IuDE669zvMNRAND4OKaedKzfJyCjbSwp
mHLNxF5FWwFg0AK6dRCXnuM5ia8Y11q3z3bOfFyWObIZbGVoR50VYFGd1zzjEhk+CboEso98LU/o
RQbfuz7N9B7Br6vcs7N3aW4cpZ02vnr50w6MSPcDObXdSjPBm0EBexAtysp/YH+SkWoZSR32rUWW
dfI2OmIPo8WY6JuJ0wExiK56FxBAfBBLCjL1+HkVDLR2AkA3uvvzTd63d1l+3Iig1bmOQD9OdLsN
6Kgn1z+wpzPGpnlxfYTkn7/7AJvmj1m7FiG1ZeGQhmTmRNG3WYVpdXRvVBYhGrXj9vzVHR/0Jtkf
+wNu0la9YUWQedJjttUfud6sk9fES9vpf0QxHloM/J5e5TqQm4zMSXXNZ8g1h0HzzzJh4NqsKjHJ
3ZlaF4/DSnUgv0f/Bjzhc2k2ZoMDpIpgy4iPNpwt4cxsFQW0fEij0+n6OVsAhtTNNIgnqHallfRW
txRufXsE+ctmVdsDGkgPLGxOlFlIb8tWmUVIF/pdtXrj8L1SH15i0nmGEyXiR5FcI+EwB2qx4PpA
QSAM7wr/1/Q9/pJMFhukBpJ1tIut06b8WO82z/Lf4waKJzZokKyEe1z7T32qGVWY7oxlcDY5RbSC
GKBiVwECg2LPYN/efZ0meBjQLKJndyA8tfJS2nAPC1y1v6T4mW+S3O/vbr/kvLUiUKGFD5HzwHCe
yhq5HL4jL/6qn3sWfhZD6EYwSqs3h13wIofSBa7ACuzwDCxiollL11Z8QVazIPm4q0Wz6HzJnrkz
SOaonsdzjUYYOmpVZII2GZ31uJyaU4c8UARYohuelVNOdQ9muCBMI5qSGxukhnNZFKVm1mCteAol
uI2tbrs/vKv4HjUvMi0By70+ojU3gw+a2HGVENzstWTrzhn1R847seXJbyL1G4O0Wi7r2URc6twO
PSWaPeUdZJorFjfB9Bm5VDvOP+Rg4rVsP2W42pGIfuy9mn99j7twqyzuIm5lXthKb+7eCcDVB3Pw
A/UkE2m10TL4wKBbsE9b9UzUBDROsbxb4ZkZ+DyqO+sczkwFvnLdvtjwMiubdv++iZDu8RoT5bu/
7MZwx8EMwBdNn1Tco7TDg/lU0CZDZQbt9GkGDGInXTxsfEqg29E2XAIatrHImZs67yc4hc9w7MNg
d6ZFPSPupamCYNCYdLEUMZkVvArwm1bB53D5Tu+1XXCcw9zfhHaqrFH6R5sWMD+yhMbuOcaMAhUH
wmmW/6Xm4sM0Ml3GLd5ALKtph36MFyA08/r0DZFX3PCUj9QzJeU8kZw96k60y7jAkv7dRrk5bczu
DF/eqw/V9NPB4u+ZiB1CvYadvnbz8kttOl81kn8O4jM2utU4lFFuBG8tJ9saa4w0zFqVyz3Pr0xZ
ZA6BGlBfOrHusehuB1KpMbTXaD4oR5HPPWpNwbuaqNM2DIV/weL2XEfa3hTiangH2AlSHrttJjz6
j4jjIU4ZDAp6dlAhYvEoVc0rM6bvTHZnmL8jI/LPoCXXx+QjN5BVS7QnnSUYCfhQUbvGiAON71AH
StsHIO9VZi4glDtX9LldDo/5QQlSxJRxQHKnVYSI6SlmBmGN80LQA07f20FhHjM+uzhZB/O/awVc
OKqgo2AHXnaZePl026mypqtltmZ10adDIs1m0+7RBRPW8fJnTWLzELmA0j05dzgcgkDRfA2cZmd7
YuaxcKjFhhsQe+5WmFyvP13laX00AAxDRIlSomAYWEJA/SbtSQrQGSkEeTFCiiwfYI7i9YmmGGWi
/55Mn6Rt+eyIsuUkQD2i1f2xLRIf3u1M5iJYuEHt54tgC576gAGaHikILc2DYHu1j13Wedqe0OKO
3QXkAtnjdHwkqSoTQiPjtqs0ickTo7ozPBWuDPOMb4lrJfo+tWIBOsjSRUevjXrx6JIyqEGpWXEh
7UPVsgKO7ryPy8Zi9ZP5ZJTCQ9Bts2lvEVmr2FqhlqBgFORrC8i5HYpOkY2F/6doZTzZY/11F0Gp
YwYUNW6kJbNG0+b8uuPMrqmR587R+Cy16YeW1nXURx+kdiinj51jvKse/uAB2G7+Wdk0hiqKna3p
6DpTzc2Jzw5lr/mqn+1EmV2EDiQGmBn8OJkT4VumQbSYIlNB4pQHZYKH2hBdDjHfG4aPvCGsCLJy
8pACWO8N+YBBul/xKTn90fDgwugCKA4hByKArj9Z8Vp1c/dbKisAqIIbomYYSL+vU2hF4WKY1usE
3krej/0hgsEgE+MNB1i8jkZv+ZYDobgSAiOKe1PYA8KqhBRGosMLpFrnRwPktlXQ6f9p+Ci1I038
LNj5l/patcKYEYm/ANEK8L9/98/enVd9954K2ZriNk8/yQpiEXeS3bYFV8m1vnBCCN3XwSMglhHj
WImWIoR7IeYjVepNHrv7foLqbHcpO7EInD8uMhBMd/YwUbsFiLz58Q5qBZq4+gPneFGjFuHbYoEB
/1IFkVSMd4mTtBn6SE3fkcK53gtptIQ3Q33uOpRfuPZOPLDegIUxEVQA6FxmlVWEshywF1CKxInu
LzjPXn9L0xcDi0r86eGvoVJ1jPR4jlrdXy5UBkp7VgcCuurb6OeUkshoEAVhAP7bPxTo87y1iuxH
LLrUkePMvgWnjy3ncW+gNaPknxJ0rcD265V+TauMCiPc2/z4fmhdFTe3O1HJ+lPnWD3P4GsUXlrb
0kP2qWAAWVnvdeYTr2Sn1bXEXxu3b/GOlpcQn6vQpvfldtF7KgQordzHI4GA41LUx8xJFutAYMUF
SSkruLGDIpNpj6NfClt0/2yp9VOTK6avUXD40Awhl6/4KM+MaZ5j2HSMVNSUUfjdR9g1pBgatd1H
MB78sk6fBb/2Snsftj1KNxwnEGisp45htwxyZD4ghPzoHKmHMVKqak7FePdMsDlEt+urDGFNIPpo
ric+sKF3pHgG2d6TtPviieDbba3Pap2aHCOPxp8sITUEjVJ49H5/UICiFBYeKgtCgUWPHcLglvmw
9bbD2Bri1RKOVyZIwjTIPa+9kGxGc+EJUFK0IGnLId1IztszKZyaXUfPqgGANLZIPStjAFVIcnnz
I8J1UnmmzS8RHxjnW6J8ucZmcsb/ZqOqfmqnycVqUnmQnkWZdudqKJqs9Ykb7/RZ2+R+qvA04x+I
KRO6ooc1LBYmnzAxQk3iC+PA1j9AXaENcN758noU/4yszaBVH6C03IBQb9J/he8FlMk6owTfhOnn
7KwmX2go91+6doTpcUlgA2fYn/PPmBgMW7XKAN2vZXPO4FZrCu8wMZ7Ad7N1GDIEdHpERZcuCqE7
oAztrBjrrj/DBSOJlbMZa2WTagNfPRo6cV/zfXc1lKRxdxw2Hxd318YNHw/PbQqpy8Tv0/dD57jD
sKMcjWrfH5K+7Ft6Hrrn1sFhkbuI/fgNSLgAbRvSjnwT0SCsv7lrOtyENqcGMN8KHJNwZXFsddso
za+LTRB0TevRpKOGJX9inOlHsLtvxG8U0bgvmJkiGsATKmr6FxPa8Xj1sU2zhfzOEUxBbvxLktr7
scOfNK7c6lWZwZ/qKC2E5nro60qrVPoXjB0XjdNeZec4V5O18E7XdTRGrE75Di4FW7v0I77pFRNZ
OVVZOdiZWJcFREPlwyjIxTbmIgSFLt3IUZ/WRaiDsciwGWINIpnjO24uNC/mTqu7uWLfkp+Qa1Of
B0tV71DCoCE3USHu9Sk3FlbYu7GN+6aR+G6nPV/ViO/GMhmCRL7uOZNpKqkrWOq90l3X+4bcdgGc
bI88MoDAhc6LEr2ZLZofHqN/bztaMXxQemtpwdXryn8R37QwtqhjC70v6De/3zBJM98RiZ2a19Aj
n7TTgPv5Bb5CHuQmknBC1DKNYpv0Gum4aPvTExehgeMeHU0mEiKOXNoCYTSfj9fj/ZRNrdYxU7e9
KljX+gnm6XtGEgE6e7fgBHXA1EoHzhRd3Oa+nRj5I/3Nx9+xVdUbHqDFAMqTW9ib9+7PXVArpPWz
4JywgW073rQRTwu8n3FPrXEAWZh6IptVMXj0XjKGI5cIfBMw04JKgQfAe+lbi+5jT+8ylPIe1N5T
04UX4s4VqD7SDQ0g33rmzVOq7nK+Wp/nEWtKnUQaJagpjxdFWlt7iZu0HONMExejdsa2HteXEQPG
HYZO3+TRlnrgfPjvWcUm/d7HhVD0RafA7NeMozRVfY4WbSEl2wBM83QiGgPYXY5SMylFKF8fjIIs
92q6jPRhMTyFcoHKBeiq28vRwAIrMrtzZNZdblMVMGIG9Wp7E0CBkCB2e6Ec5iKOio3EEeLLsQeP
/RTfTBDSvVsoftsQlt+u1LSBj8Bguqu96mPsUhYX4ceWDgHUPdMVbeuHlfZsgaQh+rtO+7PqeoAe
wFnEEGvnminLt17b/ObtWkseIb3SiX/dV2StgRPZNIlCdiCSoKAnmnw1heUdX1wITmwT24oxP/OJ
pF9+wDu/hawaJ9UqPuYNgiY+YJkw1imzECk81XhTt7qd0BsPm6/4ZytxJeMlM7HAvomfI1ShV3W5
vOqfXbvM6yuTa46xHRelrYTcNJPdzhU6tm6LeKldEDWwp3uo31hmuePqwi7ccf+NugRYlQ0xiqeX
TQyd9xiHYCZ3nXn6eMRm1g2fdb0WPBVf5zhvxHjIrt6jTqSgJ2ekxRuE1xfli84JSOuodNXJX98X
+rl7J06El+qVaqQ7FE+EgWOsKhu+ATPGNRhG4nyuY+9Ztf5LKsmaxVLxV8BojBaIumGm3spbyiZm
tHE6ZFDz1AVXQ/HNXRPui8H0vQEA8F3uMy6MEh0iMRSRZZqkYTfSoX7bdEh5SyOhlSi+ikf5QJIG
Gu586u9Fq5DKSzkpPBw6NYWvyw4Ige9r2rfn+um9Vn4uWXuiyRJ8EgdVTmGhET8fEF178YfeNAhS
d3CgOC3xgWW5uCuOvrawcpOnjUFw9pDtvP2jNaXPmNP+hhurAnSSdKXQXCLCHc1w2pqBhkqkbwj9
6QpPsFsgfzDQnCQSzZAr+44HlUj0Mmag2W+m4MBzS2Fo5y1Y4af6gYpaFeibM/exd5br5A0cghII
PyX9YZkYlydKm/acbgYlAQsxqgndfv9pOBH8Cs1QGhzRlPqm6k70xwRNI0RidJgsfVGTpvqlLp6F
h5xpf0aZUX5dyUtioaIeZZAeyh7Q0TWY2GUdeX1EoTWQ+vzk8jfSMj4FA2yvdGMezejz/dgoTlFC
zWfHb2EsNF0GER8H0JsPm9MiTbGAG01252O3vUYAFVqQAZLjy3m94iNFsVaT+WC6vrMW/2gwWHFz
Ghxe/7GrzmFrdynWSKvb+vbedhENl7F22L1akE6qnRF/H72ZsENd4g5DYxtyTLngzhgTSJEUvOkP
hwJaU5ffq0Isu55CxM8D6543ju9QMr43Dm5IgLa/G+vpvH60nZWGFbbyEKMfDXpO6BpDm1O3LpRa
XYpfykIQV4GRrUiEhCM/pvJQWvRZ8EQ19UUjf4IbGErgWB30KPI200KStUKb3/qyjBHPE9UZABFt
ji7vIuLotlEPJvlnZvlJ/Ykg0YuPRVZCnWVa9MHe7aLy2PUur5JERnYjrV9al+dY0rGgHXc6rco6
28EUkp9OKtO7PyXtffJu8DeTTQWx1V/g9IFyWtpnUH+kKYD3dch1z84ZLp6l6cHoDKiPT6jBH/d5
cBDTiwLbLw+DtmlyqdmI5T0ElWwQOIoyLNBh+epg94pMAuAZsGjxcNNG9vDpA0wr+sHJGojjJOev
7icJxvtgzNJvnD6bwm6hAMqGYz+XOYyj7n7qXwE8CDPJmVKJCzFFM95fBce14xWjnScDcOTjZORK
kyF80pNvrpDfp/caA8/jDyEcVmyY3F08jwVVBRzWMPovue99q8nDH4WPErExi3XjVzU4MN65Vj5f
l7KgST4PRM84XuW6rZ5vXEWwtknhcXBnRY65MU/Arb7bVLFx9Tbf7pcIBSnpNgSdZeI+lPAlTxkt
z9f7gYdM88QrowCgUq9aEB3PepgULF0y1RWPI1QH/nh8FDruqP/LusG5PSlZTsvJ1gfX10CGlqTD
xQqLeUyOwGl71bem8JlD3+mEtUNL5OZn0W/vMn9neGNccYXh88s3FrsS8fl+r4AmLIipZtGK/8sS
/muvXKDPlaXgss/mQez/o9d9SAotTFBh7SRFneRTa1ZTt/gUUr12LTK2VtnwTkHsBkZYB+v+5JuL
deF9XXiEIFvy73WYw4tlW3wLlLq34i65l3E/nm2wZpJsu/QuPpncbfgn9KQAk9Kq+Ls37r6bw1AL
5+Q0OeCzeOOO8NXlxv+zvZsUfX+ylOmR7me8Awmr2kpyZvG1ZMVC6rBrkuZWuhYturzsFpU1GzJV
Jmn8MTwqRe0nGFFZK2UD6s1ae3KH3nuylzeaFFLLbKzaarqnJFc5Y8786W9gkffiwsmGhx2ObIAu
s7GQe7SCmqj/QOHHKPui3NnRAyiRg63dsGVmh3++NanRP5epXWVT0EK2UpoL3z7Ijjyq7TCHBFxN
5mkY9iT8QiPPwrgsKXSR7JxoPKpC29ZOHJrKrtkWrtYpMsRMxbzcEAkuWWRO8BCIiPa4Lt1typkW
o6GXQGEq7Y1vNkumfGQar7H4v3wmat+VEPrqYKcjEhYft6Mxm/wUU8kQ64MBld3Cg2GX2IvmRHJt
cnEk80XbxtEch2hOMBJW/gjsTSZMdWDlULQpm0KPTTKYdo0rIh/EL1r8PtAZfWgrcET6jIPWwbaj
wxt4R59klYN2lCs7LOSBCthJjYKkIIAHZ5fdCM3n2+9t84HHC/pcKeegZ/iyM2s4XhHx33a0kB23
nIIJjcHOAkexMx0HooxkfJCc2VH4vJRQ4SWXZuzzqVJdFRxGvokb44jUjdR4SKiBO5A7gaSyvGHt
ViXM0/kMdotHEsbcvhJ7i1hUKaDwbIjtXuJSgr3lDawX5xfd+usuwo/y3l6VklL8TnsxnvPIVz2v
KbUD4s710y//1gufFhFf1mHj6EKt85UdMY9sF0ITLMsu318oN4aBXatQo17aGB9c8aNeq1ltFJ5q
DeTfQysLxbggvC7VD4p+tFUko039cNdoNnAzELJVID2ROjScJjdizATmpch/ZHGvN66oGPmeiJ6o
aJLQ7L7REqxjaP3qpiQWg98zK4vv917iyYfEo9fVr7DgI1Fz3Q5kWsKOoY6oX8BOdPL8bEz+iNyI
2WwHlgjKcDF7LsAa61z+d3O+qZSVgjYMNXdsp6VWNSTLFzOkwdQF/YCyDwlkXOId6uF1zESYSU5Z
WsUnkH7Kv+gkn/21UreJZSitbRWv85ugZJpdGxlBqO9xUWORiBQvQJwfvMEYxDiQQhK4f+M0Yh7N
1Dae5V/2nD1Atp+gqX11Fg0uJtVsWQBgF8DOTkvaeP+EBbOVgUrsm4v0W1EY9F5IMOILAknKshzj
opWAfR/Q0nL7fAaYGKom/MabnVvQiL4Rd8WLTsALHID/GUEAX3kP++clk/2saGf9cqNquTe4q+P4
EZNAsyCw8OP9x7MC8e4usKcsDFX3d9261aHwdzRmlbJw+O3uhs153nOe2U8jHxNigjfjEq/580y8
x8fmWc1XXUlP8VbkLm6aIqbVJEXO3iEKLLet9zbqo9wRGDW/mrysj0BOEdb70YUXcRBJ636awNh/
hAPxHBs/e2kNAjvHxeaDXPUkiQRtRe/HwwE0KaFNAbmTtd6If8IvCSRiSGUpr1CxMYazpeAAwJRd
lWuz41kdT+ctwS4PxfOhhOsBAxK4D7OLOPuEmzl61S5vZzNfOW+DJzs76CHSqLoNQyZ7kxwrjwOG
ytxQIzTry6tL5F8v8JXgMc++aLIpBuIywcjMuS84AIWMJiZxQ42Oqb+PVfy2MAegWF/7W4K3zzg7
JOVVAh5dNt00HVp9edtnHI/kgsQM52uHz/28AsAXbAMm/Uzc3mZ4yhBpYFdqUQMPEaa2B4OQR7Nh
XbFPoYy5UhdKlxS2HtcJgzBV3xyiB34lVOxYnZaTybytwyTXXyluXSsNYxoohdHkIOHA97JetjwA
uNGGdRY0gZAt5dc1qmay3dYwV3UjxZJY8q3MeArSp7XfH8av9eeES+gURisP5CRd+fLiTW2iPFX5
3xYGPkUFA6ulnevoPFgg0PhmkIZFcV2zzBlPWQPLu9RTJdLdWssGvjZAh4MSDKm8UWiGFox3gaKJ
0k1ycB2vT64YQQwr3Q1+GbBoQIwTNg3sZt9qYu0F88OUzmbYdQJp/FkrMv0Ih9+GdtiNPPT76rlD
vbe1179dcXzv8JvrJIZ1v7dw0JROkofBx2YoB8xhVpUR6Q7GwoqVPJpFAln5odXcOGY7fMi5mHi/
bUE2QWSZ5jxtmb59QzX4OIJMtVaWpozDH82VP99lZcznMoGtvO3TCWsK0hqi+mN/aMLh6YP3baAY
oV7SEC4A+OwojbIEfG6WHXyc1gSJqbqH8HE8Xw+/UY50fUQ7gETFYuAQ1C7mzVyNXw78eZ6RfnMb
JLSimQ+pvjrLfaVZ2lYc351w3yWTysSElHa+N/MvYNsvpLoyuVtbQj6AJeWelO6rSPTC1D5aEsRx
B1xwh1eRNvenZVvKl40uRwXEsSqjOFJhV7xA05mh8lV5tNMoA7N6Sl0Wnguv+waknRrpapuOElYg
UIVWlBjKMYY5FCQOLeZ0V6pqNbGxbTKfb6AgbJ/xt30/lrPfieK+4wvV39hMVlHMSAt/mEgFGfEK
wPkYlKuZYQDHFm7JVDGiun5s4gsPFZLJbGhhT7R0nb4ko+2Ioy+zHyBtr881fBr+2jR388QJ2L7W
oX2y7mYlEd273sx5gLDFQNRTwFJYUtIomQlhEh3CbxxmU4nQqoUeFFht4R4/tFQyVF3auxjEzvMZ
yNZitOUOpypVvvDfX3CXFwOaQW3fsy5zhdfFZMvWeG/PxUgT1M6ZmKNxD2RVCj3QU6+JDinRROiD
4TF/DkU65cA1V8iFKqYoYgxpIYuNHxX22bbQjepc6qK7d7Ix7znXt56+TrLRHUCWLELSQzskeCk4
l/W3WGC/o6WhBEWa9gGYrl0tJdD3F0AtJ4crcYMrq6M/pqOjSi6lOfE3GWYHyzNkEseJM1Xf9RVB
C8gMqQ5pJ8oud0aS6QBdTQ+xqS0KDgtYV6GQ6EXmqtBoh5m/NCX88YAkcLAspE/B3Ldm8W3FVMj9
pSnk0iK73y58FUUkk6qJwYJr7NopjxRCbEV9kPhWq0QEmcDw8yadXzmJ1ZSvQJQghRQDpvM+a+GV
itLzvwfBwGr6EGRG0kbC3bC7Nl1mY8/N0z9c8dua0INKnFJb4gSWivxrQG1MAR7BlIxXd1msj0Hk
G3gNFQxXcpSrFNbHV+fSlNHLquUw41F6K5q8hSx5DvzOkQHK8nCFbmotx1a+1A9EAjGMDEkHNzkW
UYzShWMOKkh21z9GPaQ7jApQmgiN8GWteZqp3c7GB+zXe1kho6Z3Omd/tgnJDgMcQGmfTPP8YJhU
GK8y3ArybMjmjp3UjEMd/4dZi1L1WGDfS+byMkMNMxIg9n+56gMjdUjX2GeuIHIsLoG6THoM8Q73
mmk0AV3c5IeT2ys+mq0PkzBXDrFUHnSSKrVw9/nhutm3HVmfUzkcGLlLh4CTNUZwEdQvC+CfhyKz
Z0pHrDXfaq9aGs0aGdeGhyOKvqTyHtlwt27XP1MPGcCSbBAL32FO6uwu+Ociu3R+xVBXSXVawnI0
kJo65qN2fMEuI7t/vDqY5wxUoJrK9zQhGwR/2siPZOeMdfhcM15CVQDiUaekMocFK9oqWpntBtiM
k+UGkGoRuuMliMYHFVqZhLrddggPjGHb43tcHa8fhDeDY8aN510Du4mFvUPfJ5Qovw3/0anvbW4b
xkSYieq4R4Siu2hDsr2kKssJEm089xSluRJzmsPuNToOMYcPyxvHqsXOdva8c6fFV149/G+Dnkxl
EmM82x+G5QTgbY/5Vdb1qs5TtDMbzJZy5zyvPz/6mzdpEyeWf0m9WwQnigegBgYX3oi686uDeoxH
mz6P3UoE83luhCUvHDc5AX+dTaqXzEDqiwgV+GxP6IChHgR8RlEJpSLnDpxrZlPGQwiXbYEFQTM3
QhNKqeoEtlnU5fEtAhYIsn1u184H52V6qyUlmvj5NXjDzQXzwuPDVTL2VqMeZXyecnIcQR7upJJ/
gob7ijbKYZZbFwR3Wbs1te9T3tjlcYPgFbUC6uaelFzGzaCpjFOYVJ+cBHybjdNCHkqCWQ/hl7rU
CEbMWMZrVUeEnH724+H1dstZG9GzjlqQHbfYgQ7LRwl+QZgISSR7NaE1schzvOrUgrumntd2iOTX
6lmkEdGMU7GM96IrMDkx/EVzzZRipnnCeRKABY/WFMNSDrtCEnbozd2d6Gw2XYiEOBLxk/X//AiY
MIFF5lW9NR/3DSBE2dMiHMln95ccaF7UCnkScqVY5cZdJckwnbj0d8WI9Q73LqGEsIQVDv8QX6dM
bc1wDc/1Z2bVNuNfxuu8otWGwfpWNEhvJquEzN9M8MAr66OzRVrwRq5gEIkCbAmUPTLt9P7aFa8J
yxBLE2uDLCPld3dYWsqzSLYeSZtWTOZ7ySXU7jaafx9O557SuriBbQLuY3pcs93Ftog9z0NatHZ8
V5Y1lP4TSSFKIyHSe1TprtRSNul9I9OKoJlo7uNaezlfkxLgcL4x5RvWN0Ov4ZJNJEQ0cHCWPBbV
hyUKGSptwpteb6PTh6FbIcrEBGq8CupqeSNaLHSQ4fBnaiTe9d5mUlbYiKsEyHXRigpP66+Wna9Z
+h4NY3mtMm6w4Wcp8N39RSOMPC9e4em0a43jAtPrPR2JmaPP5Ycrj32HlU9gWahAfUfGmTizj9Nx
9Gwi4pCWL+/Q3drDIGD2tYI10HZaUxFqgvzQ7BXZK7bCMmKVOcYsf+8y+lE31YQt+djw7oku12k/
S2YHjLD3O0Q8CfC7+HJNiFdkecGNubBk39PkPVmnFdVdpaJtrciGSr9EQLEwC+mv38Li7XBZTImO
RiR8HEFERSoq2xdDDQo2zDc0XvIyQVLYx5y0xthHSok7bWDww94LKbIMFPefKqfkKC0AwyKYH70g
uQ4dJtcnXrP/iYsLb3w5QMn90DDtWnyAOP3O8g0Vy0/4fU3cXSzA/7De1owUd+mFAluZ0exoqat2
KRE5dZNWOMCRbbs5EwxI53z9JeHzgiHRRJ8MgH1V6g+zxRUHWnXiSxOOq0ZZMJS/9nC2byVmUmot
RwnFkddrf+gsdoDLDI9FSMHMoG+PxNZ/60D7aIgiAfKKN4Htt1FqBwmoB7M28OOfia8nU6uqhyJ9
9iWnKkc7iplvICC077QH2mWEazqNx6Pn2s45otPuFkiawceHA0fu3pIte1Q9NnUM2avZR4uTjz9j
6jOo4yTmY3Jx6FR1RgD9AjsJmLse01pmYyV3nIhrrcX5Rv9512RDI6udRmrsK8qb3Z3tJ9QUvXEV
Ohc7ckuPlIqy4Bof6lDMMBcc/OiL1NWl8nBdyYO8voaykMafm9ToDQXTgtpXPCz87NWyBexc70W8
xiHGAgdRnTYLifEhUAyJdtNtUAvA+Vs47qTsr+x80nl63rXiBcSzmXj77LnkLP82p07PzA7JsSXY
wagykGWrgNIhJVTbGappxwWnNmYw7zlIkyZp5w3y04SY0L0PAC9xkP6Lp2uydC10ritXBRRaPE0v
aW7kfghcWjLye2oy1kEFo1oBuhpN8VPpdelz0fhx4/tF00JUO0TrjzPam0uFSzZoIYbytlNW0puI
qkv1uCP8zgcrDxIG2dnInXCds7KP5/jKLNnVCCxEANmfG1doQJrYzvEVTkw5T7DJpxUTM3fnYEv8
BM2IDAQ9xvQE/rlLiAlnCBKSSVX+l3fa5QI2WYzg4Lza4OP/tk15kVTFefQ9nHK7Hw4f+k7ZVeFM
VY5U2ttO1SdB92JpyVQ54FpNGMWE+bvUiWL5nG+7mqeonEkVG3YruK3sg+g3ugRJmwyhZntCOsWn
eZkCuU+J7f6OkoD4dvcW3g80KlSvp5OdQDCiUA1QfTsY7K7piqf/m+glgO1TnaqmCw1FgYqPPJc8
Eg7RWwW3zqubwgu8Y6VHnY4pFyg0MU3QWNTHkFPQAQoGz63wEZ4f307Qc6QaNOvyfT3UyFbCC27V
hFgmcd7YWWVLrq7rt+XUCjzkObSH9nmoF6a2wxcnqXY8RSKm3pwMTHIg6hVRRK0U2JGB50mV1UmC
zC26J1LuOghKMdynSj5P3ehy2Q7lGZhjB2gR+9D7+Gy3Rdt8hYPP1+4T2e+pbXmyHpubL0XJfCGI
xD00JtRix9bKouomyeWjQBmmSs6zKarYGFGNOAbYvEUY8AQRXmMrZSN00s/17YmRMw5KHbSmpiKf
g6uUTpp5fIjLkFkfKBPe2+mz2QxIyI0PN0f744FJ6bp0pZfrKsbMezTqOQqHmJf+b47Uo84+liy5
hcCV4/mfSJdUvNxH4MKbq7cG/Vb1pCuCJHag1NmV2aVstre1kXYRYVsSkQ/VXFKe+JZmB8fZ3M1K
1pINIWGSMK4cLqGCvOER5ktmnA/MDYoj55PXo7Rc6jhKv/iTCO1lmAJoGOst/Ain5jkLzCvvv8Jf
R+UOcr+CvaI+VYLyWEt66/CypnkZk35BqC8CMS2QXZjwW0EvaohmwOH1cgPZN5HJkDSKp1D+MzSa
6OGPiXR6EMak3cjklLiuxWY0HEB3HIENQRwienemZnLoFlcCQjrkLJxA9KD5v1g7t5zUERVsN7Rn
6/Tbo7hje1tviknPXw0XBoprC6T0pWvTogG6sm0oJ07/8yD7NBbYJXBK6CIDW0KWWD0bxUzJcEDW
7ruhBlw7kbEas152kzRtOCbi9wytm2WrQ34Bqy7lCI1P6ItbDarkyZHN2radjfn1/yVL5azAn/bI
OLBHzbQuASJnUQz1CUGJX3rVMEL8v5haRwMQaKtRAyDXuWc0cOXQQBPI4XSsTSjKC0+wgHxKRonx
vFc0NczTFiVHz5HH+3qobC+YEtSCBnjgxxLMumxbONlXuzY/IdmNC3VmUnK9zMDf4MNhVv1UgH/+
dCMqAhhSeReFulH8Jc4oHHE1RXmAi8x6xA1brmgrvwSJuhK/7Dfg8yHbXKztcakdzGXj1CImjgwF
bJGGRMOQmJvaP15rTd1h1aedJaNlwPEwt+tchqf29PttVZcYXIFoRIpiYdOaP9gVj5h9kom5+D/D
uOZN4Jss0y451h2q9p+IMPGGXvwxwHq5QtAhprt5/u84xkok7dBd140rk2tmRLz+8+1tqfgSrCgz
wiFnwZH4KQIxZdznmSsC+dc0TdVs8+xVddwUJtWeMEEL38qe4aGxbsJfnUKANO2OjE4nmeq7FcZU
T7xZr3NBlfjkzL0mOO28p89MJLHlU6ecTd8X0cuLHgP6Lt6YXFWD+DWESAMdJI/cJeixtiMqLgqN
5pmMeeyQ7qFoKv/6nRm8jdb8kFQqv5pn+40UUwDC7gTGdHd4qbtdxqSMp8o03kKLijwF2QgBaeMM
I4dyzZOrGKuZeI3QQ9qGul2sfPdFUjqbVtTw4XNyoxcSG31ul/G9WNhPAykYuZhRQ4WEdlVj+3bk
WlEBCQ4vGIldEwXo3ScF7P+AFDxAsaYgf2+TvWum48fwgGxFWny/dOFy2f/XyH1ojsk55vWQHn/B
rfc4abUe+GSooVFdY6nqd6uiQDB+rU/Zk6/n5p4Z7jXNgd/sjs7bESGOGCPmEz0nDEHNmji2nAmV
Mbh7b1cYAMVU3MEXZvTpSTlOLzCv+vyz0I4dnAqDQPAXgL2q7mUbf7BgEOB7HBYVELppDDTrtq5I
YXKdpnrSdp54OGvByI5ENnV2Wb7aK5WvNWkovvHYQTAvvThrbCQMFG40LPt8foROV2U/9bvSTkdQ
pTJiXZLBaQVT5dvAf3S8cnnil/3LKBoIYAnDc+jpWz+TwooOYZeaWAsVVxetv9TS6NKCivVJAl99
zSubCnaT0IVr2Pv4vtS0qzzufPNoVLEKwjXGjw+k9lRSQsqQ7/Pb3h2YICKUFNPEBqmOVdIbq4bC
IDj8nuqKQSGLNnci9CJjU3IquTKZi1RaKmD9AxKv9mgjyTpc8KcQ3B4lksOiLmN51Q1pE3uBuZed
ehHOx6RGgjHWOWHJ+nkCBlRrfBBWk9IdtxyHE2UEPb3UiguKiHtjFNef8jzWXw914sJo0WBbm3pY
OzVa2HspRe6pzGisMZ7am4y4Wg+RTdRas7iFhJMCOgGA+HfWXkFq8H7bfemJyHMrkjgoG6rbrZwV
5b2BqSlJkM2Lu5FxKmY7c8q3t91D6YOpVgzJLbA0j/lTm5Utn7rvgID9IsY2Xr3wEbhS0magfH4q
7TzU1Xal4ni4HwUBGbdZiyds4avaXe9IhJUMV9EDcVhXi0UQ8JVc+kEaLMD+QhZQRUUKnSTSTSbS
jdYpkSFUwW44EkiYHRqqAzsQ2tle95s56IUprZgxyGIfhIL1EsYbwfzHkVyG0icVNjCrW2Zgw7k3
iNpJMHpeJSEbCXNZXRjhOVCndvEuL4sTDtKhmIccYe+J7SGOw4R40chYVFoO4FZMZKKelat5ui8g
OI4nl4u3DCrMmZNSbDbyYy61d5LpKnEvXRJqhm45tRC44Gh0cy9nWjlRH6BR3msf1KeVCEDV1sg3
ohM+Nba2XRW7Hlqho7xZy2swx4zaDawQCPByHCRHoaWUNn+u3eJTqZmrYfw+gvk1Vkj7lfrzD4Ki
LufSr5WxnwH8B6e6JNhuhLr4DbULxzodBuf4jWJQ/J7hvPMDjQUb4QDKLHG1WLEPli1je+JFJfsQ
sCfLuInMZhp81gsomb/JZZcDQZP4v2dElCgxPkJ4W28gMQc/iepDp46X7kSp/G08BTpDAOr1HD0x
qxo7jYt8VC1g0hI+1WMVu5k16y0Ke+kqcKXqx5DUeTafUpSJwxs4c06i/vV1lHTuiVDwbUgYzeYU
0cKFqBgDFmN0n1TQGKlvPKUp7b3kT7uG/XrsSjiUxu/jdlTS5uPDxLHyPrSG5oBfUNj6vvAr4dxB
F10LuCstYXceHT42yFNWpHDGL84IBt+tWb2EIWCyJXVTqbmJoE4+C9zkPsn6etKrYKF2aPC2PBSJ
zGG7w0JDAST5HhYvLZGARjj7DTWIbf30NDt7ni2uWGyevovShROce1g13ZDUQKJQe/6uW6I9L6OM
nS4HPBrTdPIH0JpQX2+EmankKH/wgpY+Nri5XpkORK8fSEpUYTJJO0ZlsjbnZbvEUoZ1f494Szdt
2OvQp/RId6azw65ohOON//A1X3eihri9PnqkwepkCoKU1jKFeeKJK54v9knr5z4lyy6OBdEOKwWv
h0j5G8vPtNfqx80y1KBjq414K2H1Kl9/hs+8fE53fYJCc/tLMHnoqpEdfXagKScl7oLdg3mC7oyY
aC8SsmGcQZDSkLqNFjX6US0sVL31lL4+ni4UgDH/3uLm30P1xyG2DOw9j80gcqQ7MpCz0VmBZLZm
8BDN43EUe/TY+3RpAfFOnxaP85s1wc3ZrsN84XbuKdQoLHfU+061EWRKjZv3U6i57R5xFfagbpZw
HYUqEnLRyIxFC7d2MM+W8WT7Ht7Sd4Nv7KRGkyrLEPMUtYJErOvIFLBg/LqVXizaQZAS49Kd1erh
DBViogT3yfDSLk0S5q1OBiL52F0MxujPx6BWS9fvhhvqYb2vilqO1fra8jKiqU+xHOQ3ymq3t0ix
GEA6pRaXyq5rJuqSeUh0G0X+g/DzpT/PPelkzcOhsgaghOeU8JDt2tzSTx4ZJIIWhNi4o4Qv0IVM
6+MGmR51mi28AfU/wHLhzSbEojsZjg5QY4vsnZQEjEixj+FMko13bOBbnsC+WdS2HT3eod0rFQT8
PhgpqH49xR28b+5mHYeBK/a0+T9iUD6J27inHrFyzaRLJ0YUh4xM/HKNds96a3fsVqL1PL5TRiCV
5ewLUzdPKcBsBGbGKjakuOKaJ3Auxh8CiFD/o5rmySqCjbNU0ymewgHlwXi+hGufyE+zb7agCzsZ
n/N77i3zs9pNoWkU7TWkZoLV28opf87JO3wd0N/ogdHncv+sqP008cBKwZCktGxHr/37Gi1pAJnN
LLouIZeO49PAbjdyTJIQtssTmN9RV2cXzNdmaiT8R926QKFmSS39x3q7c4trUi4+2B15/hjptZji
yqmX/G4RftIvzXPMDhsUO1KwlEKLtVv92HFsqXi1D7U8qwf77sQ2ZJ3et74C6Ss9TmpF9659GTIy
CctjYPrunfWvxbdPsfUrPgjYNaZMqh5K+dZrj1OmIL+p3d87WrLEc3hPvFiGI6ECCyx2xFrK1K0m
g+QYMUIqKVuMpPARACvKMAFAbvac1m7k975BRa4oh1v2cqzgKwLytGQPdK4vRVF1eiSN/2ZN2hF0
3wxytVMfiVIYvb61FrfGCqVDQh8bEfxgwsME4fN/Z4sMachqk+HRB0vs4frJOmIX9Fbpji8PUc2+
iCjVhZpk8HptVVCt/Aop2u80xRzS1fK3VnU9C8RNQC91u5w2MWjeSWGmRHcDVd3Xk4cb4PtKnQTe
OZr7l97wG6GijPphSUZ6hbkcSh4xmzOpCW/i3M5NbZKZPNro5WwpKIqONNT1va308d/gBU/Ia7nb
X+1zKRbrMUDero6ty6D8Qjr456seasRvGwiFXgEh1KCTU6gS0qupFmXIShS2U9B2s9SJQHyUz6wx
bFjlvMJogtfpafcfUGcmP4BA5EdnWgWNgoQjnDo+rpqpA6MMmovjfmy/ZYZ7TCClVajY4HA3jQZ+
M/m78NGo+5XuxRrG+zlg1BdwpeXHZNtN6yxEZF9MxESABPkG/Hb0lFZxdRPAgyAx1d7ALcsqHZ+A
wMGML/x0ZLin6rKvWp7/bRmcQUdeM5ICSpbXp+XOxVra7WabdOrb2rdC7j3IMsb1eUoI5WfhDcBK
KOlhpVpEL5/7DR8wOclgQnzMDD2aJ1IYo4X05fjnp3O1dH+TMl3pK3ZW2LK+p1YWH5rsUmYvfbZO
tTtfuTkp/sgnBeUccBtsvC6znK3tt62+NPl0URJat7lJbR7yBaFzUrmlOayGn61XR+QUtxMQKxMC
KhBABPvnWy802HOfHZ9umcbHjLTNxduiD6+3k6/otWf23Nrr9FifG//PPPOvvWI56uM1WZe1XuXD
Zh1k5gtp21ifHxupm7umpndZzsigMdOFFPbx25f3U4tEZVNgjhlVZnyKV7XcadJgl1r+obR23wj8
QuhbahM8dezHSfRxnYbkcuLvXWBumXTvma9Al2ZXUyaZZZ0de2AUVBE0qyC2bMuXiyJdjHsR+wZz
ZhwEiPwvi8nzcP1lo9NjsHFsaFW+hVqRZScrL8qkUg7bD5bYX4yrwMWyooO2XYXKlY/5G3Ov9wOb
bm0eYASn0MLDvsew11beSRlgD/0QrDHpuKhFQV4FgQa35PQc5ZaYZbTWY2FKsgSLUa/eXthofO56
lhmo2yYLnzupIZLnH4P0oorjsbDs8GQcs9R9QJM3LrhfJBrRxPsXSTkvvaUdqSSIFvnbVLiXwsCV
ePN/VTqoceU11kG6ONb2e3UDvuHYnitPuwyxZNRMmiZPrKFVLgRxy2EpzBe2Fg2Htw9zF9aKsz8t
emT9Uu1Z3cHjIPwMdzwiCEpK3A7nA9cIqHlMChBtXsm4oVYmTl7ELvTsubfbA9R73hSLT4e6lvTW
pxMKiC5P7qDcH0P+80AZpJAGrY1rxXInQHKsqbmUMCDa6kwVP2zEg41h3ubAC1u1IVVlTwPC8b7H
LnQtMSeDMN+c7okg5DIk0n/fiidv/5RpB5EwL/MS9Ljj3lzEoXagFusfh2hKRdqKccJqlMhZ0hP1
1JNyTZ6hlliYmD4DVy0smFZaRc5WHE+67siiT3nffV4YTja5nHYaTRgoJekAL21H0iEEzxy5gLEv
jE3ZH8KUq7FW8Cl6oCGlc97d59YkjzeWqFANZyNdLFCwvXtE+UA3y8a6tu8dkigE+YIUPa8Z6K7J
Vg6fGjP3mPFbnECu6rqjRr8WbG5jlNWKws0N1u3nxwDVHm7yPBRZv5beGjaiJ4ghHELA/v9Il6EJ
wEda5ogekl1O9YOoTmqxbkeuTZewdXWgelLDb1usSjviSRv10PhUF/tJcn5SraMp9Et/egnOCeYs
J49xJ8IUFlRGw/so05jRceP9gFh+ugXwrLGHkOuVXUKCcONxCMDv29gEkggbX6ccOyDhbMr4Jhma
CWonpXhlJtskoxiROt6YOW+lEh6yvYybkzPxs2PkcG+4t/XY+7UVum+KET76ciwgPgm/GCptpNgG
+2P6bvDRnLeo4BJhVLcc3UXsfNy/dnAIawCgQYDAgeBeSQ26redEndZV6dZZreh14fUAlW4CanU+
4vWhZGjXhKSNgffBeYwTYrz3uwW40E9bJAhNr0C1ndqbFJ8k/7fKt5WapSwfD05x0h+LseGjbxVU
wBAufs/3dO+zct2GM3ICmeMafwern0ljygR7v2eCAxDDGI1ahLXo1+firkzF4UVQwxzrFAC4mSRR
h0aDzHFFLClrD2wqG4lmMZkn9LM0eevuGocABfYEGxni+cIVluaHtS8KZHm0NC8TlYJrQGwJ0T05
S/+UulVYiwS3mklYzm9zGnKm0hrtshReIU5s6yU+O0ytPEttjimReWeN9Won0dcKtT1rf+QHE0gW
elLuOQabzu9G8dPvopysnDGOcUu5tK+lq+OtvOXw9xLrQyFSwvlPjfnbNfG63QICL64bXM1J0Kgl
f7jgnGiXmH+BgGafwxZ1+BB8hnEezhiWlXf6+7Ba5sVhCczWn5NODxaWQls/O+A3/pHzW8F9oHbw
8XNA3wMx26KYgyXyUFtuhAaGGnrImKXTvDPu9P+DIt6KUQbtmA2OHALdUBtYrxC5R6jjbEhg8r3L
aloeKAeBmZTwAoorkLk8PWwBoH/nue2tJGJ9JLHkYinTjCb9NZHAMzLGHU1gg7SD6eLE2jSfsFoP
q02SzHYvTNOVkBPWsHRYgmhrll50Rz98NCnz1eZl1xwJj5i2y2sc3Zm/9Aa+B6orjMWWvsDGTq8B
4G1bJT5u/L3uja6hfe6k9fYq2RRPlvtJzUyNNmZU6hfy4VFejOwkrv6K0iItJzAEiBU9KTeOmH3+
Nuoa+PA3I9zg4nXu6zxjAxOCRldkarYqmF5GU0G0fIETLd7J56/fvK9OVE19/3JVX6Wf5Q6k4Ix3
of7PPl16JZY/WnxCajdT5Rgo9lAdRcai+1GnlGRzf9de0JJhaJF0Af80b3PSvQzTQlx6w1r49bBe
b/hTG6iB3YWN61vHgL7Cq88eZ2Bnmq/2O8OfEG3HieZUqwJDzxHFsNc7i+Pla90jk//t5ZDx3ax0
50bVhyGlAFCnFJv5T20g9hT8FJjEev52EfFev5AsOfyZOZuxJ/meW/dWfyXfdfZEBjLB4fVNAM2f
EwFFhZeC0AuEVvR/+Io7kSq7+D0WgQs/1IvaRhxXtKZx0aKslIZhUxzlDlbJ4M47re3vuKf6yFYf
va/OhLmXt4lvqbzWKjF98gwtLx8v4VkgFD1E44q2aZAVQ5X+tja7Y7Hm4LcKuBEUvuvjWwb3+M/2
YtQuInrFRpE4GtGKFtUcsHxm+ZpUcZ3jGhFF0jXAFy55I7axW1z0+yzCBToH6mrpQsmOkih5mLzg
GmH45OXJ8rQGmSHtXlCU0HMTRbAxD42dsZ4bdRxQMXpsRufIrPBTvBLq9dpgmVCYroWtFkVyCyEE
Uc+GpvNJY31vN+78F+VLwQKdTiuzcRvipIGb75d58IWN27NXXLQeFPnVYS9E2wtlvssc6/hamXfN
LPXsMt54z/jjmuJljlsIw3VIW+VlNUrj8fDMxGgXiGhT/S/N0GC6yJkp3nFmShL5ot7Sa1LyPPdp
xDqlL+RNGnDnWaRkwn7kB31OnD+qpBRnQSHgNps/oi6Ps80nfMKM6MJ5KB8GHvwpzoF8cmzCZIS/
d6n21RxkTD3OJhHxBTUli0/wVGTTlUGnLQVPVmskgajbFg0q8fAz3xaGLVl3+Xu3uYil6ydnDAQc
JZXp7dAIE/bfaMpurJA9uU06iFMEOKETNjlGLp09qCHm8KMe5IHlYek8fjDgzHlXzu5dIGrCQF+2
nCKXa9HNO+1g/x4dF7ql+byWRe6S7fUicFMIaHTdwo+IlOERZTbb0f7v3XD+hhOBqYl6jXbRTIFW
ey+8KZ8hVG5X0GCBXpP4YwmfOpDsTBTqldxsomaggCSJkud749RcWHJOLT1N4/IwrUs73yuXuojj
WMk36br9osF2PXHJqQDTFZZ200O7PFGF5enWSJzpe1BVkH2QhdFyxReQ3CWG2CsWs1HzfcyezHBL
MyiI8Vp+xOKEfU/Yr4enjhYehqlJiZ1sk+XLAG+fxY32ae7Jg71/HLpy560XJYSzWVwlICFLEdkR
lxAUT55NC6P1zvTsCDGbSyE394PntgafqawOXMMd1MPd0MlF1mrVO4jAW6h5nhJWsJj9lKQGkz88
QmGulSyh9/SzPIKadnnUqflzwaIr9KWWg3SBv/lI22qtDeEx3SW9kM9D99Bv+5pOgJcPlJ3uG47w
FSEWPpktdFJssuRu3uJopVZdIDr+UiCu85zPxEE/AjH1cfYcgSuDjxTCBPs93F/zqyzfUESddfkk
e5bV/mns5VyanMpVhCmTeiCbVkv/wTpjAGGKgX2JmcBrMU0VPzfnQrzFoCYJ0pvYiP8GtkRYtEKu
qpTHBr7kB2iCTjwkqgdOLzhcQzVKC7HG4dKANCfospyDuTOmkI8hBt+dLdg60Kq0yxXJYbGfXSna
f+u45dsH1jWZB4DMIa8DygHWNUCdkR0B8j/mKSRKMIOaoSNsmjeLKVex3WqQV9zqabj9FdUajr7m
K/z0StXA9eVqzvV/zd2VO/+pyva73mvZLBThrJMZUwTYn055uzxxK+Jvb4QloTZ8RN01BhcRf71A
DcEwy3bHGx1VtNUtgOWgU1ciNjIEZAHfdLQnRERY36ycsVu0pSKwGMtVQlwAVMX8WatcOZN2V9/s
YHoP1QJ8WJnnohPah6EVk8gUjGTXq9Rfu0MolxRCv32Q4Ubbg0ZIaIlMlt6s98DKU+L+dvnjaPH3
eE+N2lz60/nnbeZXA7QoRzJsHW8y4UF/uAD6HKsDo4G687eT+OtU0BAWYC+EQ/yhE1afSPj5DYdI
cEijHOBB7ExoAaCzv7W4O88xhZUsLMiaceWfb3+eWECAEZOJNOznv5qqs9qUFWFgT9vb51f6GmXH
HQjiz+s6e+2T3VZByM5jWxOLx/4BFHobuFiCOokkDrn5J1DJA00d/bwWlW73SWYuFjL0KcDrPUnJ
qBe2svDMUEIoA31v7+Ww0UDexgwOAi/he+JUIUt+5MZvoQmHUDieSysA22MRt8xBbmaYAylGNZPL
PElakk2bDjEwEhYKEQaPEXwElo9qNl/8Q0IQaYhRImORgfBU11Tbat4WTFwyjK+Qnn9pJtyfSaKV
VEPFTILIVPtVWynTqSp/dGCMzR0X+H/PEXLVBHpyr39AwVxQ/lrgHvOYcLqvRy2z9nAxT92iBJB1
U+tm7hZ0dkXDWEAjrOdmUUKikqRk4dEink3vgohkfwaXuMLXQbos1z6LmIe9U19qN6oYXB3KP9qR
IhBB6cg2CqXP7b0hbda6Q7Evy6hF1BhzuBJXnms4OWO9fvDqqW+00WIDUpqTQB9jPoocAtm665g4
XpOI9HW/g0hiLn0aEpDdjxI6qdAjpbrWwimHE0AjCF2mhov6dRelcNMRIZ3gwMh/c+5FZCdFXD4E
MRccsSn5DwaUnCcQr88rRN/RsWMMlmpaP/yunv4060yjxANrTiXtAv/AkFfyJkrYQ1l7iCrRai36
FnxLbWP99EQ8G8FLb1kP0tgf20cJXF392lIVHD5ST6aPIQwy8umdSvQQ1DNkJ32YgkrAROXeTeA9
BqGFMdOMIu88OBsoZchfXSTN09nJURoSVVvBIyygIVhIC5gROkF8tKnBz5rSiAFJZv0haF4zvX9I
QYJJeqHlaOq01lsmxn8T+JiRAaRd00moYJbnl9l/9RJcIop8qQDfwR5Bwl1WEBc1pH+GHgt1Hswl
Hb1YMgIgtns3ozNvVLnsg/mgoBUBVwX4tDC/w+8N/zs8tasOBegVCr/g+aKMz2RkKjZmaVOagN/X
0LEU5OV6outYWlAlqhQNa2Kk9BEWTSY1Czx7lXFvAcxqo0RCQQS1sYY4++i1ajJMFrmnT3hMMG82
nNaN0R1vyBaUjuSGI1DudhBZI7Ee/v6saozve/tsn2oRJqAQE7PaOO39sVCgPBReebpSuojhSHxj
Pn/1A1tFvS/P4zvhXufXZhKX/7QEk/lSiYZAt1Ro9pM7Rr8xH1kVIVZnKDD2A/msQXHj4jjAyia2
qioylmpXHGZB2OSoklia9FPE4yry0w53WL1EiYhB0IO0gpM3sfBH7dz+e220VxcXOuJC4eADFBDL
dOOGSpwd2HE3pTUOWeC/o1TgMR7AtOTUwunqmRijRKaWKulvSj3lT5qoKGkgJzY9BCQzFaq39Nl6
xTGe6crb2bXhczr3FzRuswROUaaj/7g4j6tToqI38NKgjDQ0p5y+9BDPe+d6dYp/St/zB2EoLEou
LXQnzJi50MjehC2+0nP56/ta9OGrcz9ZUYiprGHnhQcbspKKpKPYxZ40wueEq12rE/X0BUiIlWOc
LDlWzkxJtlaRekSa0gK8dOburWtPwFp+/IYmPNamXFvTmV9qPpGC1A6T+m9y0bCj6SNPXAtHmRLG
aRYaQ2QCGGLh9KmSQWnkhEJO6OqbWFgxF8XPRk8HGe3ftPdRb+3mxTmH8NH5XreDBzLxLm5Zi4PZ
h06Sv6zZVbPDTEzfC2kbjHgOYEp0LuB6L3NDZ/8d10uUuC6st90hEMfLkC3951gj9g6X6iMUebii
LCSu3CXTIs/RorLLi1TvDREs4s3tc+5BQf1R6l6pAfVC+wG42gMAW2fIDcpPPyM5RxP7B7O7mK1l
yN/6tw37ZvnJRA1GzobkZgGdBGvfXQ9t618xC9h2sj1aXXx9DMh/Ru98a9IGBQyfXGrWpcqgxH2P
4GqE3AKvxkXKG+kNuDCr8IKuvnjJwTojqaEGfCR0qQMqtbUF4dWAtKQvLlfyedTSqrQ38dAncYgH
FWyqlKxBcWzee1KSbhRnNoNjgPwBc/diyOqMjojKpMHzjqwwAF/B/N9nY5Gn+t+SWoRyhF3Tt//I
/RlimhN19bc5iaLQBMUcTD2+MaWvpIpkBOfgqGWFomYNSBehCatHC9rrWV3q+fcjFCH8lbZxqsH8
kuedg4+Y2qXAnC+jsMfvjcMc9BWB38i8C01AHydcrG7VzVtMJq1VDIcxGwuvJ+UUNeJdk/LKOzcC
rnHXci3iPszP2wqZvyxCA85axNY67QUJCfCeFRihxsIR1pgFl76aKoJ4uMxi66qqrG7ruH5B+nm6
G93/07fQsgcfGTIYNKW9ZH8W+KV5xH+suZEYHjaMDQ0Qyzs5OzWbtg6zYLwy1kzyX9gHKuTxO3OP
JMjp4QU+/0iBTb6Fp4OzMlqoF8gQDa79LM8MSc32qWhIwVwRtyiLW+PNY0jnAo15sPyZJ/u9zYHd
VRTDRN7QNzdyOS/LiNViXYbdkAw47H2WX07XBZmfzfNXGTQOgGtgLxaNThc9Z+bM+SacCX4Q+Q25
BPkM4S3PXtLodBtFcOJR+Co0oSm0nyXkg/uSksiX6TWgHS8ugNfZnxLMARioh9fQcf8RRBi1U15l
mTiwPK/th3Os8ndJJ4LORqGtJEzAxUTzHEFtxi/ff9/qvbpC3winmIcVGLytKyE/1xwJu/lsxt8D
4vEky8O+U4HpVSsDwZy3jym3r3i5RqVThwW8p0OO20arxmrG1EqYtqqWqr0teoGpiVkYRpf1Ou4O
YLiQFJ2hCRAeJZ5m7iLB69FJJMUuKbMsEU96IfYAU+bAeFxTV5LdoNM972xI9gcXXGG8gsrrwbVi
Ra0VqTVCr03EO3Y/OJS32fpn9MArTQv2q+EoqN/f+1zsEENlLSi+RHUaRWZ04wAys9ePj++IEr9l
RoOtKf9wa8vCH0qj3V6x1k4vFWlB39K+A0ejJx6Vw5mxKh/fR58msaYnp+qjHyUj8iv4RtYoAiKv
VpcBJEv+GUdIQOlk42uFLoyLoksRXHwiny6BSkdON65ru23suPMY/4zzOCNY/2c+pRhEF6+t1eUu
nu8rUeOK8oxuTGivJfVTwoc9O8AGs4f3epkcXrRChAfkRGDrO7C5/a3os8PwMPvoomkL9CMFdf36
4z5XSkDiX2aGYQu9gq/392e2I549MiRFOSBcgg7CIs4KZCgI5478zPoRjAzX10SAAtzku5Foqq4U
0Haf/JW5WNHFBlasQZyhpLf3cIKWRCe5kIiRgb9BACzVOWh4xZorEgwYdChYv/YZ84880CBRjamx
rSUCGAsDvwnazxj4oImvU+7LjMtbFyYYw+mP4wJO3S6sPlwKnaZshDFSYVvWZMo+zeGM7+ouVl6f
BGaXDeT8q2iZaiWkLo+qnXMxrS1YyGwYWKVlHhyLpOKxLhX7incfxRcVFHmsMXqySe8ZzEHEQcCJ
GE03J2wmcG3E/PWWGsBX1b4VfTtUNWNJLUoMmkeXovtIySq/OchqGK89BVPBpkmPYBWRqFRC8sOJ
Srsle2C0HMRYjFZOaAJHyxkDljkIamUWaOX/QUxezpGhWnOECLC/WIoI5ftpiWyoTlIDF2wfxC/R
SbgTYsrs8FHQFjxgxN0ODrTcMXjhYiWLpd4SqMRacE9DqA8UNuoqbBJHjWY6ydFsTUT9EmqywFuH
2mImRq7jlLtkAcc7Yf7+f44YjTjAYE+E5Ceqg1de1IXu9E/MCGuRB+VvdlTJfMH48XzwssQrFvb6
bRer/8RYjoWjdH4MSYhlfeI3inVgMNkqz16Wh6GAva7PALjRPkuUzyvxHzzSCAfge9YEqAPQb0t8
2E6+t+5h5iOPYAOJvUnItD/cVaaBWiDLVw1yCJipBjAOCyy6zwKnODkGsPHBb6nxkCY9rlcr8DjC
Lbg1FEFCFsdlSxbK1xBXNBJ7tHBq4Y+RKjAcE8lkqjSBDbJ7j1NI0hQ5NX4ISgHbAunHdpEU29fY
kwWDmWU/mtUPvJrtZrWu2dE1I6OuyDZUWhmRlgml1MabWrHQ7VCTSGRYxmMtX0ZgzkaLiD9LhaMJ
CrLqMMArB3tNqcSWCJIY8nynXwe3nO5J0sa99R1VVucW8YVVR53X1BeBNRNf5EF3FO/8P7VFqjjf
dEmd7RRi8W5yRN96oXyPep+zDLPK5PRigKuRavZrHNgdwh+OhjYr9AWsfSgLnMeB9fILXMIzP82P
CqAbhuzuRfmQYBa3/3r017HZIjdkIJJZ2Cv92V4GT4+jkv3c2gDYIz5gcVuoYNVyzJlwtpxzm//h
mSeqaB0XHNosKydARVZE9G2rsHEoXuDSytGt99jLAbUp8phlrG9AthRqxHEvNyIaDZ6Nh+PKYsr6
mVh6na/HqctQp3/GhvgYrCSUivFQxpIwKngJewIocDiZe/ycVY7u4QEfqUorj7R7MYvb8sG+KWBH
4vnI8CHzR0sIJUjMNMg6oeQJzRCjNRLO0PJuoxFAcBjU3aSA/fQQg+cK4YFrRU+OW6E3LHJkHO+/
oXqj7YwcJD9kcy0VYoq1+H+7wo/ZmitlV+MCkletim1paU9XrVUIkfZYOx+CmBuk+iT7AEVn28RY
vwrOesbtd/A1YleoaCoD+sZX+C9cBGnQ0qVu4/NdqpKMr0QoaZuvo2w2uNmje2SeAiZKqc04hDQt
gfe+Q1unTrCJQ1bSTV2dc1whwMhEmnvtLqe/m1MESI4NjXjkKlnpFv5ZNt5wPdFed+B+W/ebuqJ6
1vznDAFCUgltFf88AIZRq+xsTaTQx2nk17dJIYPoQntLM0pV27chn30r4qWzKudaqQY5B2047oZH
ZknMtDXs+RYo7jNtcEoJMbNwMn9xWE0gy+7kGGIcg32hLyObbNBp+hU4ODw6HTnZ3gUfPit2Vn1E
xPN4d5+PlThp+XOc2RelVNUYUCbsyoEYH3Y9gp3OdtPuiOSD76VymKSkZqrWSbB+mbDVWzuguyVv
S+n1UCJ/Zcb/CPIBas2bBpQHLt0j7MKXofgDnX0gUpd+80U6W6/Kf+YIHHfKygyDZESCilkl0khR
J22b7N6tFIhtTrUEF4ot5wkafwVpa/bw6TlfMuO2DLf5+JJH8d+ubr5Ly0zMKrLbNdMTiOJN24NA
MNbX4Cvl6al23LmcpEstSzR92iZYBP0/LSGdhUP5jhAktoF8IOujkJiq1cEw0Y4QmCwJjMwTcJ3b
UgU4ZZ3HPPC+PTh5PnnGNXmdGyWQ6aZriRKbpoXjxQXMz1hHy+6cXxc7VoFypg8neQHSGOA4nNHW
nktd/dkMKdzQU+pYhYzAFb+Oj/UZs6YPnG3C70/kWbUOTgQTWP2ea7XqptvHGPvo5QaIduWQPXbJ
svAFozIHt+y6fhh5zU6sJ5bsBpIFZJuNUkVBIwa1PZ0OlqO1kHuoT7Nhd1YdxAcCnBwWY0mAIYi6
hERAkZBbX5dfqUG+8sv4+XU6AE15bC9CCfIhcOoojKFwmVS7zB6mExgrrQSHmMJIjfumdqmXaTia
LhncRokWxVdaIqnKyw6boao/Ti8ouMPfxbRPFrZ75sdnJkcywZq2OKxBvDVySt4sUgr46SmAFfKG
Z7kydkYbb655LF6bG0iXemnmmHR5R28TFGsuJmdiNHurTkktkBcOcX6NKqgXrKBHnEF9r0wmQ+Og
316frSvupuxJr93EznRvc223+utY9g8tlTe2HP2WTS8dZtWpftO0eN4oxyO6nMLiRK2mkaG4e3Vx
kZC2AUcPpgFiTSGYCEmIUgyD41GcYK8sTQtkThzUjjoedI8aiLhf754RNNWQYr/9bbN7VwsgPwsh
FVPPX3kkyt9fufwDUmZEfnJewSdZeoRlIFze/kmouW/78nTWTbX4n9xLeezLTKYZ7746yjaeDqUJ
h7lx/8G0830wf4BNUrjUgHbo7F1DkVr+KmV2fidFMiyaVWrYMls4u+bADQzZ42ATxrUNXgIjFJtZ
Bp9YbBWsuuDQ3j1e+ziWtb4dPS/jb8snG27bGvrsXugLf5K7WFZv449DxtdhAde4lH9F8I3xL3eu
OVNa13NmB+brZYb0lRv6QDyV8pIMjoK6vdPe7x9Ce9VLXtHxDrb/W6BS6ifGc47y+gVCR+CLl5p8
uX3mxXsmlfvC0kqHZ9PuzxKDALEzLPLhCxocWBec9iJfHZzgs2mUJwcStfg2CyN5pd2zHVv4za1p
06Y4DFK8r1+TFeWKwORsmwqfQV+jBjiWeeDOE2X2fk9FC71xQj/Yi5OQjbBbVdgE1fucNRsRgnLF
NYwJycN0HfAgymgBX1FcoAfYqR/4u7CQtZl5LS9eHQR8CBPXRih6F5UV0NNaaRx4gldYi/RmZRWP
oDXoczpCiLRryVIDbnQH5csy2clOB5+iFdNTvk2ntR1jnCIq6bQFtEVbn4iiUD2nyfN/Lhex0Kcz
1ehsL9vlqMlBVucldIZYGSfxU1tqSJT7xoWO/qBYPCmah0XjMCfp34fecCus09apq+65B6l5xpxP
cp2j7lNSHbP69tjZtBaL8hJARlYCeoUty3kIOe5V/PX14EZRwyo3fTvIydDZxAqkBqFpsBPUa5uu
KpLdiML0qGo2S42+F/554KIYhJWgZsvZghYG/sbNc5zTB1ls5M6J7dLrcS6JX6KKM1cZAatD2eha
brV5Oa+rNrURawiMFlTda9rfRY7YNINJjgnozWepWB7iO1pDlfvXrihvD4ZlGUTgmSlw/xAcLO/5
MY3m7APbNp4wLcg2LNgLoEjSt37HdqSp3ZhxXRAOsOS61rpKp1+w37IoVhzjLxkuRo2IdwJqwj/4
8rP5WOdVz7Wf4TZuTH0hafF1jjp0s2tiXH+tNoQndXYW0kAqu/hH+6zo3KExnYLOhUrGRZI+xpEo
AUmAlYgYHX4ozCqrG831xaDnekm3BlKSHOcox7Dk1Roi/lhrup7T++T68qkCUvQcFxB2nHn9W6wE
q43yTidXdPBVmi5VIvLxV/UhpRGlCH8Y8TVQiZA0hGHbeRqkcsuy4MIHpD9KLvMlDkWnjli04e/q
xMqA1axWsLVASZUapF0aM8HLRXpjHDeb3R1IzDhpgGuexixgFDu/3bygickXE/YfXh3L1ixYtuCl
7hL/gFEKB6SR7N/MJd5nYJRiSjscbjwIQ2YifMR6vUBXhb8GtGXO6CpQhfl6mbeAqUQpVRsb+Bsf
IQwao/MJimj5bPmQ2JOM2/k1EIJRLG8Nf0eOvXmPB24xh45YZKqqyahxO9d9IIorTH9+l7k8tSir
ReWTsq3/A+0hcbgymLjQHMcLlmZoPNEcC/phUO34wj+0rqGDj4F0imBZSzrQDTIuXiMB8+2iRDX9
y/HIJLv3AZNtc96q+TZYGaZeGJjrtg748B+G0u9yIAu5bqQW2sKb81NBpRZ5o8XrIUBguUHmESVT
Ky4F470J3fFrl8NT6TPVsbHpOrw5kNX2Si/pJnyzp1f249c2cfe13bpHeT0+Cu+YMqi1cHfcvYLq
q3DbAHA2b+Cg8Nd2qCB5NtUA4/CxMcna7kC49iXvrm0PW9bjWA6F8pZ1En8Ab+ZU1ZPuBbP8dgs0
0pGx6S/hN3GXwVLAHYokMxwYl52+FkR3IvcxZmAlkBLQlUlxkX4HXhLm7k4ApTJXzZS8b++8uS22
1CrUQe2S2mpvVxA2aLQPE62SK2k8l8oD+HE9PwhSFY64FT+GGmmx179iR825/EXDbpBpNmug0aT3
ji/wr6S+WvR1R1AwF09dh7xLuSg26d9UoW6vOTROcD4aJXbi8pA2AieiJ4hdiERqsJ5aa4q1JCcX
rsffpspuq6ik3auwPXuodL9DCT2b1y2MBeT/o3Bh7KydoKaTu4e01e64T+uVirhe3okrKGBthm+B
UhwIdKPAVIC76IWi4FAsD+Yzs/wdYCfw+Kw0ES91rA363wTNoaghKTVdrZk5V6O0++HEUcbUPaIJ
RZc5VSUt99YcxzYqgV+EChG9m4OZ/1Xz0t52//k8LEORTjSIn5EUW2ppDNP8VZ7gZf4cY3AxJdJK
HwxHtIbD9aGIyML2ECSwOPOTz0wOmFQCmdRRP9yy6rz7svu8iYTLq8wvp7Zqrv5AJzCA9mMkXSY8
036lVLmuUAwQuCycjiSHxNacMWREzZQHZL/iQflzK3c1Dl7hucJE2SPdoMHViwlmDNwCgygkMo8c
dKoKGYAcPNro9u+d3xJHZ+dHcKLl9gtYREWKpjqwxxPJN2CzQLkUolnolVoyjxSnoJkgAJdGNCnA
/WJJOLBqfk+qHyYU46G4lMy7F1THSJKm+zG4UAQHNO0fho8Zw62CP4wbYJ4HiySNqsBo8HHAxvp+
bM3AeS+yvK2ZuKdnGNTvYFA/v3loPQRBaVLcSJk1Vf+DpxMdDhuvy+QjUqcW1VLPeDtwMMlcKmaX
2oij1QBGmGPkRnY66glpbJF3y+6ayAkbL+AECrQFNQm2mbPVYEXafKdR+5ugOWIUhGvLIPVqOcvo
er28EeYy3d9janRB5PORcu9wVYwygKyIfaZc55Y7ytlWIcbscPG8jkxvcU8M+3VCmQpOfxVf9G04
4UF8QHmka/roIs9pWPt/V8UtzAVbMRZFzX0NYdbTUEISXEOU9gb3U363FJjAvA34OlvMKyV/Ga9a
CkNZxQlDq+SCen4OR8W04ZYRFrjtw6tmOnE/4rluaGdb7+agIJTNdBREqnDB4MpPdbTi13fX1wsL
PELLWS2mIc4iPInKlUZ8xo9n28xTX41nTA46ZsKQk1BX8sF7HejT+s4rOJs754v3Js+x9wrqr3S6
R+2SC+dmcsWiH+Oeqk+xe9b/ztAmcJHBJh2AhHSm6QSoAG+X+cvVZ+/pUu0FCj0vHqXtRn6UcGHw
rpkxfysd2GpjlivERbOe6F7ytRTrzakeaKyufCxBrDldxkCnqJl34RNUXFgjhh0+2nX+STdARtGX
Oio+jeKrQdylMrFdbyXjv9/OB+13IEr9NBFxA/aShBcXGs64g+Ni57EdZc3PzMnNqcIpqGrkVfKr
1SX8zXL7gtXmHo6BckzVGY/yY/G91yv5k/ME3BOVtxFvP8s+Bg7oDtOSeCYe2jMI8SeQwbW59BMk
Rf5N7vbY+JqaikTKnznuu704wFAcOvE5Zj1sA/2mehRMwDbECwNeKe1jONXXCs5KFO0l2otUuvYM
nv7Xdi4PiwVM4FnMGUGlGFwKMMsd1byJWsXxHGk+oEPqyYjOxGmL/Jsgi2VQ4ERn7Zwe5ItjIuqD
+hWVP4Q9BXdf9fQi/Lb3Hr9zdms9m4fzfZa8Wn/y/g3CBi8d9QszEOUmv4ojNnGcFucGOllYv7AN
sAUJQ0lFXHy8Izh692nGzJcQe39ngLVB4JWb5Wn4kNVZ3muHyGqid8RlzvOUS0fbJArRApEW5RIl
9bw6BRJYOqgASCj8IZBRTYTeVdPF7k6nHSWpb1iBvc9+Ef1Yy78w5FTbJNFdKfDxHYZWI9DlsCzW
dDcSMerUDN+dkMOwaKtXd5sSd+IrppBkSrYN1qoLDPO9HW+a5/5n9sCWNQtm4/6aZ3z/eKWh5K0c
GYmQYQclmfLIRKXFHjzc9sITKh/f0Qgx8mKKLIKakWbTsetGeBFkL+sa8YdyHM5m66ZalAv1Fr0H
TqxEeG7o+oQsE0i8KLotzuUXraT9OBGUBcD0HI9n7qfud67JyIe9zRiweETob+lVjDYZn137zgjm
GNNNP71AtGs2v136ywqFtecHItwvO9vBt4v7e3FO0g8d6tzFN1ivWjrh2CF/pbp+zMehBHI0x3r7
j5vbZjsJKpZCGgMWmF8RRTyhHCwzG177/c4byEk5o5NcL3chLqBSvKk00zYrg34M+PAcZt7zWDH0
gOOjyRscKN8FuWEW7JDSRlsEweq50/27KPPfnI8e+Pagol0Po6cf7sBnm1/am+QFs0Uj9KDZHwXF
QV1Qg4if+muQXyhRhO5HZgYo78YYnTb0QYJoJlhyOpSioJfWfjt96js2MIfLUgHGkMoAYkL+cGbI
b6oDkYNV/dknVkMBzmKvmH2Y5+Yo4uTcLI07QfDVRsjAS+k7NvCXWsC3QnnpfKlMbbcZI75RUiaz
TQ/K1ZeLq5XugEyp2Od6jlEF/aiVtBTVtmNaHkrAJx6q3SjSQepLRcwb6x2kTGnncmaPUpi0e4je
Ylmtxy/vEkN1BLJ44zPXa3sx+w7GMjys+Tt52rXb3tet1QmXbcj74sHFzDHlUtdq62Sp9CtTWeDW
RBP73vcvBRE8AOcQXk821kqbojZLomI7WEGpjjbpofyqMLqpmHiPee1ASy5cnvTQsAkCvCVbZ2K1
mT4TdrvmvAzc406rV0HInS/pVi2pvfnMg9ROvU4Wxcv3VC5Yy2yocqHuZdhN68HP+SFyTUdH45Mf
a+neB8BWvAbQYj2sNpMCyYVvdo+IF5VeBrnhCXrseOtac+7dbTqSnCg7p1skT1ZpgBPVU0HOQ2HQ
dfocZJ9RORC9Wfl8PDWDSq030ASGHWDguM+VajW598Xo4cf/jVJI86G1Zcd9l3caLjKR2UJXuhp4
6+CrJ6M4Bfvhaguo5v7O6GgVsMvARRKXlEsUJ1hC6v7iKXtP76+C3ghzZqMjLm0n17lbXa2XCypC
C8+7B2Ws1Lpq5pSI6ItV/mgb8inJ282Nl6Y2xYzRTkfQjnIaf5/dP1tQaG51EQmM+MdnGfkMn8Rc
xFVFUZYl5GNqaLjWsyWKCJfyZ18GPMIdwXs0Qd6vPg9Pnuem7pEyKr/8uHJAoTpZUwTQdBLmZQWT
gHd3MLl2uULACSJesDtBJ/hXxBhT+qnJ2pSmAh3AuKm53mxk8RfhfjMpiah4aFujTllIA/Pt/d4h
gdPULXDK3GQd0qvAUNWRMEWanSLi326lFTjeBzFVFBu2mpPE97CJPPfy1+85F1YVwe8z+xv4A1mp
z4UVOOZdC4/q88fQ5G3q8esftMO90zq9cConlr55DrL6KjJ1ujYh9B5gy7RNIvDtsBPwYVrtSVXH
wtUZ1EIE4LrnCN4e9TcxoRry2zQxbrcn6VAjn2hxkLsKuKUaZjUqUGlZghPMWof6jKzShPmYTt9R
8uLIaMAZYiHb08CoBv3SdGew0XlKA2M/8rvZRYKP3iLM+PvQRwQVHUFKOWwt6LAX2ZgPnU4/RxzP
XdxEhfjGZ0lyxhayXXX3bQS3DpiAOS/76WU2Hz8O7C3pNz7NNhX5a4LwqWuWjkwk9QZD87Mmkt+1
Ui/EuNrPUIys6hvdgAN9EnwGRCEXlHSVwNC1OKBcwMtKBQKmvqnSljJzTbGSOY/bFC9rtnrGdAPE
zl6pEySfo8fOeZLIUwGSw7fzOYBdJOFN2bNW+n9G3lHpip4JMCAoLsXe9KyM6WM36jRcuUSrKHAa
Zh9PNBXXTRRlC8byBdPHDJ5jfbm1s9gMayJbcxu3W8R4iSLuRc5JAFze5caSE+aX9KXCu6pSYDBQ
crHdzeDIQWJr/rqJJc1+eq2rS+1QimAM4Qc36he2+M/7Aiutq+ODOmnh4zHNgK6ydXMc904K4J7h
7QvGUQncaaE1erpR0hx66QwW468zyz/MlBW2plaXj57sqI8Q48r0ys9RtMiDUJ1l3AMm5BbM3u15
sZOB34H6GB8m+60ivUMIFQSCxrIpPaDmIBDqKf9Y9GAXkgkrKn4ina1ZN1X+kNMb7X4lRpIDGhqp
XEfqMUjCoNrNs8VNawvTb6w8bpttQ4DGxkzI+BOPSMx+2TerO3QkzpnVDN6bWjg1jXvf6J3utmv0
bQbQubEcd++onysrIoJFqRFYw4Aa0OShc7Se/KLjfvQgHwRNM5gM9BXkkUGWLPxJqpBzNATH5C77
JjOFLbYieg3JRWYyxByMIMlP/BM2MXBgeRjOycq0ERvlPMweIiRYHAkPhXRoUFBXGV/4yAtIJpdt
Yz2KMCS0mpfCs4GzzJbfc60w2vTbbd1irebCKHqNcC2bMNNZvobrzXVM0+/fdgbt2ihKgtXOOOTI
IytAMvRKDittZXG+3wzvY9wbzEIjBQ1CjlXeM4aucQZKq1SdNwzKMvh6LjNez2qgMFFKNk8XybH7
bDs4KPJaFobrP6iSq2V4ZyyWdUexNxWsZB800yWDdnSdN4kvHg1K6AliBk/XRgpZM6YCOAYenmG5
xjlsGnaZmhoHOYLn8/ClS9RYr6ZrktBc0KN316iPGHLeJWDWedGziQIZiIE1f+/LdUKG+03OAD5u
O/3mFxy1NYzEvAGaIufW7TNVMJfES7w8C5ruT8SibXIYvLpsVt+jOWb5M1Mmf+4WsRBm+wo1bGWz
iD354RisbxJNfwGengTAuc8FhMOSJAx0BnwCSEcT8E9KSa0bHPU/VcBdE75UXwH4x5K1mhTseQA9
DuyM/HD97H9fZqS01/a8HNy+lUU5W2/2s/Q8e1xbtN7Y87rROZ254Gf7uzcSMJXk/ZjsvfXZYNM8
Fl+/U0SQyqvZ/mGHnS2Tc3QuuQRzjiBIwotTVajyyJlhlGZziJtO6VPY6mQlxjOf+EVgYdmI27Lt
5nvFkRuOtravM0C1dEpkm/AVDs6F1DPGIezQieRvE74IMXVrxJyJiqvduhOe5JlmlX/vnQEJm2z/
Ock35PQ8K1wjAAQzzVl2Tti0utgmtYY4XKGFUCHN/BVKi+h4J59jI8AlsqG8Jfw0AhM4gD2J2Omz
uJw61GFWVdfkdVaIF1jnCPde417IWeJMCdx6K0lJcnGis2P+gd//FI6IMlIaAUdbYvy7nS7tJhCl
uVYH4KrVPvPcvd5XxIvnNqIU50BElnYrSfsiyY5DRiQiCORKmTB/Od39S6gRhZq33yYLAeMkj4jp
DlKmBfn9uCK5QNvgpgRvSeGLMVae49Z6tFyj2tWEKeoxT9ctpgCGNgu8heg8CGP3wlYjWUVLtpyb
qynvTt7yj+Vp3CnZYrbjP3ksF3u9HeK7m1viOUONCbL76+7VEbjqR2B4TR2xoJ8LljfQTQNjfVH5
m7EvsYWmbPFd4bgq9q8q0t1q+TjZIasl66IbBGqt865s3WADvyQdLfCSUOJjKhNadrKQafOxIyR6
v+Yu0lldYGNyHgF4KXzpJn+bDgd6fZ/UzH8JYka9ReIKb4dTRYBf8ITY2oIrMvnP/JIY0WPdy7u2
d2C2zT4HbZ854BufyACnTPFYujrgLcCZaEs34nMzzrCj36r8ga4wk0KG0n9NizUBl1J8c7sawLY6
ofKaFuC0Uo5hEe+GDypE9hZQZZG8WptrEzUYs/eKeqemZDqIlF2pBvBtTkRMBbcGN1woq/ZOhpiH
+ddi9nBtltnAYSFTU///vDFksS4B4MtRSJoDsd6Bzb8XGO6HGFBoROG/baOadu0vsEN6jGPwI7zE
EausPRbas5Vt/iA7L+mPL0fJjQ1cvLVP+Yyx4hDkAKI4pWWpZjeM8SxA0rbfqegGLxDut/5D8wKR
zUImqAm+A3tprKQXLFpKGZRxfL+pHSdOomE8wNF+ZsM0k1vXyVmJ2N1g2WE6xEKgVTvdXsfo0IyZ
xXt6rxYaJIdkPgVk24GbfydwLO+ICft2VGoJoeRvvQoKmMtgvh/FYprf8a8UFw6l+4nWcgOxxEoH
5xIYsTJ9Exwo8kptxmKHPtZgzKBZ8myV8MlTOdE4FeFWKdLJd217zWD5lNBZU6xcC2apKNKrWPdD
1o/wHloJjml4/dE+IyR97lKodcc84uhO6seJplQnZHn1qdpQVVEoTO0vYUzkWL9GiCYrhRbu5ymz
K+YK4pDimP+DokhgwAH33ncCkwbVlOOCzpaGh30X69MZOF9CMUsZZQCVMGWr2glNAapyDd1qR0Om
uf0PL/b1Hd5hBDA1pHloqfnur8DRmByo7IATtZL6A/7+SsJhpRCOfLWHZaqUyGZK4FEZlcCxqcj7
8nhIwyCyW5n8rkR/c9vnPC7HgV2v7DrA+egpiPbL7aI3NnsYTmAcpjv5xGtrm+tKdfhOA6pjJdfX
gBANC1fJCpJxZmTRoFPCyB3PN0lOw+NXT91uJXldLRhOjRmoLY4lhcbuT5zTVW46jZFCaiGtfsGB
Mcd3VFLmd5EXo/NCWKXqO9hMkY+xQGdhGB50WSt0LDwPfNR8fdNEHcoRjp8TzZ0agFUsMx8p5MAY
Gw8O7IRnX/cGRM0a7B9yOwZvqmy84u5SFJSwKxGwwrnsGHV70e3rCUeP53n6HJm3hNyBYaA+PhPl
yGXY0gNIktrv3UAIzJuY3OK2Ons7uXn8T+v1GYaxNHIeypDrei89epicb/GiY9iIoR+8Z0JFSMQg
mTZ3quh89879oWNVExei9vZG2fQyylqK+1YWCqIQztNR8U3tWGxS9Fj/Al0pQHbIOjvs2/tHB7u/
HP8FfFh93CMzQ4nZ+rE4wGWqBmTQsLFSPKq8Dq4I6zjGg9cSyy33I2e93ZDlWuTVCEyMk6JE8OxU
pxt5+d/pxbz3x4GzOawd6aFcpg/kZuthwgdlL6I7DBkwCN/k1J1Tb6vFXAD6MyVVn1N4lg11xcEa
qjX4npIw/kcE/mACm03pCw5HbjOCngXQfX50X/CyFdsXe4tJk3CMtVos7oETr36URVR/mZfKakct
taGwBBkP65oU6YPS+W+a2qz/ILTYzMRpDUWtOdvxyUpkor2lSdK0HljgZxZc1bmZzyV0haqaMBDw
5BBOjaarUP3kHvcn/puMKOThc5Uie4Yjiv/siYVhJ+l/Gu4hzALSZmKQ89qRJIBHOSpBZylh4fGZ
Io7ZyqWVjmZ+h/z9YNZVlAf6RQI+oTLIJi/rwhcxXwChUWBzR3RqEF+UjM6ymzy/ygDYuAmnEIrO
gBDNW0IH75noLzUIVASYuECiiJXRGkskHCw9o9Z5G89pUdMtjvsGk4DvH+emYcR4g7OYIKmZukW1
wDVuleqVX9Ll3NfZ/vYeiY+rQmUA1C6UJg+lszqwFsAUDDTSGnRL2CKEdytGZ53SvN9UrZiqpKg2
lzc6UkaXquogLeIzkbYhZyXC2vm1VXiIATK/Vi9UARMKWOsDIQJ3K9yWXQH7uSB8Vk1Cf1cRXAPO
nqFpChYefFESZsS/Y0H7XLmVlTh9NjIAUIwGfVluU9pwVjt2P5/6nmcc9v3KvOIm0ZqrCDyTVS80
pMG+Goh6vldEtbzxzHjAAGpTVnjybgVsP4PHKPExznjgMlAQ1wMbG7FxPgOXgxVg75HqwRqXnq6V
hifoPMQ4lDKXW9f2Dq3G9thhyA2vIfMyQBnT4Gs0+whCQ6DRQkre6i0jwHDSpinyRqWuPwhUU0Gg
UhacAeFXaehWafx5B+sMtSC67US69xkrcWcjjYzFIh/j8393eil225xkdAbYZ7yPxd9JKN7Vg0pF
8JRiOJ778jeopVAsPcz+L0dINvPwpML54IBCSNzajt/dbTvXw2BbrKcNMgsYWKl1+9nwkiEceUcL
rYqunW4P8yGbugXOwz+U3sMPIhaY2L0aR0n8Mf93FDG/6M8rQVevS8JTy4H/LG7jp75YCX0YHqfd
/Dpuuf6KDkfVDJY2qlOdPuu8jWmb44WXzyCV4de7M5tP2Da+Xm8/jTLHRPts7K1CTKrE+nhhssY5
onxAJAACGW51lsJGKt0eyHJ0s3U24xhCaRikzPibj46vHX3clMmuv92T2mu1OOgq8+XF9+20wkcG
SyNACujIlFus/PTv9HfO74mhA3V3Fy3gcMBHv9ZLlx0DqNRCwHXGtw2eMllNywq8WrQ/VUVlWbjt
eeIoHqmqOQqLlm6N/isQ7IiNbK8INKLSPh5Neu1qv/oOYy5pHHyyT44qTX83Nc1+OD0N8Zfs9Trp
O1rEDbRC62jlZMOyuUwuKRoiBaQhExelOWv/pZxwpR8XWSIkucugF8iQsqT8W8a7Wt6172R4psib
bsZ1a9AnWDRcjFi+2yVyYRReR0yIW8/2D2t7bmRsSErMVIX3TmVqC+PKI35b1kqMunjre/2hNSrx
zhVVqwWZTYGkn377QMjmDOK0ySjangKykt1H4E2bn7Ju6ey5eLZr9B2cCzgTnt8s1Y6VTfOodZ7d
SY48a7VvMp+DcVH2l8vdU4LxssBGQnM7Z7cDDROiQ7o6g5SBj3zq52Pnc9njqq2wL5/YSFI9eF/+
9XJBhRtd6V41P342sqrnuDkJ/q1faQCyj0ClXvvlyVt0YU7P01+5+XmcsW+uwFQvxdXh8nHiQOS4
njHTU7x5AKJsUFoiLI03QjWgI3b7pz7ZMcqFK8Vvi52VWTpv4EKeskyL6sfSHXpRr9Qb5zDpxv7J
iyNRCfEHZqxD0gnnudG0mUOiSQqBbt5Q/yKVShoHSDTtsmhTIQkB0VJ7wxgrNYLISyjpWzb7/sEC
o0wK46ObBiKOE+0Q3C3lEVoQA0LVu3jXu6as7abYy1SU9w/DD6MIYWuEsfewnijjvz8LZ5e8w4Bu
C5HQlxgUcNZejBO+kwmCiJeOoI1HH1i9fr2S9fKTfpO7CMDK+FYAauFy2FsPdnhV0NaZgyV4GqYe
ZJn8MqACpfjRwFm85N9xru9oPvfL93zUhaLQyjQA/1nRmuGXmWcMf22mCFM/28S4H/kYa4QUlXML
yWpKx7P5uIEtQ1Ay5dA+QnVH4kHJFrUPv/WB+yc81VlN1nHRPBERl4J0D2u2vacYSlvR9IbPdOO+
EmznzWxKqp8LZ7wutSee6nGaRGgcZjH3M5eQB4agqrhKti6XmGyPUad/xdZk5ANXeqKWLhI+HQTv
BwNbLyHSssRHLN/Ege6vU+ba7IVGv3omFKevCew1Wo4+0ccuBTXQVOUFWO82vA4ufCsgTWPIBOMQ
HEwnpWmmMh0sva8pHdSxPEdhQePtuf3LOhots99gldxCe0gPF7Tg60BEsoMjXYe9OslCdxDceKsU
fRUHEXPAhTvYUfub1Em0tI+qZDfYrxYEZmO3nSvChuEXwB+YQs2ia8JxJAyt9eQj5bf/tJ9pX6RL
TNw/4V7YpFBYM/fbahXYlE9ASNmbaqghlNIEl9pfX2yKDfo4x9GCz36tl31EyirQAExg9Qx04Mk0
sTapwfZBhQdO2MNkbeiPEy8o9dS99lyOSfPXpo1SssZsjTTeH+W9MmLFoOywf/ENcOdM0+rrCWGS
3e1XcJE5zIhNf6jZw/JqdD54AB7v243uFAa7UKfVjKrpq+K2cWwsKypR8lUz6NHr8CjH2MB5LsGQ
DNSf/Kck/4kcmczvbTPX7g3NO6VEQDoW2ezztrrJ2sMxer+KFBh+MabPz3yeZPKRWjUEly/+iDUe
56wT4XpF1R4SHz0oluKvp1grlprMLYSrNgf2Dj7AaI21WSZvdjxJaSj1Myf5hCeHlvKmumE6M/OK
FAoL0P1UtBov3eLrZHKzr88p0WjFrA9irJlTvaqxZRd2DJylfI8GwP/f9tB7nQDhSQslT0OxqjHA
LWlzvc5x0UQbh9zveSthIlVbhx/NffEtxIgUrIXhL9uJ7yQEIV28LGIhJcKGKH9EosAa3B50IL4c
IcOrH9zi3TavXfoorzT6mHXWt8Roi0wsRhr5+jWDTY5HRnizYm6Ahj24Kz8OqJTCSuDU6GAI8Mv+
970Jd/CyCF/8v6xpamomKvhi807TYsNUqpJyjhBnU3kL1o2ozqsRvJ25VJPA3UD+VexfyDd1Jrsz
0gzD8HH6imTHMirBrzk73Vz645M8Z17f15UQjlRPMUeLWSN967Urwv0xXxzeF3GfSteO0yBGd8Hz
hbqc2ayXN8hMKLrcJKbjFEYQP0+uvCipvfzRJTu4CQzG07gv9XFLT89c+7OA4fgwPbj9dsxfyoj5
lT8NmnmnFjZD0jNmm0J/dV6OQQt3Z4m2u8aKdPtSkGtTinOGJK86zFwMUrcYi89lhJRCoE59tD2G
uHXJVkcDhFiEyemZxwqYxq2NuGykkhKiebu43QKiDkRQDTgzKRwcmg/Ua2dDew/HZ/BhKc4Re7Xl
I1UlOSJY3EYlv6c7R/xEFgZGCIwTWzjislVsA2ysfepFTrb68EL39f/RiaXbsOSe2r1K3bnek8/5
QYULCQUBe+uG7XhTeiMnY2qEZ/RPLvQYydtYL5ReawivdMQCveVGGWwJHiisRu3C1FpTS/6jVwyx
1CdlNWp90id/Hg5b7Hc7jFb8Xjvmo9sefTCAmr7VBAqqy1Bk7L+SxvyWktDKmc0PTA4mtnKsojNl
mvwo70fDDo9g+bOA01VvKrFQzisuUetUmqNMG50cNSqgH03H1/cigJ//bKDfeh/rmWQyOeOmyxoc
ZI3kA36NxnZUcKRBl8MLTx4ApNIwK1c8QnmePrM2K1cuBnNVJZCQwMzSWpdHqrBYd+LvBAOT3+jR
6L6zVuE/jjed2AqUkxCCsKedH6656ZwWfKu+igAw9TSX9IwEDaL6dY1p2Gzr48sWO6LdQJyjr2ej
5TgwxtVk2uKMBJ4jxFMv8DUe8KnWK1eikDnKBjftbm6ovuT8hZyfM7PHEOgXmW0wDWcQESLK1JW1
aGnRdZwASgiDfKMknCddIGjuhb0AgAwSZOo1Ro6xL5qP44ENNe4g3yIsWgCkVhcnk3tVw4hvMLTx
TeXJAHU8J4zFCn9kIPLXnJeZ45Tk+vJ6moSTbHoxEv4nK2yMUmZyHB6ikzekU04jQPCCRWvaKi7o
C9oOSnKUrJFuoA7jjtmLcDavFKVppqev8AM8zzo3vsBPOLD/OnGyuDI6go4mFoNu+KOsyYlYnFud
lEFDP4yQnSJSF4CSiKtJxJi6tIynTwzVlm7s+h2f+ZipCncaHtCZZAF0mt7YK01SM+zF34hsrjhI
TPEs+ho52XWTuNxBwiKs7MWJilePSTkQaF+uepTc/KHzOIEb8uAI5Ww2DHInQ6x6c5/hCRzF7SnR
5Mz7U1OYw/q52UALVexXA5Nqw0Qr5qDskXjor4jEXcrc7DZD2liy3aYQgTGhig6JIzniC0rG4Ndb
AwYTgjYdkNccrBCZbfuWNSCBuGootLqLPBAOgk1jCYTg6Uqss/0APu05NneuX3EV+20T9OLeTYEe
qlihegXqhbTaFfC2XV19FDkC2s5kD1xrdHRWvr2yOtVkiz4t3C+aAaW6yR5wf0kIaEGqAEzoDT79
VR9O46e7VwnTEkZvGnSKw85vBLMyhZIx0LwvRHDnhqznc6djq54XX7+BX3Gddxtq779gByqjzQ1x
PIr6rLa2G7mXxz9tYxq98KJilGDBujNM3cMtL6bMHDRkXILb/ghOUI695sIvMjVOJOCuzY8s+VDV
DOEWVATBUWohwBPo08FzoSyKihTzi29UvPSFnp9TAbpDJcAsqrvPA2dfpRo+i9KK/QY/l+czNPr2
fCx/shdfzCJPCJVbVhtVEL/1movEYVI7YpnMxCMM+UN4LZ35LVW4oWqH5Pv0ATfN6nGDiQG0hUNF
QNe0FLOxeufs58mdlUJti3CVt1z/mbPgGhLN38uuKFmgwRyrgSUKKpu8afaiURYMAKmONJ9YZn4F
IEIZwHqEBpokH8JFSVrFM9WeQilTiC1aQVs+mUOPnONJizu/bJhjKUQ8oEW/RiKkDgLjOCXfcjei
YALy6M3rIXQIgxbMO148kme74SoPgBBntKUlHoGKOx81XjWWJyTalLK6Eypyjp3tmIaDeFolxJOM
raNgiLm7FElFZOrt74lRsq+kbOGbVbYkV+RkJFGNRaPJFIxxv8Btupg7sOdisag2MZcQK9yNGe9q
snIi8wshdI/ZuBt5fqiACv5pzGHw5DBSkBArCjrj9VtFX68lrUOPcLXZl3YGb7kBZvmhHo6Q99f0
sbQDu+6kgc8raep7gG/GZnMXsbmL9lxTPc4bs27lG1YVihYfA3F6oZt2osD/lEH6Q4HU7QZcL6/j
eJQPIbks/WWvC+R+3zvnuIOXv0p9shj5atFnYRKDotO0e+3bQpFWx2rfcNuoSb1T1vqX9uiUEV9b
mA2wMV9GtOKH3fry1I4ehV8xVYmGhVbbke5bOSiYB3YGSELRjavhIbpys57wisF+KZ5QWFKT5oox
HsAAaw0mkbrISx2OrEgiouuckIEJh02PgcCb1Q9PowkLwe52+ikMT121w674QXnADiU7x1+L0W5/
Ut3T9i8CNIcpxi2kXlAUv9P4lJjLjzbr2pGcaX7kuUvo2QpQ2bRHHmCzxPbcDsgYZUQiVWLUS7eS
X4UWiBeLyxX+GgBQ5usrRvPA8ZdyoQzy7hgeaYCcI0//GJE37Tw6GZ3V/7bhniKNRSiBWl/gAV9O
8PSFfcJHONNdLGnRs27yQTZTzLzSIwKhYekF/h1oEFq35Js0GKqm4F1WDvgcyX/RJeUDOjpMlRTi
DTJ86YKYl6wqVA8bYsJwhvP38mPs6Pax6JqSBwlOd7jO/dksdXVp0a4SjtHiiy9MfEDjLoRQgx7x
4qlyGm5mS6smvlg3H/4y6wKF2JNJP7sL8Wpq+hwSs5UI48QpcKXxqU5Uu1v6h/lNepaP6S6nxbbb
9F0KTHCAvkY1ISKt72igUr2+0ZgRLeqKL6E3wZWZVQdsDm2WMXjIogtn00Hdbn5InU0zQxzZyAb1
4f1QOGsnPcFMrl2J9CKtVvc0e6Pl8hkwVKgq3XboB5yFv8us+lqI2Vn/U9T15zaHA4Lub2XzBJyE
2tyc1Q2kCN47Q9ouoh/s16vTabqgrpnLJGFlU06Humnbgs9HAtCEDwd1MsmznKx79dGZnRjEUvA+
Pd2InjTET1w0S62rn4Ly6bvDpugBfP44+10V4BsR9iY4E6txB6xxcPfanMLuY52pmIaoh0XGaEx1
1x7S64XeYwum0Q47npABHIFf1eDr/yvYUqvc5mUUetTyJdZwdNiaJodd6X+FHmclAyqprpGOsVt3
ZBctPFyYHNibgltPZbPN67TX8SilyJeicBHvxH8L46+OZrRF/vrJoFmxDVUXA33387hflpwaRxnl
4ybtOOoASqiSqA0RrEVnltGpYT3BdBweedKJRPqlNo2JsnpfX72Jc7RdO4qrBnGUqd5uJPs3JsOQ
qhpWZT/fptELkOmvUYzqIM0iJoY/UemNExQYCP2DJx+t3LIoxNFzZ7w1aWKQ7LbVViSfSNOPmUd8
2EBCswKNl3a2sH53BxTI8X6h9qfPwDjWLqohqSxPiaWBeJhlCmzU9xB4QAcXyE5rmt/C10qi6A2X
/Sh6xDPcbOpbA9h5yxOpWvmJT8mWzrEBwMJDYsgN5ERG3fd2SNj6vkR7EhTd1qi+hAPCYZ7duvPe
n1AjEFeNTkgzfnvmiudH7ADCXdQ2CIhd3oFvDi7QKce6Sog/vCqmqXgkjetZ79wYFzLlwDKm6lXO
r5m/ckmiicbhAIyYLFe07jUNNhz63n77MI139BFryJRBun60xDT2SqqbHpVBCup0JG9D8UyPFhlf
MrhDsWVkT1fuG6/l/kMRUbRQ6FR2n+DpN+qJ8xVdTB4ysm25ENrVJtbICjwZryCGrAUVHPmELZgC
9NPomPoSoqtt/4BuQnpYn3OhvaJy6PXP6dgjcQNLDzsG9MwXqY5jmaaHgpFg+M7QDkdjQaVdzKVL
FlYlpImJ8phYzj9JMWlhz6SMwICFxHmeJTjtyqzwnI3CoKzSLVH99WA59pDxYVaDtt52rKozQKZS
plVWfsHvvzowKUjkc7/JuIZVXePjh9qV9v0v/fKBbzdXb9mCO+EdzkhqqU90509DYIkJWjQ/W/6t
3wy3V0nCLzuslWsL/0b32Ak8fe9CeEQukLU06S8g2YOaYP+7JboD/LpmWMMalRsYk/Ajey7SQFu1
5MUplSgVniyfyRhunxDvMliGw93KE3Mhz9jah7XZFWoTwgjJjUgZFJb6PKhx+FdTaUD+NSP9XBZW
CAw+C9wOlGyu6w9QboELCk4VrJ8HBfYvav9HiH1qMUID4gVLbiAknNNlufKojOBSiX9hryg9MiBl
b5999U9sWR+OkOsHe0u/y//WjPtAcqMbf3N0zxLc0uwNBDOtze7iSG0xLZ+B8Z6ncU7/3fGZoGsE
6jadITmatOFXk8QAQS9I4fxVKXotApCOpzjpWHvXsKf0y0qIphHTGX6RGPzaQP83z7JyVTEv5ZXF
Myv3IyPBETCzv0yHhCHzypXsJxaCeQBMbkda/RrVGm+kjv5T5PMyexzjvZ3NmBdioQahQE+yXdyJ
XymWuWwZMKEh/gMbY2arbR6J8IwzjBHGCBv69zixgnWgKYAtChiG21ak7u8Xn2Jk04hdAK2H2GJD
lNgvSqodQBApkJEQc0RQV02nG1zIRMe06EhbPdFhKdU6tRfR24gECtX90aHRfpXE7E1qXY1Iu0u2
K34xekY6/sch7+7fyXYslXvWTTyjPGhJjbjhAcfBn7mVVESQIByYMAJ1TIvl7Zdr4BMjKRND/eGK
7X5U7tq7+11+WujmcUODAPW9Rj8YdrE1K1vOo/KDotF7oQv931ZELFH3lqcCFGOCZNSZeRmEG6he
jVnvFpwbLJux/vhAB4mnO38AWghBeWOgNHrDrYrU609MO8/mGIOGCP7sswbQrN+iNBETRsflHie2
gmoGpHzjGCSoyE30M88ZibSQ1rgck9daxZ6zUOzPsYXlOnqXpgFFBzS/eWxADp12dCK+03poGbNO
BbZMK7HBTK9OQd26UVG2Gi5OtLxIXuyJhBlIzSWxYUVbx3FC6MYNhcR3ZnN6H+ZccNZChmjM7Sdn
uv+c5sY2k1ATJs61NB6Cj4ByqqVxBDNGX+P+0DiBvd8aX7vpdfbYuLLkFymr7tVbeVS6pNME2fEh
H+CpDmKXKZ0OqvJ1vLa6gXbmIMqctV2ROm3v3R8E4fmOwpqMRMRBc8YsaFABd1twgtHODcLpa4Me
uaLdQPXl08tUhx7dmdHIuIMu0V7E6dHWrG15MbaO5y3rcSlJBz/FV6yogkYf3WtQFBInrhpyLF1S
pURmpKTpXrNukq77LaLclP3n8+K5i30eneEMAJRY+ZD0mBq2b1qEVVbMSDNiIhYAFU7YQescWkIJ
joNoJaIE7CRhIyIVv5KWUwxenanvqa1WVs3K1QX4iu7mMEQckm3YaiZ+Ri9IQ2HPcSUO/nCAKZfe
prdzAfNyCxQ6osha+iflrf4xch7wL3qAoo2zqZTuwT+DISprdMMBOcfLeRT12r0TcVjRN43UpSi6
zuc9aWEmIInC9W7QcymWsh0eTTpq7boK4/dUjPg1rVs+FUTX7nMCMk1TKS8J2xwoQzweKlva8ywB
O/TqEAkEVgfzvh96qBC3zm4nft9Brw5Qefxmp4ieV3VZpgp9GfFdSNizPh3XQFJEzuhXKC1ZN+Fq
pV+RoS1HlBJgGvcwc9BybcTzPiVDHOTwexi7Wga66AsUvrUhH8vwawcihQBdjKbrBulyO0O5VLci
DmCDxmAn+pHl46IIU3UvJ+v3ZiPoW3owAKNEKa4RZldQNt0LYS07pHsPSYmYs2ELdoglQSCBvtZT
5ULHgXOOpvYtDmh+VJqbs4ZPSk0QJREG3g6wccaWLFqEFGoOjo49aSFMFtHkFEnFbTN+Dc8kYBis
uif7rCK93l/V34sZuDKDElp9N/k6NBzjR2QXe+CHivovYdFZrm2l39vL2lztQdMG8rV+i+47nTq/
6TJsVBF5ZXQ91cckPG/xcAcgqG391NlP67xR2cxTUjRpYuzz4UhYDrILPR1Ry7ToApeW2TqY8kiH
epRXj5gDmm+Yes6a2GHuJXGchiWCzN0pfBQyxxXQ8hSGJM4ZjnZbDfZ/+N1U3BqDcaGEhmSFLrFE
uMTIDe7cyNAnG37VA1eRD1rXV55h1raya5eUYPWfC1o7Mnl5x1chbYlMI3Af5uxHSVD+ErnrHwPK
c2oiKjFpTKHXz0RqlVMhDdcfWPxyZtf7AStA3J0gxBU3sqXsnzXfPC7T+bdTbY6GHFhEjoYaChsZ
vBNNcRrZ6IKSmvGQ+pELS7yzJHtM/ZLJkJRCqRXMKMSkNHDxa5i97f2/qF0YmLVq1gYtaFaAfgUf
GAeohY55a3jXnW3s/0+qyFknr2ofnxAE3uH07XISWirCXl1liz6HFbnouLBfrJXpD1uUJMrisL7R
jTB0R1DDvoSqJxIf+4eGJooprb3je6lQtBAI4QGc+Hovg2PxQ4dZ3pfTRV8A+Q70nedlpgXsZS5M
6U1tXZjIxg9bv+kZ0q6AdBLh5A8xRWH3Ily8mrDSOoHicrjl5m9ESbum4XhvPQ1DNn1Q2ZUJtoCB
QzFYDVkpGRDH3Tlq80zkKre7QhX8oGNo/23K+YSd8bu7fECYQy9mPL/5lBBNEDVN4ggUQnNsngaC
zrT9634RE32ms+wd9wUXRIaqitZhZMXY6y2pIxknHh5CgjnLldG0e44SV+P5mqU+VtftNKodegQu
Ho+ks4MUBdSkA1/nM1iwofoDzWXIOebH1qXPtVnA01UqUjCkpA+P6ee3Uzu68fXoSV4QVuJZBGpp
CKNMv2VOy7gcMFqCMRAy1LForvInp4DHy/HVX2NSKKtktUVHjs7JSfACFBxkm/54qlE4dfd6LKhT
pNSY3vQnXAy3795DoOxALFS0EqcmmyHGgfMfglTVvkolUBRHSMK21CtBJPq3ptM9Vnk+SXGZuWR9
bGjaWxk816DKsjMeBFj0jhWKuVabTrpql5tgmYoHdBdSzct2/c2e5nCLlFSFiLtSa2P1PWWnyOHI
t6yRVpR56E5ZdXtu4Hc+B3HVxbdWskmOqCzmTjk8iDdWfSLq+MHG2qftQhR7a32xsM2kX46pv/+9
EJd4aye2SB8QeHqSpBUg9Ximy3hoxXTSl2WFEUiGgyk0fKiPtVEbBgl832kNEly/4UX7Mh6Vs1OV
TtgnuN1Z9EXLE+N7uRxjYhmqBsleMDD0+nH3QeI5uPrtzTOwZUg/DTNSm+VWfvSjlsccqjz4Bght
ANYC8OQU+WXBe9hbzG1w5z6nztC6r0rw6yUbwt+gXRTSlOhLnFdU03/Qf3Up4Rww8XCakGAEqeHF
iPRKq1At8TueW8/oVLnit+KW/bVOxPSKmyQY1UWUAAKsbwNxvyOfi4bB27k3nBY8Nwpk1KlgDAU2
Cb0A0rHDYsKm74auY4wcw9rm0Qcwnig6Jl8sGL0XgaRAzj1k6CiYtEyJIJo3dUn9Tdox7SACI/Gw
syppXJTpWQJHYnYxB+aNu/aTrxK7EdbJqeR9ADpsr3iW/bLJPMvBJBOGp64+MoxXSs0xQd7OvGVV
SeumBxJRHHgvTSIyH2+woh1t1WqsLBASPfl1xfWQSdQ8tXK8HCAdRnyaT7CJ1jwC9/n0FDoujvYL
GOFiREy35RRZ+YL7h6I1XbmZYYaD7CuY156+ksPynq4SL+zJjdckD6BahZrRCE8REpHsdvE3rHmv
dhyPx2oQc72mB6yHYWhn8jWX8VA6GaKpchQ7XgY82LCLsrwJF7YiSG/4kfbRkJSr+F2fnNIQQ9pt
9dFZmHoQYoC/I4A90G6T2CIpQPntx+OTc2PBBbOtB5sPuubEziOoj2XZTSYRRq0VntP5TyMLcBlH
IoUjCSCn2hOipT24mbAedJr6WD9fTu8novhChBedG8e1X3pyu9ML6cSBBv8esiWA2h8GWw69CkES
E+KqJ5o8APjLyY9SiFD6xg5gjoTiCxyU1HWIUvEmxTHjiffP0qSWv6YC37v4Rf3nhUYkLpA2ntXN
Kwm4/Efx1RVfR312bOBpiMTHc0zFhMVEZHMjRVJ0R3pu56WA9IxT/U/Ou/t6P2L4NyC4mhRCOmUP
NUybQPTWtQmIRaraxOUkLzCOywCJyg2/cZBf95QxC031iIncauCtOtRIyu1km1hCCWnUQT90kVO0
rB1Ks4D22EV0wlaXVKcSS3i6VUwuOGkTeggDWcwBHRIGMTytmQutpTKcg+cnNWygfSGZhyiCMV5T
26f75RjcVygrr3A3Cub/JtM49qMg27LpjdAobhrzzH6MGGWBsi3VPri1CZFP22VobCxpYT4eTNH8
OZR12QofdBjU/8ypyGQuJl3dZVB2I0mClKj7oyUc5TcZUoNhidfJUmi+Io850//gy8hNu9KlNwgE
3bZBjtfONT3oU1QWSp/bwwW9lR5usBj9DErNo/AojizZYEE7HoQqPpMz9xIUE1x8XszHVdUdJ1ci
fVK3S4Fnb+2JAZc4/WelLIVtkZcufL4YnlZv4Spw1vqCCj2HjMR5rhib9fh++enLLpylddhknjWk
p/eh//DSYZHpyYSiB+G9XEP8iSiv9kquaCXnD/2fx2sIv6j3rgEUh2zxO59SLdAVhf5lpzug0LZp
8cuQKGgfnDqlLtIkKaupRQ1pswro7+L+h3oy60ZpmO435mYvMALFEFSBGnRzGoRvrOaKUvVtWz3q
WP5m/rOQbJyMg0Q4cLtWriKOryDF+KcNKWQO31Fb8f4TkAT0qzFGsJHc7sW1OYXQK8P4cJdXVKs6
kzrWvGxOd0ZDWcbkT2/mG15GAMo/mDlLvxDydsC4tuaCyRPrTziCiZMfZJFArilzGqAPlLbOPhLN
DXDzgpoKJyHQFXigaW10c9Fjx+/cXL8Dj5xj/vlhlM8YixUCAeDGaO8RHW0CnulNtgre3MwjcwrP
SAq0FDdI1kxmW6EaZcGaXxHRqN0t/+0aAQZmrM+ldshE5DounvkL7QGkc4qJ77pZ/72en5Bg95xJ
+N1zWRHdSZX5IgEkdWEs8Owm16pzLts55aPeIxZ+kfNRlqnQvWTIdPo7DS9MSsmf4vFw90dXCNG9
WPPNXYr7xGkI8Z25lNbZ3SVKm0VN/YHQRAUCzso10KmYGxkvveBfJ8W73tbbbnT7YvO02TLQZ7Po
11oJRXToYCG4Bzs4LvWfoskDQ4rYETOCXNVo3S4zBTqtfaZ941Xx7Ie5WCjOHs1Yb9QPPIAGvoqd
4voUbKoZ3XVzm93GggNbKRHbev52QrJBKvGNsvjD7MrlpCbj2I4A8kG/CblXpgMzodgcXoK2tYRa
1aNi+aw2vYPYXL1BXWgn70k7NTjxRyTZaV9EjhYNFAzrp5POpaLKsnC7tza54/ErebLzbGWm2a4W
k/CixOfsGKxZ2OrTtG3zks2pXC6/GxgcntR0JHdMECzkgdCNu+zWVHTKBfKks9x5qUZRi3MCo8aw
A0fcI9XwvMQ59bC0NmFzXnxYom79wtilTZuy/wfvY66Z7gPQXTpO/6Mpo3cYCqXYFaqDTdKKOVQT
bFdOQsY1kmu6J7eCvo8MESc1JSDTFwhW81aB+cdsPZ1C+wqD/FMufJ18Tnkl91xbX/R5Jriew0s+
8u7GRFlogS7wJT994g+yFyRE3DD5lEsYr7arYn+epa3sYQWvuMyLcJSk+AZ/ipqc0sKADAtkPTsd
J4JSwalZn+IQzykmqm2WCtBPu41RbHlGjh1p/92O6Hk4fxiiapZalKcOm3CY/GecnK1EYJ6PTcEG
tCb7aagVK8s8ZLpuB4x1kz9m/rYwYil/9Lut0/2K3rZXvolvC0c4NkYH/GoyFU/U4Rg6ZQQ5C4IB
9KGeogywPVZWqgs+6QvGpBrThLUishiNEL2DSiwnRN/fZUpUGdvi8XyYDTAz//cqseB1Wu8B2/5p
HG20FJKoG5x6VQRRvBVQAN6L2bh9lZ7EVuSEtB9d0hIhaFdqczssMrQFkHPMaIPjVlCh7UA48jTw
pr7YT9Ye77v1WijKafa/EZ2IjNmjDgq1B0XNOIs0qFvuIvmHncXdZa9E0kSrZJSbb3m3L45B3/u1
MCNobX3QeIwfhsmVEMYub+BEYBIX0bUWNezb9LE/qkSb0UjY4oNOGNNDaAtfCnZt5mEE1qfKUgNS
4Zj5G8/rS4lXrw6wFi+42l4Ti+hkI08vK3Wm3GPo3pyRAUYWJp0ssBjFsx0CIuWATgzzHWvYv318
aGQnk1WreM7tYI+0zG1pyLHwNUTEN88t3NN3L4Nmhmabh4VleuCw+0gJtJju7CUdgVw3XDDwVzGz
MM/FbLYNq3pWG3QNmM5mznqyZw7QjUYlJ7PoZvfY3udrUokfb565iDBMI/xsjKT8/EV8R1VFxPnZ
B20pUS4BdeoSdCrxRRVaQyifvgaboYG6KmGmeOko4APg5aWYO/ZReNawW6xYuNh+PJzOeRJ0Dqp4
6aFECI1oYbNOzGpC7N6XfEHW+a6PvXT4CgjoYqpylY1d6OzGylIb+DQ5yOuICMYzM3rsca9Gsn23
183TowzNg8EjHpKZMUOMUbfBiz/yY076gMnFpdxdcqJ3mZD0/lcCDItMUfAHTLJWULgkO8nBJJIT
z7YVKQBojLpX3k7BNDWI80VLALGRzYTsKGgtFhO3eaXHWcU9Mb+p7uGsM6UnENPjjehe9XTSDGC1
DfRhV8mSV5UaGkbxagN9tTgj86pOgR8EUCXdsdOUAfjS7yB6z/ajZ7jQIkA4queb0y5f8ujPmcTn
cr8zK8/RKj4d9MKU6Z2N5smu+YERZRHzQ9NeamWQUO6uQoXgXaJ+J5rUvUzY38kkworPHjSc23lN
kTt8/w08OmxG1sIOHTd4OWX3cAYh/zN9gf8pGuGY4Tir2NikrfmxQFmAx+QirhApHJTO5VjSbb+2
5KeqSaSWJzFT9znsriFnOjL1eZ4DTnEQQCTQSAzMjBgvi4xwwrpaFrC52gB+qB6Ue1anLn1t+Dd8
30wkRj3I9GHCEMWXsYR4FLc90xxX5mmT8jwfYM5en7pm4HqNsHAM0gghFUB9zWWmo2k2i0OTwUbW
ZYgc2eYQTexki0Hi7xW0HI/mPmxBsJOdH8QHW8zZcpE9kCoL8RSEyY2y1tsQjnXgK380MYgAaM9B
7TNYyLC5rhAIFz/t1XG7q1FpAh10F5HaSV0h7xgCJvp7fTuFMSbLH+OmcumzHLgrvrB40OAAUImo
eBV4nqfnCmOht4pKe1rTTVBg2lO0dY3BiURwR4Pw0pyP8DVDcZV7IG3oC3GFtDcwpzcmqvxR4jO2
vdeLfA3EaVCM0q8Bhlcv69ij7GNdme0xnXZoJjQ1T2D4g7WfdaxV27zDEw4ZMzVogeWsMmDkmOas
WOis3rxRpX0d5d8dDhY3+BauOecWz9+LfMtzr4mBta/g8kyaqxePMnrEtwGPRrfKjUEpToayjKt6
Jyh7eXDAkD5ecZsCvyvAxEqCFy2R+5FZ2A/0fnUonW7s1gWzT6BODF4vJBe1H22A7PicBeW5TnpD
xwoflmajsRft/cctCpP/rL5YhHM7BmVPFwH2LHQCHn9BG3LLpjiq4QkA2lSytlX4o/A5WDrDYceh
uJdHgALTu8GLdDR6uJc7fwlTKDLAqD5kPFtj2KvUrbyE5kLxfdJBEYGOMLEOPZu+9LBDrZ36H3BS
4pm63h1HLL2JXJWWVXU0bKmBLYJz8pztHY96IqCfCesItgWAtsrq/MF2rn+4bRpBbRZhUb4hP+0E
EeCS/QqraAp2Vfokmq9QE2XRAefjGLW+t1GVmmWXa/SYe00yYSndgzIfHKh9ql0VDvtxYFvotB7v
s2IG8dCizZUSzeJte1wkqHXCBOcQGFdims21vILZWoePsx7cMdPLHi/vj0bMeo4JmzP+sR54TSjG
ZkWsB+1HWAukrwcxPRYaIyETEUKs/hMZglvOCaoBWdfV+VQnJ03W3/gExc5Wpbnb+4gr3to4Je+I
3VEduvVa2UCa7hw8nGa6RQVq7gdhr/1N4sKYRe8JCGO1Y22yhcV1/RS8cQ8I8zVzngoOvwoSyUwf
6BF4wl48+RhE5bx/kkejoDzwhKNfsDX3GjZYesxfO015+EGGJaKPznuiD25SzF0nqgbH7yIjrrbB
qP7jCHwuq42ECeCHqIfHirLPvgL3LnS1ozzdpeEpupcvHQWSN4R8dpKC8J/kmQ2RZ7J59qrddjWu
B+uJFtaik/vYp+ABWHEdpumKpfxbTaxHL393FPwdB6WgDnwj9X6b7UzrwFtbXM4JTo9D+jobYIhc
hzEiCj10japBYs1aMMJkCO4tkRG2zjrvdh1eiJab4+kUnYii1BqPYuHu49JrcqgYM0YvMplqciuq
24RRJtkO0K5yEzd3i5zZcNbFBb9623+V4vzeo29AHlBwbadT7ffXqp7bvrImNz62yCw44Y108juS
DUs0G2CA/fOEs39EfVTtTakmx1MFhGcNHJzPlstiikyvad8Htelr9wrY5iRVHXgeHomvdzbQpm6h
NwsWJ9Kg7/O3TpQdRCd6ib1Ylxmy486MkAOiya1CpUjhRsaV0QVKy7WkF36OKPVvHfbO9lrwENdy
jZwVjYdh8c6+6vTAiyZJwfxWQ75/Y3ANEkl9mAt7wOAXqQrrNZIQWxEtyMopgUQLQpGFtR+gniVI
e7NDZ9hduHcH0xArjtBLIM08Y8gOfIs1QIsQ+VnBWFNDC86G6syIOF4uZbCtOQxg5gr6gEWPwwjd
uM+Vljm7cocwGXQXVCV0EuZ7GA947/V+nvXKzNozzfHsg0Li2YM6yGveGUUEAUprsaOkyZxyYNUx
q6zKbi2NmtEtQw6fy7C+MtYc+NaAJqL5uhYQ/3Tb/Jj7Xu3m2QFHBZijhOas1e9buWYeAMd9Kemc
7in8JKQ1fxBpFGU0S3Oj4LgbTzTpydmdfO5WpGz3Nxc9d5whb/SXTqYLQTqVbPqHmsTgzPcr2QVz
rXJUpc2z9WWdYEpXASePkxRWSvJ1u/Fdvk/qCFk13rKQqGXSeVRPAV3b95ur/7FGdF7aX+/wCntd
eC6eGKpDLWVZQaY4iN12w/GJsZq3uT2jFC9m40NIOe6FjghYlhtAKjV6Ief5woaNXlznNhFWVvyx
GiBl4+/CRy0ICGU/oO/v8aIMctoZekDZGymn/s/K4uRDiZYivsp5IrlPhQnlUeUeNfgci+gODpHM
400UVuNDukj/qioH5Grw5o/rDMssAJ5HEi2Kp/xxmob0O4GMu2TFYrI3eANSmmk7MLcPvwilUUkJ
rR2nJ79g7nrAcL7oADumz4eLy279rGxfn5hxi/6pamGv/OkuCfz6tC8sCwJCo1+huUGJ7+cBf/jn
SCiB4P0jqhK+wTyR5McLj1/53pYSqQD3MxQp5UdgmjiOVPglanr+2UQN3C9vYPBw6sVc4UZZYIG/
yl7z/aX252YRiASnaLbeOjkHcCkoDAfkRUMLGBiF/p0KhwJfPVpVryte7Z2TnLeZLRfUTvMsFdaG
yZmq1yQCI9B6G0tRSbu1JEMQbD6Krntq2V1gWA8DXvGkZR4HGwmfyK70FugSSqnGzP9nmwHuXUvo
pq8cRmQDiy5sxWxK2U8g8igXAEsY71PYz+BjiU9I7YIJL3WURLgSOvQlhbPP4xmiOQ8fIpDqMvEl
saLT9X6332yNWH2Qgphf8INKzrvUcuFb2Xh2EFeKYKngMGwht9P3RleVgqVoex4LwUZrEOhRPglU
SP5CbQ9nXpf3zZ4Ofr1OCdFCwPy2Pc7R1TlrZIRr2LUAQDP3HFZbziw1PADIKkE6UcXrAyx/jyJr
DfdzKf6hT3IkNRylLk5jjmiQH7dXMVROIX8cH9NQwl9CxLCiyUnNZNb0c6lASV4S7HbYcC+Gh6cl
YspGSBQAHTqKmUuZeU/bU9Mzqc+bkUtTWUErTAAc8oZn2HISZ20NpxaGYFwEAWQfFj94heMkoSYL
6kGIsrq3ApJGjRIMgfo4yG3PaPMwEIFI9ukvvEngehfrkTj0UPSo33GS1UaHHbDetXIJiRSQzxOi
KdG2AVi0WP77WPVqj4jtfvdYQguM8YtL/dglkjXtdbGTek9RUOVw7MuV9zIh/s7h9bSvbmQY+K8q
ruf+ygeT0Boxk8R1Jgab6aaxIf2L9uZtNGfRf8rNlBJH4oeiL0I7I0cyyTnF6T3wDG6ZWAPa+4DW
+2jRebK/hvlQ8f0+8ziRt+90E0Ae297vIHv3b1mFawkuX1kb5S1Zrck4s4hHizG5sfjf6Nhvr6YG
EWZS9Et8EK3XveVw0qrXnfLvN9l+nthnWsZkjmrVOWxg1NScfOlFfAitxQO3kUaink0rttQ005fu
WII8qSj8ysiUntcMMsG4q0+9N5N+nyzzueDgTJIBd+XxJXalYkcs+SiglrlL+wRsNL7TZc/82gQx
auW3FRI/eRwV4HYYxhte0MCB8LO4/sqNs5JMl0OerD/m2Ow2qyzybxWjwA67G0kqiKsUc0YUNogm
8vXX+vhQwvD3ri2q970uoINLr2JG3HwMWuVkT1XlmTAS8YK/BV9VC4WVG70tg6sQfeG3BX+lTZLx
qfLrKOVRsdOPi6obhLDqH8TPzTfr6clZOED8PhZDS+TLRhjoKAJokX0Tg42Eyxa3AuxRWLoAZhiZ
odv+HdNF7ixZkemzfC2bPxyechwmxz3cPjgyjeFhmOcBYRAEntLdBOkeerUz0v6CBDbKbmsELec1
BBxZU0lF4jf/BbET4Z7V6TqqPUYS3wWfrGCNopLx1sfgfotdXZQqHFuHN1EKI6LgACRrVHzKsml0
Jo3cT+m7Vd3BJNvYEpUXI0u0e2TDoFzeVLPjkqiQiISP2Yfhdpa5Mz4ph5pvpO0o3wZxGlMKChtq
E1rzWVhKGLBcPbwQvOqQjg2Xo4TlNQEBKK+9diDjfbzHW4zyldkWAhHUo8DJnNcOq4Ym/s3nwZ6T
EixjZx50BaTAzr2QuFvWhOei0wccSblPDj8KLGqaHOoEmRlhJfkUwu+owx5o0feAdwD8EZcN6oxJ
/1VbcKaGla3JC+ZK9pD9mRcTNB1/vdiSr0DhMjxG8bQRlIMtrVyoULckRYIp62y68X7m5j+BxgsS
4+lpCUJ67Fc671X6/qmYLG/9Dg/+W0imQ8yp6xjVc7LHGEvI5Nv8GwXxpJ2tiqOU/HhKFsmMenWR
5E82f3seeV6Z9awz05E4dpXogTUTgf6ELnLPMRMGXSlq7ydZQzHgCqdp1f45DhCLO4bEMLASOM+8
IVIM9C+IQHV7HAMya5U5Jz8uuMbQj+t+lBqDJfSdMpo9rNm9cJhJcpS7Uc94FmPs7pZ254Ho/rT6
kSJ9MuUsMLGQtZEM1VP8kqyCub/Gr78VC/BYGlS0VeKBha3P6soSPDYBIZJIGS0S1jCM7ph8nBiG
Gcuj+oihGGopYfM6hD3uPvopCi5Aep7VwJxc5Z67irfHdzAS6n6vz5OExUlZ09iEa3Sln2S6NGIg
bzmawsQR+9dNm8O0gCOpOP44eqkW2/B/q48BC+wYQ/7DMemaxJbPbGYhUzu5A8GMOuU+wLDq383C
e8MMgXwaf/MzSoaGHdQ9YoazGPfOyqGwuxEA2lsiOHuOA/On6ZPb+3vl/XbHaEhIZstZN9qEIvad
L7yYC2gY0KXBLvKoJEXxCRaqqajBq7rBvxXufZDtWv3U9PdHZGR71vcZPcL8xrn2qsbfPtBpvq/B
aMmDIBcHGmCzhhCOd1Y6h/vAOEg2f5PAwlQX3wadg0eMipWS/stmCmnBH+DdcrnDEsgqcQV2OQej
FchAHHqRy1prRQLSGMrc6Wu+XdcBM0Bco3D32nd5fvK2lPk+/OnXJ+4DJOssg+RXy7gMsMjzqzmT
xIyvILLxhAsVaLp2gGLu8Pc/7EHT2tWncU7ouUGhhEWyoUon/hXbikwMMEQXR1akq7v8mBDVszre
ZXWpaxtyErBxW4aHlgl+Zs0moUP/1Oc8xMdVnDlocQL30d507q/2YRxujBEP29JgtXKzzb7I1udM
lOMBBthO59wEzwAh5+ZkbD1AwkjOabvG17AAxlcXc21w8Ca65/7ksMOM4ZR40psoQ6nV+W9REdiV
+w0UDqkIt3aPLBZ6dFpXGBbspKNYWYMngka6o79YYHZWq+nA5FJn9dwDDIBUisv2biAx03VFA2CL
Gj0h3ifIsSQjJXQBvYxkqzAsyUDlJTRBzlomXej9cEona2AC78zs+ZdjkWfgVo4C8oVoL7IQsCd0
auEMwapNbFQLPL+o/mzHYiOZhA826/BETfLy2ELcf1mZOfMoZUJxriUWzXYhnv5Bjg6Xccn1YNoF
2RE4JyrT+GSrMPOCiTXzFNqxUEb9PehMPUWBM6db5vI6Fx3ZXYm5nPai7mxY4ETI2GefaZOWNIa5
jDoeRVAxbai18vt8/oaMuceLPQoTEM7OyJsfJPt6BijYQSYvLOXjPoSTAIinGg4siftPpWmNvaHv
zniVvH6heyPnEpQ1zEP/aycM4oGQ4s4slKlxeDTq2E3vFROr/0GylC2SLQ2m04CCUFaq35ZXFk0Q
f1Ai2gAMnnngTdBPg8PS0sR3eDZbRq6syLd7O3cXlvYj+DhTF8mGLyU2/DFto0pNSEkWOvarkyEP
uwifWf65kdQc5opE69GKkb81l5vD+fGncKnkdCUYsdx9dk12Vhs4v9rajRMAY5Y6FnMnY+KaRZwg
nYPwf71yPFm7UDbR1/kQNTcwjZJZNqoCJWUjcbExzGM02upCODNgSflxOKANR83iI9rr/pIdmryr
mTZGMtmtlz7wHs9AAWi7RodfBn4tcZXH5xuMHevhEpa0/hwfFpkU6Mko2H3xNzO64iHHr4dL06rJ
HwIaCRNrEACu/BsBMW05j2hVPepsP8FSTbEqHoOYS9moQoXJOIAGGxJnGWYgxc/O5fPLs/5I04/z
qdnhMTRi2BqVaOZSelj9/cV4BafFVC9KVWU7vzfrok41tZJLGwaR5mZDVSozy/XWYo4cgZZR4dcK
++axlg7qZjtvJID3nccFQHUMXUvL+VssqN0asONG9JFx1nxUxvWUUeS3waTBs2iGCx/kaYYgJ2Fv
IVrlp5neWN0OLmdEimMz5BbreavSykSXBdakba3ZtJD3CQM1FyAhotTWJQpY8O64MFAvyWCABBBt
FdgG5lG02BR9kaprDPEZgLER03HnY2kVDTdS6Kz42whdoHr8yle3NsZiXxTnom4NKZGzizjrzGoL
8sqvdJozKWvqJsCvY4Ysgp0gLNagwC82pN2gcH/kJkAJIT7wRdc4bG46V4svbAC/afhyKX1mJHkg
JjhCzhVS2fweSEvxC9Vtg0150N4laJBDU5CqvgQNIaCwSrnOS0AUH3HrE5bCzKOSMSLDeB7Sp6vW
5flBk3m4WiPfI+jM7Gucz3Ex1EsLKNW46OBXvTU7R7e5TT32x7/qLmQp7+XIeiSMH8byApINMKTC
MAO8o8to/bEFIlFzIVlahxQ2jKsH9Whpf+PVCkZ+GUUCFcvwoRYI4RlAoy1pWcgDXyJw+Qq08kBg
2GITy5IzE4zhLBNmrNQzJybfewbuL6lPblmC70oAEkq2IrSVfKWRTCK6CFTALuxvaa/KJoMAGcq3
kcswXFz0Tt0XjVkxL1gbEznMyPa+xUBr6Op6hT8GxdPgxmc15U8uhiwD/tsI4pYiw+Pj7+uzK/z3
8Qo6fhd/zvx3LJ1QmhjfQR8dfiMmy7XPh34oN4mbIjCvAN/jpbmIV/JVIkZkjd0R0XXjriwQiBvI
oEdu8ZatDsyPXV3aV5jsPF9a5D6L6oz6PHzBBm5lRTtPv/l94ikJc6PvHfY/rqA/E0x1F3aGEYDI
ikmH/pxlQelouFbukh5I8FiDlCKo2Nz2giD7bf+X7TGwAOp3Q0+JS6RCACtuaT9pQGozgS+S0Dmd
K+e4SiYDBlV/T6xZauuMrTiN6ReukbU0adi+Xvu4Oo8aH1E5bgJmWbIIYFzA2UjTpNiwaz7PjSFN
Qo40yic8yA0jTIerq8lakqBScZKzeM/2djuNh7cvyQxcbSKLjdwTavvlmOFiS6/t/M9i188ihCKH
4g0OPHf3zv+H1dH/7J87q96B/McbLYvt1aopoE8JW8ALz0mRekLTpOvKhO/Ax0v6d5eQ+GebxvHE
sdoHY7+dV1+eEGQN107BnrjfP4j6jcAdUn82XLrTSxupOwe+tOYVNIo9V5vJe3Rs5T16UDUZ4ANW
Ig2xPx9yTk/r46PLs9euICAklWH9YeLiyJ6QC5t0XPdh/mwbTWVD6oRFuLQX7wb+fx/mmzLy1NXY
EqCvIh2QH4DBiwYHc6mq7EkoJmfNnMk+Lv//m8fRHO3ZMPejrYKmEthyO+67oc7d/VQZS7rl+zQr
EEdZ+bxerHg47v2JIH66FM6RuQFAGVg8bwm7+PFBjEvkG1S9U7cvVbfLOeZIKE3TrRjAyyUXvPzv
HIwoY9vZMDzu8zGBadAE8nMLpUOfzd8gNVBSmg88UnwnYG8RHAEL9+nvK9xDxbo1KaR02ohUhg8s
gad5wsFm7HlNJ0AsFXVbEu8HgXG1ZjvlSnXujvmQVEvPtRPl6g2N+GIVSiz2W7JwACu1ano2audt
o8ZPwjKlTxmYwuB+3bGPUb94cuU8JhLrVj8No7gYm5rCyNAY892luymGiQRrtB+Zy0widoX5N0XK
onrGUQSRyuSdjwLKzcvmKBatqk7SN7JizpgMivs9iZ8EKz06/mCRAgey9ifSNd1jJwvS0MPH4uxy
FgX2Y7w1FKIDZLUHM6gK2Ffe3TBMSpCz3jrIyr82fnKhBAfwJRytQyh3QkISYRyoBWHmJ+9Nlyeo
LoyOurv9+dDGULB3HFiboyiqZcZo/foYD3OQOHY/rJtcHfJhykP6bPrmGL/LTfy2SxzxQkjKcaSi
IKLDu9YWR9CMBfpdEQw6/aiD1p7pnUZm1LXEJX30/tOm26hTROAtPigSrE2bH3FrwteqCRySYees
SbuKa+APW8mOz5gcQYAlF6jwt2L67rqDTgtQdzZxMOsHGj2juvGpv0582PPvOMyh6MJxvJFUsuNF
p+4Isria3XI6i7qstkqbc212VTwHGFPXSMyUf5QwMSR92fglAP4KLcDbyjB0V0PeaQKrPwzilg4F
mwvTC5xCmJm9zi5s2Pf7gaB2H6rV4ytRKn8p5E5lbRDSyeXLTMXOHvkGwFCouF1vzxbhsRSTY9oo
oLyTuvrpBnvoYQCk2BqknJMEmcFWcm3TEzuqeOnH5BWoGJhC3X4cJYBXsPpec9ZZZiML8UAPeUnc
wQ1LWv42idSnc8tozxEwDvf8lw271ECOWqj+topNbE33zgln+ig7sIsfg+12crBTtxk3I7TAGk9B
HQGPchSc9n5Bj1sSfb0vqwZ2tvWUYJU745FIvucgdgyMhuWO/JyZACvoYvv+qbQRxTlF9Z9dN0ek
pZuig8V8cqgsR/qppgKCf4M/gwfMnV8MwssMeVAxTtPzt/RhGgUJiRzLw/d2GSshcUA1jlZLHbAM
4h1UVsrxqew+seVDPp6CrMQ+9Z8RlG4jRuBzXnTQySQhi7GUgPUPLMmwP3btlJg9+xxvdLBs7ZLr
kuDdCaEO2p42XhIYoMWS1y0PJu7C3J1UYVw4e5XLu+36XlsLQfF+13uHYux1L0vd+NsHRkOvCzWX
dSenhS8rNdBTwn4Gk8BUepfyIolt+YRhW+Y9Hw1y5DGS0wthZDntiYp1dcqxHubIdiOWFo8Ecayo
RvYGs77/s6Y0IADILRHJkXzWaNbMHzua1vfHYrICZtzWJwbNPm9VCYnBV/dhtGNYcdLzweLAgFLx
aQ15fe71Q8RcbjHIBzCi47Umf+d7IGhxHq3ia9bNyqv9idiKSK26bpR/YwnsV/W4L+dYfzqIJwxa
6VAK7lJL6yiWAZAX8O/7iAH+VGMY1EMKDC3KeDgfNzIEFG0q5VbQ1FojthiHv4PIB1vN174olNOz
sA4qaMabBIrVltaEgqvx0mniILgAMtstKkdjBWIyhiJy5OFwFoIh1RPRFpke8AvWCoYXayTmRPcU
1qkihpuzXDkgfI4Vo5An1dN8pvD4VO/wod/2dh8ehYJcgdnx8KAIPjXOZWO5ijPaSSt5BWMRLuqy
8UeyLf4wckAWpA+SK+tB3dJ6uM+Ih0RtEPjc9o5FaJVNdjuwe9fBmYOUaF5T1SPLXKC+aeNGI8l1
QaBaksHSJY/MjKomptj44MDkYtd3GRFYSM5kft/jRcoDilapzMa9RHrhSBZ7EnBpi+RthBuytNot
+9NYTOyJH0bbQadxkp22TvY8mAe1RyOZ6Hj6tYGWIDlNb8iHx6/j/Kryox+u8R6mo4cxgAPkT9CA
UZxSfLpCQUqexwR49eVsvXICKI8hSiWmv2Q7nlCw1vQboFMT354217rYnTx1C96DIfHRPgm+ppIo
pPVyH0KKaN8GacdLWZIivYhP8vLNl2WqdjRa/K4qzE2S/dlyI16YRWl/phzQG3hRGKqLQEGKvrsw
q2DT0hfJuEs/qaMFJTqRLep9Nd/3rjrrGr2Nf++mCFTi/sGm8EB/JMD+v0z1nTtURiMj+jitSHOd
OcBEGtx5MUF+218b8HAUli4LNgygCibZNMRGv08mMzW2K5v+StNtAWf0wC6F5pHyFlaBp37qTSw4
BNkeOsOaQTe4SUcbSHWK/eXh/wpbhL6GkYKj/5Ta2SWLurrEyvq5WJMd68GOmIeSKGNrshL9iLyW
DlhQZzDoMY2lptcKlDcfp97UTAZ8eSTObT9KKorXzToG19Y0Ep1Rm6DmodPhfbjc7uxNJVZHyS1z
uNvVRJB22oXvGTBKOukWNpG6LmnADj+pRiN2bZZgDtzLykHkERhh4oGlCFeaIlBACe8/a3hy8SU/
y3pyHGyyUymQLqdQZ310fPbkxe8zS6Ci32kDvCwXny+4fOtlbAWE1UsyrCly8NxDw/7j9438tDe/
vYlnunufcQWpl7FY8eq53bhmgYl32+qJ7WeiwEQNr6PXkXDgzFgTdzgCKA7qYGZl9nubNk/K0xJM
d8I0d2Yb2f2LWgbE1p1l8odfXlahSbQR57AX3XmmVBN+O7Q4mSxKkqEuEjay8WY12rSowqXCGZiz
fTytSW38WIBqyjyCE6Y5OlEOPhVeEW7wMlk70xhNy50oExXy+YO+fu/WQLW5sSNiXccgCxCaOO0B
eekuF0QXSJq3KvkMGYNoZB7lqSiZ3L3pWGuKNH2u7NWbUcbxtHny3FC2cNE6qa33Fy4k+gZuQQP8
Dc31vGs6aNerUsOAeQCxJF7zjtHYj2HgKwwW8Y2cKtI31AiKF1mO9M3jG0lXXXqxYviJk/hHA6YD
u6g0jC3h2mYpRSnUcInGMbv3WTV9wFIChvtoIwyPqbLE8zOgaY4lgcwOMci7F13csDL5ioVlJenY
J9rqSimp5gSUCG9hZCRblSeO7Wig9Ci6fc4eiQbJ9yi0iqjmUC3BPUvOg/nBmOY3y9q6rlB3ymhr
oS/wKLYZShsqAWnmVwgoVtJLsZuFGw1K0it0dfzQIdTZ0KBtyYjulFJzPBScTzLjABLs7vUo+EIT
zFO4id2KpQtogA+C5xT8qisXz2LNIyKzBJp7c//Yfrgr4uyx+blZPJHUKMUWWrjpmWfZzfSNxkhG
66irjcWKsl/6w/aLpqdc68iwlGyyyj/g8TwNdTHs7K/ua05OhYb3la7OhbTPNa1sxEBJflcHewSF
6F8vziV4yiraLemVgbzYvOiDUjrI2oWhBFLRHu4ql1SvFGatZgCicDWHglD+VL4ZQQjRNK2w97Ym
qXEKHtotTDWPpswZXOhWgVpSxNy4TH21pWJDvRg4DKKG8rwEUBI5j7oPNnE40GR2GcBbgA9cK0Re
2BoyhEjg5BWjEhDCpa/qAmnhdmCyYQXi1w+GAWBI4U/hOHiepWYmLX/Q6Wn/u2aRDo3VTHAPqP8N
IiSuoP94/nTM9OvrMEjPFIEKJd7d0TdkbDWF20jJViCQEW4nD8fChYd9hWoWqvoxw2z1/H2LM3FE
HlAJf6VM3mF3Q57R+9oxj/4X+uCyAtgcXj+5jpJn2Ez+2sDrRMO86/x7v4ss4SldAKSXI8L+b5SZ
jNei2vBNMVo4t5u+zudYJym+FSq5vO3BkLmbTkJ7SZ1T17rBGNcMCmmVUWoHKr5c/YbG9g2Weavh
qx1SUKHGY1/REA5R7VcBXlpLJ2lhfVJbmyv6F9ZEOPZ9CEBIlIVpV9TfvfAQ6RF2OjfXlopdaAFA
3z2BdjQQKdlzKUavGYNvPiHXlGT3a+yQFxkFwj7gPHzViNAbbeYc0yKA9vl7sU3hRg6ML3T4ApTs
jHYt6CSp+JSJNmx6lb0KM2yiLqnBrCYaUHDgJVjkTMxwC88TkM4zYJEA3Yy7W3kZpYXjqgPaibI2
MBe6wg+I8jQfa6VqBI8DZW4ql6im/AizBooT8iQahH7D4OQtlvE+Pq1RE8qVJWCvbM3alvUw7FpB
Lt419ugff6TMtuwzDs8wh2WuGFtYrgF+Rxv8eTwUJnfaL82YU5iKWKrjP1dQmDkYx1osgf8Vz/Y8
mgkeCL51w+o53gbEW81GCuJ8C7l2E7j8LZcI/D8xGlYU4oCootC16wCktv8kKqM2z0jkeFyEh1hH
XB+bn7zWlllfzSrdsBK22x5Az7DLuac5FutInOeC6LY2gJ1Zcc+ut6TPaXGhx8uF01TiSHn98D/z
RAOlG6LoXvI0JL9zZ4j142ln8WM8gqWVTktpuxCDqVTkSVerfNge/KiO0BQkQRmdGiQsYmrtf8hw
gULGyUXvtJfdLI7ts1qEA1JQ9cGAGODlUpZZoJhXWn9lWYrcf8HFG+JZEqfRAYAHaQtkXNQ6imMk
BEJmO+uF4uy8fP9A+4QGiMMBEAGcUuNgT3cmiGTvwgolzvuXhZP5kPHFW0RfnTOLUBjVj4ixmx2+
2pY5MEM51FOJNrgvQ4f9rwuJQMK4KoSldmUX6FgWIaOk9ta4zubUREnDRZEwBhuReUDiIJjnKqGR
d0u2KALZ8+YUNLci5hvy15T3tflNpaC/esu1r6qcmMa1kVE9DGIoFooH+VjeKzcKET0EU9t0QX0C
Pruwd4SDEnR9/DQVKQGCue8GBqlNEi1adM7NhQmnIxhD2JQA4Cuk0aWmVuQcF944N9GaKjHV6hOf
GT6iX1Iq0TjzW4TqT7rmLV8Lj/hz1D3N5VfQJigM5Ri0yD/UbDyBF4Dye2RepBN6vgCde3R6n6eU
R4qEaB09Qgjcs6lSx9lKkEdLDE6IkscEndRDq3RDabunGAuiJ2oJEaw56eanafMjN33Rm367QjEO
Dk9FCxFAl8vIx7sINw9ylfRXxSDlPOO00vv94IXfmqxYCP38BS0M0fnanNWEwi+P3EPvAU/yrGvY
hR652At1yfPAdt1rqUdZ9aoryezNTzMzQdoidYjcwZ2432oGaoQR8HkmUwtzAUOSBb8td8wQ18wd
a3ZfpBjgxJI0zyod0GUmX26ZVBvWewDtiY9z0N51Sq0grOxWdO3CIg9X0JTSO4AbITYWbos0LeBW
7dNERbSYJmN801z5zGabta1Vh1bOh2fAI7AUhGPQOnDCPC/nAa5T8iwBEIorzZcCwFcyWL1wpFJ3
2R7NHn51P+iHTLjr5VYzZRl3qwPD5mgYaK+0eGzI2MJhHt4EDxwF4KBD6KUg0plka4aEiV+uy/3P
Ee5ykYHyvGJIOT+6A4/FFiyWCe5DATNZRCPXPs8tlDwGyvhn4ly95xK5CaXjhd9AylzzdLkFrtoR
WxkmDwngL5VH1FSIopTRPH1AliEBP9K7VrjN0YjsGItsPCSc6yaTKoBCs9IPXwIDTV4QjafUs873
sxqqriXOGIHozvZ+ehRoeIIN+tF+mDutgW06Zsucb4CZzRrUzDsjHfIqUh8GsIw++7mYZANSw0ai
C6cXvw7NRP3GUqDmjcKbPOzoT+Xvu3izb4LkYR7S4tDhG99lWC37FbjP0FM/6/xj7hbqPgrSYWkF
yxyv6aelIOmPr9WU5N0QN4dulh3wII7jqyTZ4AqwMfyClRwjWu43ah684a6/Iq0aIJA9+QNcR0lx
hGkT6ac9DuuE4phDJD6CC808haFkJI64KCHAK663SvxeU/eCfSwbxmWmO9IbEbotxFw5VH7aycl4
gr7Jjs4UbB7yIdqSBgnl3MMPYbZV0qfpRerTfVi8bHq9vBKdTJoNbQTlfJcji+1h9itW6RvfVYzF
F+QhryKTi7giOwllbgDCLIVVPDfsJueyTOF61JjTMfj3U986GAaNSi85FCBcz/6JNkTVl7HpYvgM
r1rvweidtXvrarn4ai8sRKMANDB8T0xPVG+JdgA2ruAWToojY3rYpv6FWMTTo1HBBXFaUs0r7/IW
/RT9rSf6NeWEAFTq2RqC/yW5Ei05T8t7yhETeeH5PtrAKc3gI2m001bntOHMuHdzv9gAhWKOwI89
FZopjXztgJTsYe0yj41Q6UZHTQeCht8Pue7dTYX11VmqPCXMUk/slznL5IPethTLuVUQ0APGUsqk
DC3sDJbNigYhwAR7wnvAV+IhLm4DPFFP0aytblpbFBhlC97EBAb+ZefLCSBolvkkLAct4Ko2lSsc
+JKxk5pAnqFwUTGrHFexxHEoT6NKu5OJJ7tE+vcrDcpecjV/0iK+EZ8e7z4u4/3jbT5sPZTdkO1u
ZhGfnQUPiTjs6nVdDDj0u35/drdgM/hHkHxw4kE7OT/igWYGTWfHnzi080rqVJ3kr59ltc8u96nI
UnPhID9YrNrLf04oSQfk4Rq0vJhHYZbez2Dx89UPqGHahdm1uK4eGS/XpAWrUDnqyW4nednbU5nS
3kcDf45/YtFg80AAGT7rNU44pzUPkR9cHY9ywlqRtmY0uSWnaILhJ308XgZSUFBZhqqdNrgXHN7H
57kQ86WJTcawUnjEBSWSXffVQsfzyyr/undn3rTslgkHfi9HqTADmoQr3kl0Kqx7ZLCQjvAI6+dR
n2kzX3Vl0ABFIpwlmnoSH2k6VqCvINaURArHOhuIezACXEuKTXs5NcJYhL4eV+h5kUXs55Ugb4Dg
Jervg8X8qh2sww9QDWL4a0yCYMZgMgtacQoqYBlUmnExuE8aHiAGjJGDJMF73hTMO/d13nzQTshq
KORqq5kb623Fk5m5rILnNQxyQVZJo+EBfitzTKPf/PF/9rOeokd1knKX29sDyloJYj8codfjVFW6
9vcAPEIoZAqpuIeUC42TqkHyleuR/lHe6jWy2W6unNggssftw8v+KxncQLnaCbra2HjVJ9FNO4Wb
FRZKTFbcJMJTD1z880mOZwbXWCDCubbucIvAL4jOCM0wyMiIy1tWDHT8YUnpkVBpogfMmbxXH1nJ
AbS2rKhSzIQaTNAshsnJs28431PyehDSwgNpCPMOKt7nxIPCNfGTnPGVbD7MEVwAYgIhsgeFgYfa
yrUBcQNlO14fW5vb+MEYUTeQkEcOW8/0Oac+Crep5yPoavvpf6+xiqA9H0D296Ru6y048F8ZWex7
OcXuzH1LLvJY9fKnDZEt8g6hMxJI730EXx/8Eg4TGg0G9Kb3yGtVrKOlbz1Uu0B+X36y7Y3FWrUb
O4YSaS847Z3G/eL/imSkmewbVaErkqRvkfvjIyj3RtKXmA8609lS2PpUtxfWOPm0jdAwsV5ARHl4
8y6ZZZ4oRGqkQRd9JBCzY7vI+yqwlmOswGTdt0v1FraycOPwzA/61OJHvjtDRAn794fWix7qNskq
YTJB5albvt3ZHvOGtm9C9qHC2L3aIcqhS7UXj3ycrCEAZKZ2KSDM+kiYE0VaS3nC8ToIuBPiqkWv
4q2xMrdfFGRr6F5IfGGHpVU8gwMOQy2RKkDYcC/bOfuzEg6PCZT4iN7aNdaUIrMZwPYdRnEpkC5Y
dbNQqSs34fKskdkZjcS2QQz2OGifh7fCyKYTKN0NB02s2QM9cJ3IupTdCgW4UUBUpS/EM9PJqa06
VeKGdpjtVFrYjbP7lfn5JCHqqQEv7Cs4A6qKyNAt3CP52ArKCwlsBGe0cvATu6LL8kVYPQzTs7dD
RQmD3/vxIDKkcdtOuoqfyLNaqOE/45+3XAj5hlbHFxhp305zyuJJpmxqOaVa/088CBztGeazAtvI
s3jeYIDCeUERyxWwwTmxHl1aTT0BlX+RRXpcM6YB3szFlNNLpXN6lUuwPGUEHZk9MwP6eiBBJJMf
hcflhMAnVbIu++ikA8yo5PIZpNjNMetcwWSwmAyWiUs+3fkgyj/g/4681ChYbPyAOPv3vhhYuyRg
TG0SS0tYa6SfOl+JmnOvzt7kNAJLsSwSlXLzaXaEXSnoWqUzhYZC3p66KitCiYpNCLU5xKNcUFNM
vqzlUGV19zV++Wa1mb1pFBZWYbXojrOgX3iIDg3FRAI4xlNMZwYuwdZUwpCYoWOsih4zUZuKSrCP
fkaHTsnQoG4+p4K8B8uWiRcZIB9eq5jN9EHwLfN0sQ242/s19M3ga6mlpzlZnIRyGwykbH8xlqQF
BMygX8ejeQupsCwkNY84Unm0VAG9bhcI6kfKtLmxKn5NNUSEroqzcFhiNhROuE+eB9J56mm/l9k6
oks54VDCmx6Xm3do4klLyHs363K1VW+LK7mkI9e5uOtrxU5n3A/qvm+viHCvy2190kQXXR9L3qub
+DNdJ+gIumMtkEqiWkKNkZz3ZSBnjRuDZLq6topotMbpM8fCPW0RK453nCy+4KZ6ZMaPfCsvA3sR
xHZ7hi1xD1asIKVLkEM4buQEi09j3pHHtt9y4nmTeQdjDHOJwsk6Uzk9TsiB/blbWf28j6wBmVJ3
EYzWXR/zKynsCFxb5VH6iENGpGDIov0n6hjf4AkOqqyB1hh/AO4MD/qL6wvyx6ZNspaOHuKOouAm
w4jF2bK6o6NCcTO69F1vYz8YE0ptLv6WF3FThInCLDA3dLw+IJed+5DGk4vZL+4k4D6tVYaD5Lmd
b3uzfQQ7a2P/RGRX6GeBl0vtUu+BQvVLzOoBnYn8FzlhQKbcg1NPV6gFBIYK5P/7RSYu1/ptwm+R
lzscLNTCNGdSaGYAIofxCjIPHEeFfydTJUlWJogkZQ+jR4y/vuditO8xBcrVn1u4e+4YaRzjLemo
XQ+dKpQrQ/0pDWDGvO91mqqGFDUqFMkqtB18r7cSgHNa4PkbZkfSdm0uGjiXNbMgkvKgA+iUkTs8
40VZAdStATaAxCeJWAauNRr3w1O46L+EkFBRC+lHZ83Dz+LbH8UKahcQxRI93CkgMwbOnTreqT1J
aYEEJUHcV3//goP8AdNxHeBuglnnNqToZdKwpx0IYk0qWdPvx8EufVI+dVTVYi6RXQNFAe3oocCU
mc0HB6IAf1K399tlyFZFkwDeSAvYAXyw+49/YRBkxQbO878KpOVSWWkDDXMhDPtwFrSu9QdHtlOt
ImT2dugN9O2xcnFYHvnOETnPflesYOvXlde7oxjra+k/8fzyOjbxMuvIhxXi666lMC0rlPEXBl4F
RViMsxrRYRGdI8043nK03mtmolOp7ck/27vmUOTRGzQz7e0DVeYLgH0+9x9iLnrqnZhWzspOIhUR
dVoJ5U3u+bNlb+5wHyK/CTfE7pKInEt8rQSk4HnN0toQjX7aWC/luIko8fYI8PYm/lJbNGofkNke
DQJZ67PZivKCjCmV5I6zk8Y9p7K6eeCmf5dtaMHJutrc2/8YIICeP8XZ+vDZxXjeq8DchtAoqjUv
diltL5XMt3SU3+RfI4JCAK0W2a1dgAEO0GFKOrKb7LO/m/TcXeABeEd5n752FL6zkqQcGIpvSbYO
bR/5RXDrwa5iXXp8gJbB7Nl5BW96PXuznOhbQBYeKrkAO/y+QuEBoZDgJ1XTeyVfUpoAMtO/zYuB
+0dk38xOykXeRQArn8Le07BeE8MK/DSwE8ThHPsW3QY46ydfWt5ZMlpZoEByzXh0YJ5L2hUBA4xx
BV0GaAC0DMqudXsyCKU9YMd4ZzDyTbTs4HA8GUQEBwKvhqC964ySv0EdyFHb9JDMuQ2LHneHr8Uq
A6xRaEB5F2itjPQ9T6RjNnpVffRm/TPvNgxNilSTSM4u1t3aQBZagEJIeCAmDXsx12udAriqS1xW
GevidFIUcANgEV70pbzzdvkFp9QsjsXMpIWmKbLustJAtNsTFxt16WixTGMJvCTojzHklcYk+LPh
rn98FqnmtEORIGoWgCaqwny1fGIPmZNXkxG0X6iRYYq6n4a42esyJN1DaCJQVp9YAIw6/tDGh+F+
ut4KGGiE6WrHyo9WrBZCauG3CLmpsORUeYQEQMuGsw119wK5EIa2KHmjayVHvsvTIyRqR/u8kOjc
ZNp9nEE4tVeM7eJr4Hr/bTFDJEW2BQTtEbjBYx16XBzh1CudMsJiwKI9+osq9w2dhkU88kM/E6+0
stHCk/R+xVV/+DVG3XwgoUatLVbJV7finKJhSCJCOw2wlYh94ncTAuAuY7C5tnNobpSLc92PD9xQ
Xyj3SYjdw9bMJ9Ctcmq0BvdWiX1LqxkjU4AyyL/5TpkpqOo6CnSEu//pXY4+GP7mzx8gA4pNGI/t
ANOvPQSLQrIyJyX/uGKQHM8Gd8j+awEPE1B8aLtUOrOuf0b4mU85fKPJH0r+CxJtn1odQcjQCXSX
VktnvXO8dj4ULT3YVKZ7p5w8ipcLUgToBqEFPxzjsW2K6C1TU1xerfSWKgmJef9oeDXxBlrgO745
INONASLxn8LFbARoXyYUm73lxRJ+HO42qxKMymoxEOd+fbmA/nJ4wFFqJ7wnEyYI+3yJKcrlekVn
PdsQqN/Av+08aiktch2eguN/CqlLOH0uZIB0QhbBNB+tfhYA/8kxAWcGRoLm7i/GdwmFIPBXKj/c
1Swjk+Xjd7zqkyucvUTxr9iyXhLvswDhOjDMphZvb4LCmUSUtvfRxeGdDRQtJggpQgpTpYdLON2E
8JDf89kHHa1a96c7XNh02UvXRWYMGxJJrtDQEesfOpERCYhBauPRN6elAhg6Y66lad0W6vdC0e+z
OyGwr12lb4t8HyCeJBz57bziWFZVeJ6hoKekt5BhXFsELIogREuw0bUykbikaGPbQT15VrT6Zyek
CuqYynLqaPSnSndSS2fKozzReXAutkdxf6FVCPTezVE0kl1DjoxtD4LpbfJ8JYAzSAMmNDR3nm0z
5Kov7HphwwXFhIIN1K1dst8v49I22j0kioSYSqT1lc1eyEhZb16mDIGtXV7MWgoTt6An8PsGZ/WY
X4Y5mQMCBdrB0jHhXwl4/fNsWUeKeDYZoF/U4fu4uzZXoppZw1xvfdMm0Ip006o0q8FDRp2dIfzC
V79hEgJE28kgyCBp66YcoRD8KphDgDdSaBzpAnX5LpYKR0IlkNcJyWOlDF0qJooxUK947lKws6Zq
wfeqpgjja7ziRyrrEgMcb4WRyEemhONXBnwRK7fbdF2TClfYgHFYXbkTRuWCoBpmxQGhkVCfwZPn
s4wHSwUebUv2N/VHm1lWT+UlgG1lKBp6g/PPtnoaxt51kDmXty86oDYh94/U1nbIOKmmUBD68Gtm
0REew9t9p0FKxyjcrXHqeINL58RaPI1KHiGGwHLGRvpRcduVTLIHBLa5dUre4qexSG1MlUo8Ze7H
2w3CuyjUBn+ttkdfOL9jcShnRU1ibuPJuw4neCW8q1aXYgP2ljJe+fDmukTfyBcLmErMuvqQd+Rf
stRvpeLwTRxcMNrJZO6wsgXpAnY1AFH4NkrZ0DbAhv63ddL45nlcJMBw5FZg71ZbCATchwIRmb0h
0UsEJPylZtA7Nuz8IIVAd1KPzUj3hHqWuFTaOjlrd4hW0K5GsQGhf0LqPdNKCpFWHXFQirs+OqiG
aJufeaHKt5f29mGzyaekrb3f8N3bHJ5h+gczzk/ia/bp5XMtcgiXTtZ+cEQu2N/b5j0eWHcN22Pq
T+zMbTxneuiyglPDbtNYMSYipC8yVK+Yp0psvTOL0zH9DPOZJOiY3w7K5s8urnN5x7Inl6EwwmfY
Aor6pgvqxUGri/CM4OiiRdleJq6OYJN1qcGZwIgRjRoobiYeSQt4b1rdXMS18phRKYqgkpLRLcf1
m/lAR/PgHNbTqYZN/Fu7h3PTXIPO1EMVsZyzhkawzcjMLziA0Yf/qlZ2h0dSCG4TZd68e/e+tkU8
2UpuZi8XFPPx9ICIOqOKkFh+bg9tJOxBtcZru77pvaNkkkWIDe+4s5bW2IYPXgs9Wn9zy3QcB4G+
1wmVoxfptJ9Q/z/ula7gIyBhKZ1wl126j9H/OIDc1/bbVUwOxHgfe0fHy12egkGI0mKvIMHo8Q3g
edQCkf1yV9/fAsoIRf3z0ZcBVh6vciraTUvocT+D4HxH7wUpECf07tyP5izop6WwcFksuvswcLxh
akrcI+yQoNqveQt4h+5Vc3qaaFmSst1U3JL2N7aLrljcz3KRH8FaW4gYieaoORKqG0J2Ch3YkOdB
Q3tuBo5PwU1PAiniD1PxTKGnHxD4Ydwg9asMiUhKOQDmZ5nulbdYl7zm4HnIh5NgSqwEgvfw4XiZ
N6ZRSHOAWazm1c+pR8LavbtsZojOlznBUTDGJxPUShQkJep5weOJbM4Or6iHQdZxqi9/nuiIP7ho
HPauV7zKPneOxJ+ETOHecM/kcMh7nIw/UAFTYu+I/HFQt8cv6NA8T7gf2QD9fwbkt+YSf2jDEhA8
MInIK5A+xqhaqzagbXIMx9Vxp26FXRu0P6jqYi2MprgcIAEAsjLQkOEWHjSGwhX7+JoP3ycG9I/t
gC7m/vug/80HckHEdYgVUpLcM97FOVbwaOSckfX0+3G5+hdFbrsQfMPh4bJ8wLDABcyOp5zDh0iK
mTTvSVTp3vXrDMkxsEvcq59rA+Vw2vrhta57+8Bw9kp7cQkhsdGsxAA9CMbbGPe4H+kLPAJMKtlf
4LEaE6df4E+2a+8Pacvn7tChp33RyiL0NJD9gfExs5TUTXNOhrHaS4yohq2RRz92e65+H3HpGo1M
FO1yGTVZeY8NStO2bKo/QyA39H4EkYt2hzbqMyrN5QpnKXrjtfrW+cW7k/bQPGSufteBK/03q52J
EMrDPI6F+rbZXz9ewbgNXSrS1pd01cgu9wSKd8T2d7vs+HU0PCx0rjqd5tOfkClNmgR/1sao2YLe
SNGfVE54z5+Bqn6pXy4ygUxw9wVlWrEljnJVn2HhosaeRuDWmperdHM0Y2X0op5dS+gBtZ7U+wWX
Psu/QiEsUnfh2QrOszutaF5h2k413FbsqI+uDTBrjfMZBEII05zmeNjb/NaISMbDN1r4bkO+0TW5
7RwIWyThmx6Yow3W26FlVwhBKcl7PDhRsIEpR0wjxf1eNctN5+20UktsIgKznfmnc3zacD/B483C
hZAOgUqTP4VgFAnhg8r5hrSu/GK5p6SWzhpjcAHoHq34/6O2GpfUJyxUT4k4ZwUd6c3PReJUbsDJ
tbcFY1z+bIytSk+e70VDVkxeY/Y2Dr7w52gaVjMsSxaOuEFBF/gpsIN9WGQ8/qIdVyTwZnGp+ZaK
/X/CkEgbGhuhbIgb9E7egJmg/JkXobTFwcaeFflR+rWOLSYY+PjyikaACYD+jmQvoixQwC9fb0E+
Ai+TUqvzhorDu1DTdEajnYJ8Bj4+ULKaDrHP7UNgGU49Zkb/zI91pj5c4wMYr8YkbEr1AwJFSdQx
l54TLuEGdrHLcQjymK1w2r7rXrSlnZPL8fn4AZD/gN1p5Lvxar7HPQNKOupSU1g1EBY9jfDsVFOR
35E0cellsUEJvy35tG5POpT/NkoDcJUMCZtjr21sZU+2E9pi1pQnQvMyyxaRMmltJL3BXF9WvEi/
XdSrFqQ5BDViZGV0ikXDCw6gvFwAaU6SR4kk1wV0LGCWKYPH32GEmdsgn3hpZKICspwv4Mq5pW5y
vV/6cd/0ZflqPbF8BT0ldj5Jtncn3emyDLRbVVz1/sreCZtDFEgpxU0g+brzxdkNP2I8dmZfdZai
l8WwuY8ur5XR36cHPi59sqzhBheWU7WyWN8MM5vzdTz44BPluSOMvpFoGYnNHfxPXUpv5XfnmBZ6
iTMuEPo2IPzJelGy29ssko6OGuDkUqda3uEtFAMtmXheFvPMHQ4FRd13y+FcN8+DltOii3qAzRtG
UwduFec/+FQnf9wEdz8AJD5nClkvnFiaW19W9GDHDJwYPhxnC79mx8/fTs0guKLc4T7AX0VPaJMA
UBmH7rzl8TyWhP9fgqZzk+xMeItvZ6K0e0qshKjZcDwkK4bs/IXgzml74BZC9CxfaXLGH8kZQr0g
PFnwzqb/oI0WoC1UQS96oyeQcjM2OGxiN2ZsEykPKUefAmaE9ZKiJ6ttVg385S84b80FDIVIK3RN
5lb3DiMxVEg8HnCLGEOFTqw9w2Do1zAqHyNkMfqn3raHgxTB1B06xiYR1g4/ort/bLp/IXvr2ryl
NQTGVF3ebVBWXs7xwR8XMnxkj9gY310T0pPb+SzLxDpuEHJzbNvTOLCEPxORetSD9DBKhg2loy1D
lMdcQr98JMaKjIieVMtnDHzXv4pPZZP9C0jVkTkYpJR5jodoq6F2ZnZdx+DFKJ+vYViT1EJB/5FC
L2w9CUzd5rH2lXtnsntMeKaOQ+vLGHgdSXsPhJYmf0ShcAluDRdwQmfJ9F3pJJuYmiSFz9bSeqdZ
uyjCyyfzprA6gEcYQPEBNgqpdHZ8oAao6DLMHs6ngGkFm7SCl4u58xJa0gg911bRKgBiF6gdgP+M
MwPYuh4174MPqOcwoyvMZZ1qOC4yWwHOqGV3bxQpCbil99frU+/5J0Is8Odk0/MJm7SuL8p+A6i9
KrQc/WASAN1jOubugRW/2QBkFuv0AETks3KwG4bkrbi9J4GcQ0pgZTeinFTyeh+KDL1jlfqBi68b
6rzcWRrGCqFCAnZrFxztqlR2WNhLrTzbsFZGMNcLCH77sy1Sy8nf++SYEoCRa/gBk6Ow+L/+AnkJ
0m84w1f6j0D0Z5/E09D3ri0RYT5IoOqtSyxKUGqpJcVgJR6X8C9+RSQUqxBu0O1s8/Rr8QMQWHaH
2pKGTi/fGKZjS/zrgKiHrY002203HsO/htCjkiE3ANug3qkg7Nbw6RgQJRV+1Ngte5xFGvU65ZX5
xnO+KYr+Q1PGC2+nCQYdl4E2FOz0pVIrPAcHhclGROfg+FcNsWtsS3HetGOpLPS3LsHdwSpGulZh
SstpEtRCy8sMjFGl90d7fsUVglVK9FoxACR1Bb8nN20JxU6y2aQx7aQFmmy6667br3DpjZU6e6xe
KT27BWUjaDCv4EyjmJGTV2FhgBy7uiXkqbRBCqnieVWPwJ2jic353rlDI7ejdDtLDz0PlgFQ1Q8q
3Y9uhqdynw+0kEZZ5HCKBfu21k+9aQblvqmFKYykji4QkcsLc4vyEbHu/+FQ0NEUgTlgEK/c/TzS
BLczpOYQvUzrVB2DaKiL/XwrZmVoXGsIoo/L/ECfdqsTG1Ybr4y6VfIWUgidDoXlVrtgtC2d4SuA
/NqBiYYxyqQ9enlHrHP8RlORWChJip8ojG8RCEkIGUNfZTmdCpNEhBudM5j8mWWAnudVCKoiBu3G
TQToEZiCy6A6YRc/4IwhZgXZgEgmDRja9TmccqLm5N5QrSQOF7yYhLRtzTSSrh4Iqms76XFhPB6g
z8qx7vKdldl5U++3gUkO1fC2peTRfLmUlWcEDTl74KZrP5lNl3sAFzkUboJxD8Ey+9txEIz1+hMq
Vdavmb1l2/Pa2NxkKLxqRTNwlljsDCzo2+8pa8PRRt9R2hXnlGmpPQHaxp1/Um1XC1h7lYsDcYWM
q7nRNRA7w5DhF74tcylcAvafMk10Dfy4AzyocfIVz6+bw2mal1Cgb9mg2t62DCgbdxOPqUN79i/R
FRSbcek5uh4DGpFix2K04zlUb52pWUYX+S4g9HHOcZltU1zhtWhoyuY0vOwTTvNUCEFtpI1T3W/S
ge3/XECxFH1gKTh3PCHu1MRu7E56ah21JfNhHvBcl+RXu5Ml2o8mRU/tyYZJzMuX3xG8BvEfqpPx
sLFi74LWBiCw4DzFvsfcWUm2X12DdwDziv7p4PBWHo6KF5sDLDnNheWobyisDj8nIKGrp6brY6KD
TTcGiyQLGPeAKGuki4DAiMjfH/dhFl3eLFaLpjNxxuoCoULjzKwz5IUqm0kSOIo9JPGTNYCkTEz1
r6vqnEBb/RRpFZG7AQKxbO5RshVaLVFMcG+8g+x3q9FhaGLbOIfwTFhkgtrpUyDEwmKW7VjIHuPP
xi3WkL+HyGZmOprcSEw/EmZBpkMzOugT8kO95KM56y8RsFYCwxt4afP3tF2CAybDemNME2fZjMHF
Zbv6Qsy1MMHTQSJdReGLfoNf8NYNZnDpa6Wv0pDqhbVNUdXf+YPGEMLdZtd29Bp6MwWxcqeKY3ll
qkr/IFF0eFrlZoh8cr0/0fYWbQpfMjg0SX4d5JORnn0ZSdqmd0saq1rTyFO6aSNTxlAcUNgthFXo
4ky7d9TxoggfMQNLLAAiIK4IhwEACWQC2ecytQb53S8g3nEKwM+uTxeLzqgkzIQZqqzvv9BQ/eRR
ZWOrfowiERj3LYefdMRjwthuLtisjGspgnInmyOXblzMjBPKBk9iY6Te1ruFhEHYyPE5Hi3Lz9Ms
YossfzdVFM3vHN3HGCPex2aLBHDXDgLImeg55lYSR/qfmzqqxDTKnA5oDVFUTCto1NquEWOYcP0h
Iy00H0GSuo2gbW3MYZhmtsnZmHAqdDNXxgdGfy1v5yaKzcZOns7RjJ4w46Tx9g2SFBi49p899FAG
2jeydabgZO8CAy9c7xsvtuxNItVWIpD5o4Au2SPlvJBTyNiDR30RW7WLmui5Cp4i2y6ILaZZKhkf
+wtQuzl902b7QxibSWtI7aumuY9hEyw2So1Yu3WHDwakzVub4Xg9RUXQNLMsYnStM3an5MLpUa14
w77mGPEjzGjuvVCTdWa2FdKq+arJA1EMUFWTxiiU/b+4k6tXze1cTC4idxMuxuHqFaTj/G6wzsH7
S/pPjpe54P3xVbcVU8nTKDJ7ZpVOJHry2jTyR+yHnO0QBqxlcefq0XzT8N7FLBB7hBLojCGF9T53
YKlTJ3saodbIbZSgTNiiqPqaHI7TkLYPnmSY6jm2ZzOivI1OsBNDKfxpHyOoIhr3QS5Qz2FJxn6O
XIvQ+hTcg8G3BS2x3aPokuEOvy+m2KX45mMdv3CdI9HhAS/RwDNyBi5IMBilV6UDoba+b3fn+IiP
tn2E3rXfCKGPFe3GfxgYT4clJaGrjrWBO8ZUCX/Ewlx6YQBSGB3RnpeXCzTeisGbg/5ccfDzNgV9
kBMs4VOPCoWpv6KcBDk9zqnzAPZnWUtXesHTZhmH0DkXWBPydaOV+NwFJwAweseW35d53uQnW4T5
VcvhQ3T89jVE063J2I7gIf/1EtQUaNbo+Ku6j0Ts/2wnNurTqq3R8+/khZbW5MtYmAwetEJ5U7kP
X7qZj48EOdsNLujQnGqi9glDy5ySpNBSOvxfMhe0qX7bh6+ba3LCYoJVbtLMfbb5aDhh0A9DfGmb
GUpK/YGOkeCXr75a13c7d6pT9PZrllIo/goVOlUy7xS4a5TToSyEAF7vRO+h0zHLX+vjlQktHcwm
fyj9EAO+PZJHMbuJok8/pX4tWCdgGUkcFADk612FREAJ6Q7IZB5H3o1pSCXmsgeR0WPxVVxn2PG0
bSxlDR1malRG20tyFgXQt5NRiz1CEUFYF02OcXhoQpFwWJp4A3AkfowNq4ktbaJnqSZn89n7gCcf
ORmNxm/rAUjY+z5ROkaJ9l6gUIi6LK173FOdp8u6EegnjSgq6qcphM954l5JxAL1pD3TsztxQyAh
r3rQCsDwtRa7gAZcK3peCNKaVP5YOXJO23NJmL5w+bQ6BXTyXvb72FlzYVDyHYORBNCgsS+8VRaL
dC4ySFU6Uj+oRw3vL1/Y/CxzzZ0gcQ0GX9vvP6dtlxo2MOOcTcPNmR6bpgej2sm7KfbtTVU0zYyR
na0DcN6cEXZW2rwLMvwnubh6LdPAFX+vLP/jtjuiMNa3mrqKMCPZoLNnBK19Oi/guLh4+wxAzbdT
dky1wsxieQeKELuy2oq5Fi4/SG7sKZaBoa0cm0ntX/WnEx5Wq5dm3dLyVq1/56Q0mmEEEpjb7GUA
3juaUGQ7i6cBvlZW6Gnn9r9YoR04mOi4jJtm9ETWdr4/gIAZf8bhLEZfkOHS7+NJjVLG3e6huo7v
7cbRPZZ9A/3NO9FlrrmGwxiqH2vJbrkJa5Himl79DaVsoX2lg8sMYJrJzoxS8/IJK2DkUZvDatAG
FStFuJxZxf0MKehRXV8S7bhRAvh8ESBTtlHFMvzw/LkBeb3vzdWrWB/I3eWLzKL+wE3JvBeXgWSd
81mIDBEff28HW+wgOFlMQRdDdpS7RmqgSAFV2jGftznuo1JxDJtR28Bcs+irMDImT4qlvqv8FD1R
roLJ3MKaIaGo6fJGn17CiYCHuFwXQJ0ZN2ZNuKlh32wUy83KFYbqX9c9e3LWu+0bUix/eNl9+eCK
bf/oIOBM0g+syH87NuSt2BKacVj32EFwlWx50hGYwdz7AAkomWMO4x78CPRDitkZQbbzDr1CfZcx
nPt3/YQvVQlRk0FofoQRr9lp+qLbnl+bmFL6fAeY6RzjHFh0kHq2kYKLCAbKuvCKT4BtdDGJClb7
TKchg1LWTzakJKvhW1NpqKAWal3ZOD6rPbuUBJjppBdkgTSsNiZfoUK58J9Uc6ZzigoSZondeKaa
tNArXk7woe8wkhgD0jUADyefbzVbHKvM14VUi6LDYSR2fFV+U3r0docHLR1xBV0SZfGPZvV+dfaT
bLUFdCdib3Nxl/zfvYRGh254VReUAa74Szj0uBDu9DW/SEepYRaqYhWZSlKiXBN5yUpDpA+xfupv
UozGP/CbTJey0+2Z6Z9qlYhO41T1vvP3mCOEU0Lg5MmScRW93tfFgB7NJTPpDQopV5iuna8XtrH+
5DzIyCyRJ/8n4H6yNRTbdZZtVy71fhS1MwBIhlmt6lZGJzl3cXOccX2+Y5FZjCGHQWkVmxW2EGWA
0yn5hwc0GEpuX7JS346+JjkPtN5WC63Ez8dpMvTI4vt6HZfXRkE84ZGvz2CLLVnXWUW5PPSv826p
AgZFhcQ3HbWQDJt0az1GPIqlAToY5KOUCTu5XasWI3VGglVq6iiHTCFsKAvtxrMNs5Sve+6DZ0hx
jh6qOOma0Ag+5iPbU3NvFfGTq8iUg/xYNrx6sZsjxpNZkHt1MDn8VdSZq6lCv9CeabohZg8TVrm3
VcI3JwsQsJEcl4y+IlGQrtv0QbutgnGdx7Z565/D/gkIlzFmoyVg4fHXybr0PGKmAANKMovubVje
J/mt/JeGdNrxpq7CsuLiPdcq+FNRzKNBkh66+ayWQyPm7Am/cvOaqVVfEU5Y67/CUssPFCkRyX6e
W24K8Nrko3StZzfRaOav9B9IVMRE3KtXiyLITlmCwFvSgZGfO69kOlpqfnYBwWDIccUJYqaEstVB
zQ/OVQTm6OC6klXS16LypBFYmhuU34qSi5YSOLJ1fUbaFZ8Qh0HbSLg+8DLl6r71gobdo0NLmocX
5OrH4vmilpEwmtFhGzazZHK/LFIGMBzT2HbojsjfhcAA0XpgZzYB4bm2VNksGqon1D5aHiJhdfWY
4PEuvHiu6tOHepSIZcAqrOl+dSsKtx//LN2IL1pcO+aRp/tLRbe3QtV9Et7YXBCIlgZ0zVOSuAe0
af5y60LqIbY2NRpaegxiZwHW1KZZA9H7typ7Ld/qJiEkn+s4tRLDbus/aLqSpCtMV6B73Ni5eGm7
bhPLZ/zceWjNaHD5yLxItgMgwmS8MBWnqVy2IZfMylcIJYHbeZ96CfGsguFt3swaL/C6xMVGrqGa
C1KQpriQa3aDolIdXXn1DSs/gkxjkQyTA3vhQjkLFF73w7VWoK5q6FrDJsYJl3DqUgfghpMxipjl
pdBDAP3p3hBptEFCQSyZ1GwwnxM9Cs5J+ojbbmkbb7n4SeJXcG/wwXPHw0BDTCiw0w9q1Ga/O1lM
94FjL0BLbkD0eOIqjlb7WiGFjVq32Q4+pMG0VQcvUc7cbPRfsKmRO+mEnTGq1+nEJY1WsjcoyCEN
Fu9mMtVybLSznEOJZK69dZmesWDjlfA9Pt2fyDIdM1YDcyxZMVvHlaxThGzM12YJJBKWrsBbdjo1
uoJvtNTtnhrfZs/Ij7RDRkCswJGhtfBVgtyNsFAki8hiqdqMPz96VJCbLrhYwS6Ewzr1fCz9Kp6a
0Uu4Lykh6UKu2GfsX6U1gQYRf1bVDE5V+gfuTo5eBAk/KIXEHvUf2MB8bJb3EDdOk8qOF5IcgFXe
RujIrYP49yWZqDIM59QYCml07P7NBxBwmDN54oDOhubb+i68u94QdoLIG0nidFvRV3jpAOZpqxPQ
In3I45w9OBbs6KiTx3Pkpxqv9nStnHwTfZjP5zpWo58KYke9HGfG2bCYh+Y8c5Lb1UQiIcJV5Lun
lDm/rn0AfX79ZO7wZT6V6VN66gCFpfKrbXUDWTJTtKTh53ml8+kdosX4dRCMrSF+lgbwIhOsNNlq
ceES2086eOZPzEJ0MKPKNytyT3k/BNrrO2bJhwcLbxQU3Z5qTWUYPluLx01vBV4VLC51KsaopIFB
dnvjv0lvL+u4+psv4vMIJB2y9ws4NSCjxQBVW9W+Br8Er9iQDiBYWfdugepWj9PNm+N0i3Z0aKX1
+vN9wzTiQTM2UUUoIrJdjBMnvZbz1g768ESvVu+PYPL32XI1TgA0O0q/2rkXRf/CustvEpJhDTU+
59Fu6buoopuvhhQCCNzcAc4SRYCm2mvhSwCmt7QCSzbDlUrzgu9tBpoVOl2nnv6ynWgCHYhkfQ9h
hnqnlUYX4bLEmRtXYrRZGj0U5YkSk+7JaWsbukMaNxKHikqLE6zbKd8F4sPsMK+wBhQS3ois5EDS
2Esk0Z2kEcXo+RV4vqPUmcV69q4o4WGvTjAd+IMIkQsEvjG8HmsVZNd04tsdCAqNhJ6yWri4uMqX
5P6kXyzC6YqjF6ePS0IL57llv+Q/YBcwIytYV/dKb6zrnWcsXHWvF7mcm4oeYvripbQRopv6C+vr
b3wmjaKutx34uuZ9D09pZNpTjelkwrn+xNykm65iHcAmSRWUqNQvNWdAZ5B/74UuAGaziChok/k6
Y9mOlZ+Ot+q8+nqEJu/CpC4IUr1YY3LyCU2RnlHSq02F7cAszGolyzcGESIXzbEfspsMBQAYgnK9
AllNZIVncIw30SQUaRxgS2uj5YVgM/ju3OpOuRYkS5SYv6MrxrQPoXxMqEJky4/n8nuX9JMCVAKB
Eptm33ICVjaBYhjt45eIWwmjCF99WYsjeLzfg1fGRp+3riyvnSrIYiPPmvq3YIX0/yTJDktp1Vx8
1xI19i4FucKddYslebNQ0vh5vTj/cdgPcQn1fWImF/S0uhSIFdyunq8d7kGUjt+lqVd+sD6Nt7kv
KPyfxG0PDEmEiqqa+JaaYSJ7sWTqhi2OKH2IF6hTEtRGq2aBFIy5bHVBfXg/AQCBVQddOWZh2k1s
aPs0wYmf1EGaPezBEqvVDLtQm7acCms+ByOofaCyFASMJlfTX6zv+07cNcfXSm3Fk7/FSjZc69aO
PR1A0KbefgZ5dqGDqk9fpFr4K2A98M0MEfwxGrKYWyeimjea1C2xmOsDtCIF9+XoR/u1jn/I7MuP
fqzw7UGN4eRl4vdofARqtqmeqLSA+3GKH8d/iAMixtreh/xGtkeBISeV/1zMxFtV4oPq/WT5oBW/
5CwtLFabvJl71lY67/ajxAmvZqYYE8qr6zRRbmyKChlsr4y1R6M9gkvn2azCeTN6PpOwL3d72ciR
/2I5QuRfBfhFc4wE0gQKZZ+rBoKlBqCt88knt11lRxzYoByuAmA7l8eRxtNqqPDQE239+RuPeqAD
AAfQN5KyJULbJ73SeyOQQ7s+p7RTv6g78UjokfaEKd8xUMGGLOrHRpFWzjrYR0YppCRI+OVKPXy3
zlS4ueqpYhFkidMk/8zpMttFiZma1ELKIejM6V0XPEO7uPyt9KqTqO0JFyzhzQ0C8g8k604vlEk5
iivQbjrtvp8LdIoZghwN5Mnep/5LS4V5TPUQQF5rBqOSKhM0L9Tz9BAnIoTmhca2NoCrSG3RA7Vv
8TYHwU1Y6lI9669hZPW7N+5tyeiNSQ7z2wCtel92xkDx9GqucqnaqsN4QKltpwTO28hFzRL7VJZg
LVVyqHj9jsHpN+fGT3aZrvBlMnz5LiFttpU9tQhQCRIYVny60tmxQYOUmYf+Niwc59xYD44lmoi2
BwVnW6KWW784f10ZlUrSfn0DB2kxl0vsycPtYsNuxpxOCUVVMqFCkM2NywAV8S3trEMAhJx6inIo
8YOYrn7/XXyGn37INcqiy67G6YGSWdQ93Ztlqwi8qFHBxm2IXR+KnxX4zTkqjaKwR+oHK4voHtxN
VuhE0Ou9BYbzmxjBk7ShIT++6QU5j2hi7kehh/d1LD0BT8uoWD4tl+Q950VKafzcZ1rWxgU3Dh/w
7NdEC7lAG8MAfeOKwra/LJWDBdFHCYb4QU7meBGwB2S/CFI4XibUZCO/1nO6+iSLXDK0OFok4wnU
0Jy1brFM3WwVwOzwSYd7dVl/DuciUPoqX2mChar7ZYKicq1FnE8RoDBLRWwF5Exzol51SLMC/vMm
p9j8thUcIo+9lMJMapMkR5Y/0zLq7gtcIxqrPPGeuRmnkQzfOEoU3Jx8HsM+q2GOIB/80XxVJ2TP
fJj5h7rZb2aHmX9pD9Y5O/xbg1ytef7uTn8hyRvYfoy/MxaywSZeXf+PC8FlZGPr2RZd2EkmfLpT
yQ0WvWjPvurN1WNVd+uT6BfmccYj1/2JMPbnrUZl3j0EtP5+jrB5zRont+iIpUofc+WRq/tTdKi7
XIfr9tQQ+dXFt1oiyxh77OFvfqvxpIHU+Svuwda57HnMrNEdzVJCk2PlEj6D5gUi7NP1DDjJjmBV
mHlVcVq5rHrRi929fg6AK9fsM8FVsaLBMt0toB1+3qcSOi+Y1K7Uc0PYTE9ksZAzyBjWW++x7gXj
Y+BNZZO1au36egEgYwOhdV25XFAu7YxcY+uxdCxsbuENhxANetOjevLx5twxvL7Iljz3YozNWrRG
wGTuXfErIl86o5WZwuYpAJTRKS5wSeONXJ3WkTBxoh9gAUn3L8VYjJj9eahMOFjz/fM1lZPH99qE
RzcXJpfWudsyrudf0D1TCIaW/JNwb1y4Mqj2IcJk4w03jkvbklb5qN2h17cWusSjYLquRk+YmGmL
pRg1ecz+DhuOs1tOS0JOznZZK47n0fJ6nA0w15mule2aLtHQLHVNaMLDTKR+2ly9JO0Ja6nW8BFi
GjJ6L1pVHmedI+3SA2KxlPdkVV0XceVoqOpYnJaIhobAUgXqSLz6/hgPxJT0tSZaSQhxIKKhkQ4D
fW8GVuJGhgB2c9tZoXS8+fDz/hZ34qf+WOIiVm/O7TxzJ5sFMbr5q9XNJCwP2DcnEXjNAxafiCj9
Y5L1GQkrk42qU3rWHLv307xHldkrSuI0Tn23T/XyolsPJGsEeNFWLGoVvLrI4BPJNPvAdnsNx3sQ
HAaA9UpSg/5GeO/i3Wv0qHnKwi4Muz4Edj7jUuT4v4+56ANBoHg3nK0rlyUUz7ZvhVuYZRaKJbg+
bfvBGwDOm6StcarOgK8FqKwxot92NYUgFzLmB0X4Ag8VoBAQ0DZZFAwHLgh2kCf2jTN2jhWvtZUf
HteshHbDV/9Oek/KXvZYIOzodFMDYT6NpB12zCSgd0YhL8VYTIGIoFL4GCy2r60Bri/shVzZyxU6
wxFSi7VH3xt55bjq+FKSp9DQ+ADDsdqcMNsaE8q35St6WLlH36JbgvRSwKbH6NWwR4duDgiS+bx2
5n8ED+VNAPsTBwxy7+nuEBhcyrXF92ahCZLtIOdT4Ro1OgYvbgZEWPaZBn3TrIQuxtWmhmTWqRWZ
cv2XBViWg5xBTADVNze3HjUvkfUFL/pbT9rJArCU2UK5YoF6Z2CYz8a4vAeQYyhlQtS9/K0QO0DH
kpp8kGpxwFMMzk1azdQ/v9vULEjcOxB3+mFvz1X4Zd4C8JkHAXMWlFU0w0TKfjIlMQoNK1+CQ/EN
JRvJpkRaKfLfbHqj/rDdVm2/Ugp+p46c8jizs0gqchMLuD9cadDIXSL5ik1+CG8e0wWQjf/XbGer
n0JLm9KnHcXSaTQaTCPXT/UfoqeeopRI+fDNIKfp34/mgZkrvSvN7VeSKg0B+t5FlBUNzJ0ltwSt
FRaRS1OsT3hALQ/tg7YRN6UzfLyfeVBknsYcjKFPQ8lZPihPcFFCiexM9BRX5a9CG/UtVdqOILHY
ocngf0t7FD5QJh8JWjeeOofDQu6Mpyugm9R9vCRioEqIIkjC8YlsdhcZe09G1I32IpGu8bDwuDW1
fwDcY8yfjqiuK0m7crfO0UB+/pMaEqRNxb4Qnpbf5XcgYhOOglvecA0XakQXAVueB1PKFIjaHUK2
vETtMhOwg0LWot4gO00Zd5W/PFwj58OBVC2yGvLy0JaFl+nwfQNQ5BoyP/tC/RgMIpRuhEpy+fai
OuVosZbnoUHk/JOYfjKeGwpTwJBQNHTpYdsDd0+MqQHYzM1m5zn+wQvzLUZfrJcWG1w/62zCQhYj
I5ovPlvY753E0rMegwOlrYwfjixtp/D08wC7VD771jpDsaLU/+msXrOApSgqlrn56vcs5vGo9DiM
zGvqid9C2UxBooDwCMr76jn6m2XWVksffEFyuEJHME7m3DvmVBwNiMqJRWRA/lehiRK8yhS0+jGj
9OQSnV+UmBGDQv04eDGN0GLm8JQx1HHn4+w+SP+UTuFlYch0FBEth0dgrfWti62J81moR3/LRJOf
BzfkBlXAbfQ9PTNT1k5suNgQGjhrRv0jLGp0P0FPxbe/V8PnDiHGhNwB+sc3EPmlA+vce/P5d+df
G1yOMV+rGlQrXAP3vX4YkEkYvp+vsvaraKlQ/0Haxp4tIpsgDO/XDEEPMfwAStFYm0P3elS4fVEv
fULy3vpYBxBxVUXnP0j3cgZDgHxO5Jyl/dptB9knL22ENoETL3jL9yYQ5DgaiRWg4HNxfFEXoJIH
CP3MHDK6gCb6SK8JYst++OFEFun5GqApukOarUVegRTJnV21qv3FbFrwxbj9IEU8CjaMJaMyED19
rO36u46r/daR0zl1xWIVdQpohr6QWhL3CdFl9bHGvXrgUVWxbDWUXvDI+EizeVOKplrk8vYY4+GG
Q/Fa2q4hSOh/6OdaUo6JG3eKUSnZk2OOLfvwLT1ti3waJCuwMYg4Ei4S65A6ybdMDGiwJ6Igs4p5
tltnJ+2OwPWOmlxGFhTALyuAqy6ws3Lql+5pEv/k4mUYoTvIZCjAuYVKTq7SpJITDv0x2mjp0Vhj
mYz4oUI3WyUGQP9fHE0xWjRRZ7WNO8wCjgPV6YW/IX51cXBCK8bdz483gAqONrzJqcU/zpPDRlyU
MISQye+PHEiIosdjrEff42DybYc5qF3RaQYz7825p3aP2wdNT72gA94nYMnI/IWvEftLkj9fxNye
fk5RlJKFmFV9Mm9yRt2HCFWbbtNtXdWxUXnwSlhamYC56RiyzatAwFvCeLvc2rH3cOBpcMyyv2it
zD7KcqTAR3ggHgjHayKiSHNGS55oLxebaAIBrdBeXzJFguSA9tXGJVYvl7ozyyy8+KVdC7Fsmnb/
ZDsA27leMcAt4SbtXejU6MHoaXFE7QEDk7TZEw70ZlUli4jR1eIF8Q3g3KASjR6yESBQ4BmLkFFe
BWDcz+Mqx1n9Urv5hwXjR4z05p3FYphO4dakXRVMurPuDJ/ntTB+f6JRfmSJMxr034LfBmg5pd2o
8MvfnrZOw0yEW37wLAUZPClZJZxaiYDgLA/6x8gDxtQGE8g7ktdB2t8kgihaY/ltHD5M1o1+jfDW
Fw9qXCAYL2hfjjPHg3Gn/siREzKzNmJJsDOUE3Q0sPWZzaIBGK8HUB6S0RMDg30x31WLWPha3jMZ
zk9TeB95HMgBp0n6/biwuU6Ef+rTtFi5ThqvTdKxx0lheKYRtMmQQLyL8t+9jqOqzhqoGNVJnnI4
qjjXhDSedvMYNpHG03oH7d76MsvWPFididu9XYmRp8T/oKlT427uB5AK1lV+cf14I2AA/LE5DgF+
jtQeVgEbEReIpQYB5oYdjwYRNQvsD892AmB19PoxX3ddtkQMubMFTqI8agJAzMI1UNUWSQshXLXP
V1MXI40v01oRN52OZ5+XMoFrtknIhittJUibWuVnXHgrFrH3SpVcHibSs9rQUIldtAXhKmKuQY3n
n4oUEUbCDzPVuhTWvQCKn5b5wpMdjWlVDxICT6niQ9gHC6IMEAAD6+IztYEZS+IfBnWBeXmcK52G
xMCE7A1CXCuhD1VJ7F4wMGecFskQB8CAWpKFRoM2FIlaZ7fy9zUKKBzunT4VC1LwExMBPqJKKZaK
m2vzzgrzXiNg+cSEY5BZL/A41D0U5LmqeUOWWdXAPDXIXLuVigW95C2y64vhTLFWDFH96wcUsCtd
xveAhtPSACdv5WTje/Hciz+GEli8Up+zQFHnyCH4fUmdybHmU8kF4xVrOFlOQ/QjOAZSNBr5j/Q0
WPYYw899+X7fA5FiDT9Y+GYNAk8xOZbN7yU/JoGXjhVmtbmRbd6KWoMNCkMeaUWi5mOA+qkgRP71
ghYYPMYC/JYDXeIWb0jZb5ufjYdIrMr1+crJ/iG3UrdPTW3P/dapvHJLQuipjmolsYkYKuHwOGwV
qBfSYrTu2UVJ1VlyQO2EzfzXaQIU2e4N74QEkLgD5CQ0rR9uzazTJyMvCLoiLXFUzFlZvekBBeVk
voGtqhE4Dea3NS+16vlnH20SiG7zrhIwdCa3+3WWLk9jlnRj9Yoca1p4c4atEgxoas1Gy4JiGpcS
nr+hCi9RExMuf2tpcTeCUG4Mq/YpiIFWSpOLevLQpFvGC6rmeGzOCR22YuHOQatp3NWQxqmrMjsI
G47vxJhQUUSAoB2CP5R9wcpn9C3qTRd1Se94q9nRD7iMuJrjc9UyeAVDE10o18EniHEBA23HqYoH
b19Q0SX6aouOZXTDgnPjYdXE9ImODF3q7TC10S6bvW42Zx42uZK7AsbaT+8uhlFtHh2N4mJieizJ
kR+TfNczkhMiCRNgrGVNkl8GyuBfAraO6ci7f/OoB7mqnzy2N5odSdv3KXFcVBNGjyC00qmyQNQj
yZc55QpGtIzD1npXg06ihEy7zFSaTNXvIC+iI9eA5nn5OeCccAfSOoPFbsBjRtlp6mtrVusYHitt
qI+FbrCah2uttJ4NetGQfa3fIo9bUnGpUBalxIXhk/4Fp61PtEbO4Z3QPfhgJbm+6hPqKXvSIgvT
84s7lKXEag3ckK1DDvQU/mKJ1mMlY8PbyI/+e5S90XVI05SvR+D2wHSv3B5z3IIVWZeI+uW7qfcb
FilH4D01BL09r/lzvGpzEWCKJLib4RS4THi4NLpDt5lPu3zGSJeCCf0IFX2ZbaigYURQYqAgf3j2
sXKvcfr7CGo4vq70TXoF13nPiFZkQVqidmCfSnwBI0ZrW5jNYpGoPkb9ICib98XMHRK2+HjH3e6M
aUJwnbAEKEY7e8HcMd/yYaj/dkzYysEG+L5FO/Bvkn9LymRkwfaAscuslEykVgpowZCkIcLVDF+P
TsQICbMSpIN6wAQmSAK9oB33JbcnCbWpstjkgOhjK0qmD130xfNVpQt70dZGMHSCqTa0TbhDB9ux
HwdSsYEZNkoz88IvfnN/18Eerqt8gMV3bHEKGG9neAnMSNbQZe/drOZoHwTOWUlVJ654zkA9rR6r
F+3fqb7l9eb2Seaio80Cpwe276s0cAbcixOpsgJVffKpHvi36meQpfvNV91MI8Ge/WPxCAL/jlUt
msnZGApr5+uPHmbkau3QIYuYSBysJSxPCrYEjcPcme5LigAzYfUiM2J+gts5XnyNXZdZANTlJHNO
wuvigeGrfgrr/87c+KuSRBl8j/FQhOvx9qelDzWX31z+xuUGXREcJ2sknNouanPzFkejOFd/f9cZ
goOMVT2anHkLwhg11bVFPaXoqyeiylsQSUBtQdOsjqA1xTrfwC7E80Sm525OtRVM4fN7q0YgX9+V
2A7zC6MDEIPbsYnGiXie9ybKrsCrSBAJD+FWh2urTdj3ZkQVbidRzK4JNmaC5nGgF8xgqtSPhNAm
kQ60J4QCdcCRONh5LxCDK2ctssPEQMAzudERRCmPpwrw4Q3j+a2LYN6WBbn+mo6a0+aTIL0xFfMP
7Q0Y7b+eg5weEyAYE/dT8v+YF2aTNtyrPfzIstI17doYPT5SfuWAZN8J0hF+IuzjbFUIqixTX3E7
xroMTagU2oBIOY3dX/XrJYrfrUzCKK0B0TX1oVG2WX1Oe264KgRBmabc4kJiaNfPOANe+iQ7LeM/
+9j1coV1Uhj9Oq5rl26uVxEoZ6nlR6Q3I+aJLxt3LzxQaEbxalnnEs/LuGdWyNZV6d9m9GgDnSz6
aPmSGM5wITOFXMLjrwqg/avEI5GQyD6T0l6DHDvD3phg/b1NrXEbYP+JufYWp8tPxwz22gD76VHL
RU7BY1hGhJW1ZT+/wj1iUABdRwenxjoRrtVG7Omac6aDsQiPhh5bABuewJxo1RYkE40W1s0nz/HR
DDxYcNw3YUXsQcapserZu5q7Tc3kiWqma18jJ9muoqKDrRCUIW7V20tOdy1LQwVi6TFKY9+DUbgP
HnSQY6WnbX7VHOD7xHc/xtqn5UHFLIK0EmsS09kWHkDFcAosmSawtim2udArzfF4KHxXc1hdITs5
URH/BA229thAQx3RQCQTNcf8dzIfA245reHDfp1qh2081hZDugOOg9hzFMRCJLbwc9mAsjDsNWZv
hJZ2SeNfeHJ+86FohVvwhYo8XA0OukuW8k8bjP6LhKQDVPs0sYCbzO1KDi5i6H0d8kgrmmzkzlvo
2+7D0YiVoNzBJ6lLdxbqDqsWAya/xRcBwCvJKt60BXGK4I/O23w7nL0iRJxET/CJ1znpdvGU8fNT
6GtKJkyGLxGMhzR0n+EemQr/kDBvv2qGrYT1xyg22oILRVdT7JQng+DMWUiyyStGujJHuQxU4lpc
zaLaW2yp219Cp0U03xd4SetzyCiivn59tq6e0MP4X65bTOCiORr8KRMF6KGr0n6yycQhVXPyrv4m
aA+hanCB5tKfScCBI04nLb6Jo9kCQ/AVsMFIAXFaWrvqLV46bQxNJdhy2iInfY7K1/M6cit88kmh
LL0kKJYFYEcuS7g9qSS5GBHcwXkN+Av0ASw3R2d5Z5P7C5YbFNm/jmkpUdA968gtPF6QKTYGoXUc
e89a6pzut10MRg5zCxG8bGNcT09LIf0ayyraeqfX8MiYKLNkoCqg3f7XNTPbXa1JdWikvcvUo0e8
HC9JYS6Z02QqMM/JAw3qnuxRVz97/JyGYcKx5stQeF1K6x66RfLPqVxb9XjIaEOWYkFYb6NzAPlq
vcgKN7bb/Bth+U2eNCFfKhtdTYPakw40Q1AKedidfFka0xM7/eBaHgUaGO9DpSr1tH4FfowsEYuj
3NfBvBNZVsOpqETQy7yEXedHZz/ggSIVS1iSwkAuBgVXG+3CDe03SaaL6JfDja3yGCOyMc194vZW
qYswzGfGGLXiku4go9dZLriBmbopgX6bjlpHRkzVQNKCYI3QAsHAsAeXri/JkhBE2mAQOJEHvey1
lBae0vYTbAv2TbD0BycK9gzI62tVKxtRuQM0f2/cwz5LGEHXSlJLEOfpBtmI3r/h7ZgBLTnCEUX3
j5Y/Wf08FfNTq6OQI64lO+JyAhUtYFe4Bvj+4EFJWk5CqScZEIDwI7zshWGdx3T2goE/6G5Cncb1
wFMIqgzhNhK0mHHV1eb/1WMbWgTGbBoh0YypnL1Rpy5wi4UrtbSNpGTcX7Rnr84RIQTWh/F3/03h
K1Q29w6jnFd9a3mzby3vQsxjDgs1b6vGEc4S2pUsbmuW4UdUJ0k0clGTXLKaGCbcrdjeG+Ogsvno
KvCFgo/IDw4jfysYhplT960Kwg1+HXsLd6ROFILSm3WVPk4L6myLBgTVO3ncoYmxOv28p4gMJ9iJ
Lf9ptXP9vKJVIvxB5vC5mVM7V+cWLihEEhxrHX5Wz+2G1mKSSBo4AXbjqw6Ra8FZBs2NnMa2urdI
r7tklUSUEM71+q3yCuM2mO+zEvxRQ+qQ1pMFO+Uq9vEtJwXkCcydtcthiBi5d+lKym4+NTpidB+i
lVXN2uEuW/wXdwtZdMyaLUVqSCqQlOikyChokKeE8bRhqfOXEjBNfyTTmgtKaIwDWusebXMoRDd+
0IgVzV+czZK2IPrWrf8s5SnndZU1MpLpoq4KXfjYuUSlUWqGVznsOL4Bl4R2+B4MHhKHcs4ktrc3
D8lQPCClj+xY2Wuq9ZQLvyfoIVnuJwvHmn0DoZC1wSaFS+NmIiDxXFnenKExIVSW2VOFFvpYRuZE
lL2D2N/7zf+uD9w2dhCCZcY4bLHcFTTbOHOROoC7zo9ATnGV5R62nLnAlroHsCp+yGfRvpmb4Nmg
sAMPG49fGk3hnNA8YFsvdGgiDQQwrKRBKuDlYx2ugzvpTmJSXr0ehHy4+T5Pa96v7+Kg0lPjAEX9
7J12BJjV3MQjpbbLcMRk7Qd79XWBNgreSefKPkn6thb5UtHrJy2SV+ECHLl8Pxp3zplo+6NMkIdE
XeLx45P3p8Jm8l+ZdNq+ugCLqQ3gG3zmn6laojF/eQzk5gw+vuOvz79lyowxi4ueBi7XZfsuzbK6
xs20xoiGwJI85MElNgpi2Fvf8vmewaIgnTmCAzTAzitXZu9CY6ofh0J/mkmK+jDEshvFNk+/cNPg
1j7/OJ+X6G8O3CXUo5ZHaef42MbgAQRoksEKAxIOzP2xaIdnMo5dOhWVYMasKS9vXco9tZcW/04b
2vyEQue5td5pv58/6aVOubcSAEhAHRFqbGI7ymRpGMzdZ8iqKcfAyHwVaw0Zw+DeVoUU++PlOlZP
gDVkhpFL9NMq79Is1K1vxYBtCzcbIW2xXX59Qw3USZ2ll/pX7OicY1efyN8KP9Xl3xlmPsl1Z1w+
Abr4XNXGDhWmJdrsHT+4hTyeLEUl50GeyZUJAqT7LujJGQKAKsgcvTeeknGMTpPLbBthWUYD7+jr
L8EOEmxg0PsifknNyxXe2yS5+0l6RIp3r1D42h5wkOp+pt15sWW9Q7uxKod/GK1asT7VcqL4eBLV
Re77wTNEeGFOHjdnQUQqLAJsjcCFZsEst4WyWgLYXWeOUYo/GW9VSHcyUof8kQdbKvWvwFjHtZlX
yBQu7aVocfuAAbnYlyLVd8k6CiQpD2grfgZFO2pJQ0rYmxdf8TWHQBjrT8jlD9mjCrMt+Ch/nuOQ
sZP0O5zHNXfPwX1OjppBtuaebwCstz9PSkApwyQEphZQDnSigqX4tTOkEq5o2kYjsU0dMhLrqDwU
aB90v0Wd2aSfeRsK0s9ZdW7Ot+ooC4IuByi02Ls5Ki9UnKAn70W8I/nGp6SVY5BZighPIUH+yrzf
exkZVqKTWXXZNS9OAE4pP9p82nLb6k52l9MsvnP2xwHAJw6JsXgxp1uAcZxRspSr7WASR27BKSYP
mGUYCf7D8PZIWciTIktMwTTJjXN9Dyxr08qYtJR8R3PQtfQAPtF4zd6+R7e8+DoBszWzBPz02iDC
AED9moI3ptf7nXc+hSiC8I77Ys8YK0WKZKFJ1p1BspNFBNcr6JgO/Ac+aFrrWjMMQZ+k2n2s6D6y
hKusRZHIUHRlT1TFipMc5Vh0Elm4JLjukTjTT8x8+Hj2IMQgIRgW/B+M0TU2hZJK3Dp+X923U45q
qq0vDo4nZTtQWJir+rtUrPWPGZdRqWYjyBPvEt5TiP6XC9BRF8yA/VfXSV00b2MGtN1GqgyAe2V/
qew29hagru62z2vHoJflmUwPdF6t0769OZ2D4CNNaaO50XZK7fa5CLF2LpNSic9rOtb98uIDhc1j
gyXtJ2NNOUYtj0y5s2vaMTrhm7j9iQF+y1pkUIv0TS65Y4UI2KLMSYV9X90MepBVk7x0+y2jWPxd
9z9EHgq9vtgkHUiFh+POlQg2+ycVIyjCtR6XLQtWtKEHiY/kKvvhS0KMmlDR5ETrLBM1FxYD6qoc
Fgad1HhDPanzC3XK++Wuk/5GodMjQea7nn0dgiNplj7Q5IFbijd+8vlMMpiPFPmNz04vy3AxT2hZ
2mBO/wAJwAFH0c5oEbUJ4RBzUpqcGOXgw/+JRxFv0BlxzF2npAFqQH7J/BInkTAJDC2wWl3nPlOD
697QLE9cfSvI4Z45tG4flS1z8r/wSdT1d0w1cnnYhbv/OeGpADti/ExaDFZ5nsHov03tj6TMcg+m
2phSzXHWiu6SU8TH9V63JnahLmWIeX2SvEX+W8ay0An5uFRIBWQHd9Tk8DQphP7dB3LvnFw4Wm2M
ELz1nhCm2FNpmwBTPGG7HTnkXL4+/6zohbmSOssbMNGh2tXshPRtV9bUMC2Gvu2PUMOTMTujklCA
avk07vVaP3rWSM093YgYCO5iQWaCvC0NN+QwrOfRwTGhcUvp8zY+k+yOQ5OY4Dya6B6P4IsJxw12
FSTF1cb3afhqmH3xwBO/3rcrQDYubM1Bp8E+2ANI6N4QRRfBJzeQcu7o4L6i1Drj3G3o2PLt+O1a
UvB5Hs4d84GPMMLbeysNl3rscqx2wECiNwy33047PVztwaLMKhZWXWed+WtKzGYA4vCY4YJK/XlU
uQXl9laoga2B/G5jqHAovlMb4eZhbUuH4KQDvhtUA8+4uYTF7q6+hTY27T+Y+C+u5D1/RCzgEcdB
ZNwIEF2BAITVPpvhB4NnL0CNDU5Tp+a3WUJxt5pAHXkami8DD39n/T81D+7NVQKXldjQb8zJG7z5
og3kXtuat9Lcx0n+smvCC3fS1mJMfm9lDKoicNcniN2kKLWyg+RhNd2USnOptC6NiYfOfzQyR6NZ
dw+nV0J+iaWQv3Zux9L4OCshahgx00+P1rdAFmzGQPfX4sjVIeZ1lqOAax0ZUx3P2fTrkxhZzms8
OmOesyBSmI0Tr1vMsVW18/DmDHvz0gFRL0n/ev8lOLE7ARAXSpOCQ1lSXByM6xMlPqHM/hJ7lH6k
/Iygi+CMlDkc0FOFnJbSMu7tdxHknpaDQgIywHF3+pbD3FrlxzI78w/9BTawdvCC3m1JvIAMoX3A
V0QbXEnYFFVmobA8yagbLVVHJ7dDkaNidZc4wMdheqR9c6g0fnyLqLPcdF4JEjDh+s1hNCKzd8lr
x9KHSMa/baj80cEbP+mp4eBlm5ehicXN96bTpNG7I3UJrUGSXWfiSjtfgUb9hC3VJSmcwg51b2lL
WrpEo5rYWYL0mQCVBEZs7s2idAW9dDeQNiIyb0FqeSorcgnVC9gA6SaLtULyWbkwT6yAd2hndkU/
DNyj8+xLEzvZ3XMRLZpbovMp2mCbvn1ClNgYtRbyruG2X0fVwd9wfaz9AQ3IOKeQmG7FUDaUaCbg
FbDng+caq/0e1zawEejHwL6Chu7+vgscspcW+5LfrFaUGhJDDnwjPwdxX/xXOH1sz0WS3x6ft1g0
KpRmHeZYZXcIUqjO/1/nv56oP5/H7yOH3zVZ2dAt6KAHLnbUy329UjZgq65XU3YsgelRISeIiEUP
yER+NvQXkLnB6qaPzC/B4fDxVnwVXmaiPeGDgR2NqEPrLnTPmnV2UBlqRZORdmm50ajnD2m/ZA1f
2hL2TgM5qFG6iX1A5ugDojM86vOcrxSce2DS4KUm5g7UkDhGmbSWDDVKJ5jhwCwOARBAcIEwVIbA
1Hny50BNyucu4Fkpeu6vRbp6LxcsehGizvPDrA2w/vFVcM32IxayguglA6BvhQzvts37vJLxU6xj
K84F6LNEiMQYjTttI4i5yNrqhT9Ixpe2eOW2CQEnbma30YQ1OMBROmH6ezDWAqSIOIavPMWHhNUC
S1ogqP+TxflXTe3QcSw3CeGwCIvVEyrkwlq0zyn+3kXtr8U07a65wXZ5T3661dcqyl2ukqzOgElL
sG0rdq6f9kC1Jt2aHRmZ1NLU2E77YWYhN1vYYmzeIauEm7LVB1MmceYsWeAEa8AacQ8VIDu3MIC6
wAEyJjBIrJ6EYrqH7sJSzt2LqYUkQiJrrmTSv5h2cxZqRrRxLCjpFbOq/Wd7Eo8jjHqHYXoY2AVa
ReZ64XfUHv2Cq8d0XZHWKIFHiymM4+c8z3LC6sSqU8pUo2jhEgVCHTHlTof2BEsdh83+OK0s7PaE
56M+RM2a84Aylcof6tvjK+OqNCiztcq8GnK75qJXznFlqPHQKqjlQSADrGszpDGWRm29mZk8dWMJ
N2DFKcADODUDJCiSGbv5ZkoSOCEGDT3DMSk6GsaxNnr1N3dbQ9l258VOUcd9qZtS90uZjGB9BoF4
g2pPn9zV6V4atKJ7J0GdiTiBrVMoClS+AqePaU//XkTyw2urBxVK1o2Hx1gs2qXzm9unmuJh1iUq
opJqeVTUkbHN4RQiQQK9S/NSi8uC52BnAljqzWfz9XxyFV9KIJTPcaz6O1kbsz1pq7kBXBbVqSop
ns1ee+nripnu2GkuEZe0ypEI/jPzMIqPT/NdKJS5ky9Hhdgl7CI/3/wNpjXC5fN8+ZLesfThqUcA
9YGElOCYJIsKMfSGY42RAVKF1A6WCgMUzWFL0BZKDGcSn3NZBxWwB67J2Bbe31PDkIxUziYfIE60
fZSta9Lv15TCCkgD5hJAXzxFLKsseTm8kh80ChGFwewZyJuNaPPYY6rqqnwAgE3nlttqrBcCD/Cc
bngOZ7Db4OwcorJila45pLoJmOPWZmoqdo9TH4FyFKgSKQsky+FWCQBHWap5Siv3jXjTJdncx8Wi
TFWf9qzFyU0CA8rSW/2AbRZxhZz00ACx/eNzvRHbtBzoergqx3hwcgqaWeukEaOnQuVDe1nqj2Ne
LEtO0iFWmyfGVXAwjw3tlAxwMeHBn6YlXazELyGObw1vMvrQAemp0gJGOdBONomM6sFMK1RxhJ7y
8DkqnHviE5BmdreaRza5Ty+LER5asq06Y9MqyhOyiC/X4Zfjo9MbhDxAVtlQGxwK/mtTc1Abg5Qo
/g/bHc92+/SKMzMIwATFes9lxXlybO6iRus/SA1xj4DrgnHoO3/5zXz963W5MVU2GG+li6I/OID+
/MqLUrbXWhB0MoB7VDYpWTvRhcE5dcQ98yE8wDKyz7ou5Q08CNHQI3ShTKKJ32qA16yMiYTgfTzz
sYhIgoQ+SbwZmmeKsfYte8+mbGhRnntJiEiasnbVc2Fu2v7WVcZSqB2+rQXjIZ3ufFcXez5Nc2O+
achuYqokNMPd3KHMhQh0M939f2YLu81+YXc7E+3hf9NKwdMI7YbxbYPSqKOu3ePF91OGHE9YJiJA
HT4o1pZ0ANvexlIOG1G8ft7/by1Yn8GUrHxxQ2WqgtrNi4nMgMJ0e/tHM2xsFpARZnu6xs8J3y8m
X4nxjdlHe7G+SEDFuD0KKi6Ci5O+h0hEKAo2Negqmdfeszup4yj3SJn5XkXU7Tt1zXq4Sp/9viAr
JU2IYaGQdh3IjBVn0Ax+NXR0msM90A7xxcpBxk6wwXpWEm6XKdILF4jnW+Ojcz7kYAxmXHJAupPR
tEiTIbWVOMPZuX3ByTLY3pkOW0shv4QnuDnqQ1d4vQfpH3GJIpNg4qLwW+8H4MSNJatkryl02YfN
R7WhdlOARZkTnDqrbDINi0atE5Jij+cBjgaylZ5JcckE2YKBQ8b8gRmDPos/pCXvIuYVNJuoAlUL
d5J8ofWFFZ4bSBY6vJu7qzQrtkRBW4OZy0/JSAFiP5CS6HXM3G/ARiJ2aMQ7UB/6r3Prq/SgbWZK
lLTuxFTikou401oQfk1UfxhC59YU4IUF2cJjdc/Q3uNR3+WlagfXcs2HEQ17hwO1ANxcX9J11OzX
d2QO5lg7TWqGa/2cdaQZvmkQ+2UDoJDGsRWZF7zPEyzBaYvkktYgJtRya/LwaFT43m2rI38QYUwh
scdeboPEsObPbpHJCuC2p+NRcjz0VDAHq8SPk0IyL0uBPg/qdplg22Ouy5oLgAUZX3j8H81qNhAz
T0u3EqTKMCYRd+pVYUqex0w3SrhyfYvgmVXBthb+FIFXtZj741AK/kASupAhwWXFBIOULj9ErUPK
EbqLtJOQLrrzR9ppZ8i/9x3C9G8oPPwU65y2ckDLH2DZv2u0Pk6eXydazj8JXiSwYM1e+WbKF6Aj
/QQ4ycpphVOiTM+8GxNjsLalDhJ1/ofOmLaQLTFpzwuDes+5pge9ZShQdyvrkb4oHr1hFtKqMMIV
GJJr8qyfdfE0npU/q359GYnSxGNIUjwDbgQjfKNvNg9ml9Dc5lif9Ie5zMqC83zX8uqLh8EPnhRd
dK9i0nyrO0TLIXG3SNRbHlEWGwwTx6sfF59r677aAvPKtuMgU4cW14FqED0Kyce1kh3wrBOB+yfA
YWKBB7IdAZ5EdSibqHoH/ngKBjp8pjJEJKMXEbAWCe0G9jOVQdsbhv7z0i0YyMrJ8rrM0QaHrk2v
Ep/0qdrcy0qwTF48iVxKAlgnWfTexpX4vSfDiANAJrsx7VoKTWtmSRIBIFWiaK64uLry83ogPaOu
/T9ku+nTwnIQ+RlrzSc1lXXnm6Apfk5ZEFhGnzrs1+DFcklU1nivyVatfHG5ihp8bmD1ifWhIky2
uFB/IPj6V+3ANn2Ae8WYjkjmEeYVkfYRmS1Ru95CLkzo8FJdfVn/iTiXa9tpd+/zuCGizpr33/r2
kSi+ICRuhWJLnK1YozIfHm/kVL47QrQXc9WZtEj6p8d9ufWNXQY8L9T3xXH9yi0ZBkQepaiVLoqA
P18PMXjPudlWifTUuXzf8GPZwbpciry8oYIa+hSFfuibA375hiNz2NZFt9uiw8tM4ctG1ToptddY
HPhjhJ6C7p+sIoi1pQJo3T3J8vUI6pIDE4rky45PHn1ksq3osHj20lw3qFMQZDUGiAAhL3cgvfAJ
c1RdnGCCHqo+2NJq5VU+YkiWpKyVQAVFyUaTJowJZ4cnN4giWK4o++fUmBNDRyaXH1MjqeTBHVZp
pnUmQLGMwZzTAVaiPHo2Nb9y+yp1AULq+BdiXr+quRN1caf6V+d2sVJn3HT1452wvkCIxYFSj8eL
d1P3DeRlBs2XvLLm46eUdwTcEbaH0Lz//4vEmwWQfcguRXXeJVJQ2NhR4v07xnM+TLxxV1roeuMk
tiIkHu9jC9D3hXu3FbAfUBUMmtK8qIIzdGs0URwaNUa/73jUhFBM0MFKJ2Tx4ITJhEBYmrkTVb4U
ruD6nMZ8zKIywQHMnhCN/u+tZKIFG3lzv7/PtyZ1kFapZbV/JIzQUtJ0oUkCDH4DW/XNcFGWNfYm
4nzV5wDCFjdd5Vy0lDnTsqDND7rDOEWmIE8+7QtFnA3kRiOI6bO5ruYepT7IAqTsQ1GAouQOzlw+
ecHtoIQaXw2bzKEVmw2AsFAqFcKm9LHmtKvA/FI1QXDF5/vFhsHwAbztUWH6t3nYcWsg8hGlChfV
IWvLw+k2haXfL23lGouX1nlX7VmM27/Mdd5qhZo03fTPFbMl3uW5I+EHCIVXw8ZzHwjhiYhP1GZq
HyIykP2ytWGxPE1GH0fsUQcvrbJTsqiBvWmIyT6TKsP+fYTQuEuueDGMNEKGPfR1z+cUcACw6MrM
gkddAxiU+U97QnxP/+WLsG4tiekLCKmB0fwHBM60kgC8D1UKCT3Yf000r99hccYlxISyfVP4XkKO
DmU1KmclRqjQGjfOb5FaOTGgwSwxbPew8B/kDJ6hYcaADUVws/PR83B+uvSA/i3Nd/Sd+EGlGqUy
8wztqSy+BEyuaGlNgBXb3WK+oRYwpjcLZT2p0ToAr3ii/kdTZCJW6a7xWSkqsLWzB/5o/YnuxniE
eKwZHNR7QTo8Lkkt+7TEXDT2zXISCn8rBZ2pf62+u7Aq6siwZWNy7gdfTT8wB7UzIb+BZwPBfdnx
oRWRs+x4Wd+ncjdQ1CnO9S28LmJzTcTX55SCj+XDpTF1GLCoE145TwezcFvyTU1PNtv4LCiPiQ7h
y6iOTKruNjU/IZgz5vQrsFLmx6LO74U7sgcPr62FnV5TinMv1nLtPEkB7LVRngXxQjK5C6rU52PE
cSlThyiVdjMTadsTYPm6PPRa/7wDmqtENjBzRHi0woP48w3ltqlSCWxKBcVZGGbRYPxxge3pPcyU
aC9K8iZLHFzjC3cf88AFJvUJLO3wjSJfDhAzRIPL3FnnHqPjSQbGvTHtSpymFHO8E4F6C9vziEPz
PtxWBLf9AGVGHptvCcQRCoY4L1NemV61dR1WtT/NxXLP1ZVr5UqhB0RJKQiemPLQvlSNYWhVLOHI
OftMUFGfJNx0Cq/bNWbXvb7CdET3tfFvYSZ0L63DIXHHetRlmRS9DrK0SwXODyfPOaAdhHfy0tlc
+ephx5YlezBW157wydngMd6sh+1LyVqosvJquGBICOSS89I+2b/G4SAXueLmgAcGjzCxPFD3G9el
oYzT/m0ydZgy74aMOZbJqqpbLlvHSzU1LoNxaF92br1OSFNyXP5ZYk56T8M1eXr6PyaI6EG1fSJl
WEvXy50k6yoiPDLXOmgD9pXvyryL/2pY/zj2jsgWsqZa6tItthfm+xBAhqKZhQBaBv+m8quZUhlM
qXP4ik9jHO8oUjGGasMqz3mUWn4ZIXefKVYz4YX3k6BfZ/Fy3C4su99RlUthv3AdaO+6I9MvHWVn
TeNHbcZWZ8NkHG29/ZyG+bkMJPEnM5IE9CeBusdtMFHYfsI1FSmVn5rfgu6FsWBnSH6N0Bqo53VS
sMlb2zRgHe9FS1f+35v39tjyStBqDTQ82a5JDznV+aruOoZbUHhZmtgOd6Qv7rSWBAVujSRSaoTD
1CWe3ddU+mIX9rkXM3mELuSKlsXYc/1v6Q0WjkCCA5H9+9wBxXgY7hMPQvxGbjlyaIqKCb5ch57f
wmHMefCyW4+DGnlx2W4hRzsM/yJYauxg7Ku/iY/hOlKwUGqP9rWW7FR96HUlmU+UIdEkt6UDecYk
2zTO85U17BmSQH8igx0RgA/LpMmnzSs2Yn2fTs/P4Vq/gxhB95utDpNZdxoFZDNwtgZd6on0ISFb
QxVcqgE0jqu72lWf7VxGu1kWoFgY2fszXis+8E5KCSVCODVxn1Y7SpQl6Cu0Ez+cF/CLwx/Arfff
EAql4t8SJbYCxIXTvNbULsxWfL5hQPZ1YQ+gwRAjnrWyGAMiN+52Cgl+XWo0r6B8pTxsvKvMPoFc
T0xXVk5stcR5CVQPXXEMq16fgvdfc384N9oYJ8cMHBPPzusRcH7GbQlBvmVk74WajCfwVZ6Qlu3N
p39yIQvrFVNVlOJn00BiR5nYTTZr9autqzZaA5GG+KODKdIz1XZ4WJoLYJ7fMlZ35khjhkS4QZbv
Fw+AoJyV1qk/OzNRkCoG7dP6dsmLV+qKhArrRak3PUsI1wEL1/NvLZSgRTOr7hECDy6m/lqDc4r5
0aHVWdxlGEt64OwHcQqOKZ27QJy4t7/gkiwSmragXxvvjqk6nZWpt0H83pzTwU6XnfHZnWDOwaEu
oTVXrzn74CbhFOVUog6knbb6qfj04NTThblVNcRR2OmldgZgrexI6ksRa0QSxANTviVqAv/onrO4
xe8b94WLEQif4Kd9gFov9cXv1heHwbb/MsqqI7FByJbtzmj2n0YLG++G+zvCP2WEXIRLh6tlFfCt
Kw/nhpFAXl7UrahL5ZJH6lsYQI0J90Jj4d3+oK6mPdo2G7v6JvZ0e0vgWA+o7yKAbNAhkWuwUbbr
4VR410eAwVr1svgN3EfVlL6aXbl5aQIdphHVDjuJBWnUy6KQjLQelg3dgvq2tk7/ToPRHEcikULZ
SO7/+3T1yVyBpf2yG6hFZt+6i+/dQANOwEX/NiSIB3NKLhR+K2U0C2SddrPUB1qUmGeBKf2iEWJZ
FDVbotBAanZygHd1yu0vdv66FjWbirNjCpGRzdKWsRucrF7j/mNDU/FGLqFR75l0GrD5iBIJdYHN
IWgvbOO7Xx/3TgDTtF4dUVCIRZenqtye5HTwWzgtnueXbYo6r+JBaatpXumvV53uO5V0gXpudc6y
Gqrzmo7DRNpHIltKcqi6alHNwQbeaSAzHA+8Ss6pHXCJfeNrqARP0cjsCcrVwjSiSQHJYrkNV1H/
Do7R+LCwKCZoqm7ukt51sqkrHP9qsnd+TS+4iJLJXSLVlIB+zSse+/U/MdywD50so9c+jSz9z6gQ
IRX20vXrsXojoe1idBSC6MmXfXhmcW9rm72vZyqAsRdUBdfs3t59k9Ea+LVrckt8PMAyVM7yZEFB
SR2G7YK4j6aXFzCEWlqMgt7cY/AuXAzDaUduFjwtiItgPchhM60jGr2NU7q2FBB8hNepHoiz2fIa
rii+zDHOF8stbAvOVI/9rywTjaQR8um41bVHqcQNq9tYSkPh4J6l2iKGDA8sqqplwGGnGBmjqxvq
gVrD2kMhq/3jC8LJCUZB/1uelo8nSTdUO8+0qKjLB6POzDvyZwLWdHVFhli4THZ+DtSBnf7nQF6o
AzfbStGXqvgswPY0+UxvSxniU7CxX+o4OqkH+Re7ZYWSzG7KezJ5JUV+HwbFlkmQdBMLQdpBPMH1
PIE+9xQcS0Dtqlg1lO52PxhSUtkgvJlmb/7NCUeiRkBXsYT/LGkMbjJ0URRbT8oSlTSx4svwGtMp
RYhjj0l9krC0fWAffVaVr/JiqWIRHc8L1ZCLqJcpRb/H2ViUFCA4jNtaUuGk4Sh4/9TDCZ8cuG4h
dbF/EWvmOpKKtJ1c1/WFyAVCcyHm/YNEx9Bw64i3Z1ZJBFQ9glsHPimIcru1/DXSwaf37N5+a1rp
alz8b9avoiUh2vtncKdfD4HjJgve67xqb4GEJSeLaKergwJlyWUURl/vR/wXT0BXYrrv5YGeLa77
oMegtIuL8W6d42Cz68iMdDdGewoUUrASZzPLxaEUNSswXzc9Bfl9EollJJANq7ZMhNQQai9qYTWD
55bzPF16mDnd4lNWn+z8hemY6mRQw7F59L8CI4HwH8a4Kj3EH0ubiE7/9f+iY9thWCV1Wl0IGvK2
OmjwtlqLKe4qhCQqlgwgHLUHRFNpyQvtQyHfyxuS1BH2m4q2Y5BQzUTwxCjSWyKChVDmHcFBAJf7
SfR5x7TVNOgl+iD+sRxBTb1E9LV3WoNH3jeX0ahKjqI1bdD6yOYo3ciwcCv0Ri3AIgQ6xSFQ4pSW
tEzD/mZ8CG9kSCdDvpZp2NYeTM8o3rkynhrT3ShrIT9ujFuhTvN+UWb0hi9b8/736knji4OcNk2I
OSij+shRQZaaOriR9ywdbJiFNDHMwjDJ72jyv8s1yGl7mjwoCnsXrZuNzgEoYaONsJ7322EFhDp5
T/xU5kQkjJzsSEjpf9z0O4kDDgSbIyg4SlATV8pw9F/V0fUDGG1q9GOEhXq0RVlQTck4xfaeYSo2
8g6l42+8Z8grAs3BgYTBtwotMv0jJ5K6nos3f3fdFc9/z6FQlVZaWM4zF2Az8LJZaHq9Aa0M8rJ0
YwZvK2CnK+j1UVYG3U7vHsfzT9DTdygTwpZFJI+TiykN4fETu/XTinPnzPAZJEWT8C5ne88UkM2Z
0iH/Mp1J4AwcJbdf4Eg0gSpZXFe+8ZkSnFHKLu82XwLRglO9Zj3941ADJP2OpRbDa7RGBJupAADU
4/gLgVtl7Druqtzzlks3e7s+b7gQMIl89jckJTpCUNe6QVepPg+8yDoRP94xX/XEF0SBTOFh7zSY
Mfl82veZaZHtlEAUyQc37To6bozPdv4ezxVr9f47PAjzmZYp5ZJEUBcvzSU1C7kR9FzoQ2YXrQ0X
bI4isZK6kWk7DgvyhHhHhHrli0JxLMk2ZjzLZ/jbhhEEyy1Ci2FPGGl7LBoCRKXXYw21ZWGtcO/U
Q9wLtFxGtCWK1sK9ZR4HcbDRDHFnBbiolkYzBKbdF1mp9UDM+XQEq9JAo4k6Xy91XtyAyke/uv5j
D7NVWpNaTixJaADa1chb73e60xI2LP5KEXZVBJvyLGXo0peIR/NMazqUNI3+Yp03h6d4IdHlDwds
nk33Eebcf/NJ5IN6NAQgudp6TMKqtDwWVYGMjM8BvD4fiPipyHRTp1Uvb0N54jKCR9hW15jKApls
A3/h8tAMT+ZeJRnjc9lJhxvsc+XL+4ARnjugV+7OTEA0yY9A3udI5oYeIpCUDHjY9Ri7a+V9i9c5
rsHVHnvK/vMesEJPTIXpWz4FxO0sBShpWiHTD8IPI2oNBB7CHwRWDBDpgKff9UGl3Uq9a67LHtRg
blCLOeQF4lfCZM+o+iso+gmxbv5AMBNL4OYLWvxx29jWdwQah//K+HJ6Q8bB7183guMKXW+8E/pN
M0zbNpvt7Qf/O54nIsF1jitkULqKPY9Dkn4ZFkyCPmMHg3wmWmglaZt88kbJIDea8mJp+5KzyqXr
kec4Z6h1fgQO9WUWS8QV9lZHVefcng272AfWhSugu7clKzo5mn9Qtu04n5SDtSQqi6GcF88qdw6Z
pwXZnOOtcfz0b6VWv/kEfrTNYZp+X1+EAntk4KCD4Ot5Smf3CW+LmQz0H79CnNPl6YLnTkGkpeXm
DFCNk9uuTD7v/3x4WIKjhrLMJq69Pi70TrpbFYaN4YXaMB4/fQyCC0i6JZqc/2wQgvlL+/WyDx13
hxydifjIxF7P+dvEpnzeLp0U+tc59f0BSltIULWKp2EFvwZ0V6vsmMlQ4pWYPri6ZGK0cCxALmuD
e8tDhqZHA39tdmleNom3byzc3vBZ+U4XX40y1AWxp2jmDQG5FevrBeNJ07Czoz5sdZ+XzxrCMkpb
2w8h5PksdTGjy1fMoEN0t9JlkOvvEzSpHQ2cQla6Hf1NTvnp8t5qlUISoDu1CgtXQnRhme14EUyr
M4ifZ2o2dAUE37ophl/FlONVenyFvD764EIadQgP/lyDvlbt5+FVcQF9mpJ/p9D99h1Kbr6ailK0
eDIslS7LgMctGpn7mONSV/aQgWGK3B8kZu8JuxGHbtOCUHHmvWSMgaqmSwtsz0JgiDxUBNf1s91I
F02QxL8ETl4I3hzDzzDkSL73DMxTREG5gblpwWSMJbB4MfJlZwGqEU2sppcty2Hxc8jcNrWqlefw
e6grCNfUmdrySTvKZo4nPvXM3LczHErSyvw1Y1cCHCjUapQ/45/yyZb758DZkE17ARYpKkkpfroa
Jyn/h5vg3ZnwlAwylP6Ov9RqcxJbLQ7q7/TkSaAyruv05S9+cndj3gdBKoT5tPL8B/1lT6+laGeG
VhroiTGqqayFx5CEelLioeffenGP4Gf9VZb2UgeGCeM9TjVERSVQEs+e51DB3wP2KYrjGrRLF9Fv
11T4Vf9HBM9ye4DBcqCP4u1dfpfNMrDzxh0J6KtPlaz9Cs/PDG9VZ/4kwGD6okJaF0mHhWHvvb71
DSfX8KwKziPTes9/dxWMNuCjfVQqPLPl4H/GYlrZ1RQtPYhSxNSNnPu/CvgfijrYe7MK57AIzJDX
OyvunrmTxd/R8nA4R7DJ56IiKsxlrWslLU+wQkyNwWOh/zb5Qn+PMHCq+7ZQkd80MCb/Y3gbSDOH
ujNP19lhvuk6WPOG6PbKmsfManzRxzXO8/QqTryaFpIKkO6ukVdtGYiKBx8xa5KCTm79y3QYmICh
wsDAyVPv9UVK2xU19UGRse6+//RyxmxbvNS/4gYdKyrpICx61m3S6cWtamMF3Q92E4nxpawYdaf1
PrT8APY2wCfQ9Yzoz/jdOIX5d7HreNGLdgtNIhhVi2LPaPO8zo9MGO2Ng2yzvemZsVWKr+sNbQ6E
Zi2HI1kIANh6e9oIyYLngcl5Z2bIb2YnCeZec4qN4hUXFDX2gz3MZsfEPfua+vskcBl9B9jcWGS5
sa3Z+0KmcNHBSBC+/jLlVWfxynCCMniIrXKzXIAiWy0GS5oVILfOFK1xDJWItO7KbmsgPtwSEWPe
fySz+TDVuCmoZ2vliJtYYbk3q75cWpkzzqKvN4eWicraN9aIrIpxQl5xm6q8IRFr+CFsthUSq/5k
FjJx+kKmjWxQJk4fGnSF2lB6fccNyfhgPbuo38HuOKKJmBHcnSI+rYCLHQNkz5B3q3iy15+EdRQm
qZ0CLVCW5yGz2fr7cHL5j3T3tpL2+mIi3orPPczcObQZONb7xbrU74yUMnuxIkuLBHlzs/HKXNd7
UAg2rLFWFZYVgvI/BbnZ12W7vmujcmCrmWQi8tmUWDItUCb94O4MB/plIE1ReY+REqufio1RpxQu
EWl7G3BYPheJ0nLBlr1yohZkDG8+eBQ4DvNFJz8uaas/llVO/hWbrU2RBqzX5H/kCRDBvFZvp04S
9k1e064jqTP+h1i7vUCaKARSgFQnkFgTI3v1riC0d7R82dbe2ftqKS1jEAg4eo23Oo5UBKPzRnxS
x49fqULLYVpExjqqNnoMlYgLc7FXZBfqKfOVMteSFGNHFnb159l20x2U/kjHC4tYfDvGGFH/C4D8
raPveqLn0HMlot2PB5dpEHItw+MyOBWAx++AwSTELjfI/WDE/Ohlzpw80AoLf2mVvzDD2hoWf6CG
FiUDKisvyCtacMMcXBcpaBYV0OXKIIrX1uWeTPQ8eyrrjzUPbaVUJhHiwarx/Y3r8K/W14bjVSGc
vYCyNLUg+X/Iiu5FdMb3C7lM828ox137hFOdOu0As6KZlMMwohVRsYaWOYMplHKmzGmdqXAlhUDb
5BcQSsV7pFecayzdfKVYC2N16eCcOwM0uJm7cKwGYaIlcdf+GHSKWh4GDGyvk/FHtQd46yoMX6hT
vzLB2h3j8weWoRvqWV+Z5Ps3SlQCvO5U8HAzuyzm3vrSXvX2nH1KNeYbXNL9z3zFhckZyCdySI0R
Gh4im/UUfhjPgC2EH7ErGqPKT9lm+ohvPK8SZez0kS5o7SA0WslBv/1XgNuEllSKTQxOQNEcVZrj
9jfy2mp3yEuslP0FVyToNJQK3Hd3citiodeJOxkf/Bso2CC8ALvOejF7O0q9YbSPEmSIRDDYhFvx
Yb/kELVU0Xj2O2X4IacdCviav6SXAqUJlcArwPgo7Ntq1JETSNziFNihqyDSgb1DW5BIVx1g4CzR
sRkU89lu3dfHTRpWxA///nPZdhn2ry0sDjzoCCecdhKxIA2FTUdYwQhSeElZC9ROxNZuMr9HnLtI
MO/17m66vEj7/FyKgZwxn/NHfwWJqpN1svWMJh2VYey4I8LfYVVeLIBKKxy7W8mv2TK835LsyzG7
0sifFWEV96FfIsaXLGm5Lufv2KqsVIILzCSsACqbcUYkoFUJc5SJpBLVBX34ZXSWHMAyYZw6Ly7X
JIiXaZ3aDIGwaGDinGGCV5M+lHPJlvd1hSkPblRF+r5WYI43nXzhafKaapl4nxorWrJBWZT4vtnK
pC9S6+CRmHpuwtJGB8qHF66nHlQHmLHEKBI8f5e+uyTHSBlC/AjBTFlGG/hOXnABh+Bl2BonShGf
N8Bod9gjlV7drHSdCHLUuZ+aFO3TW554N6SGfjWTVhYRgUHd9CsHoIelrn+3K+GozXWE7MM4Ad0O
N3ga+DZvlZlxTCXvSrxj+i+grFZzk/FtPziF2aOJPFVnlGy1O0ZKo947z28P+GZEQ3C13Nd+xma8
6jv80zySEJ0kzCkfMBwRdbfZRiWb5GMTAOk42OAvaj0Y7+Bbv6fu3m9K8zFw4hhtRjIRDZpzz96p
fMSBgT0AH2NAANNxVuoQ7HH+2zUm+ZKyEnKVUgAgzUW2KM18hrhCs71tSEDwGjzvdZu2sfuzzSgX
gJzWTzCFuYpzOj65xeuBIOD6MyqFhFIghy5Hv+cToCqayWqPANuCr5G7uoImIVQzTu+bfNluR0Jt
D+ndmBaOhhZNDVTB4djoWhTHf1lT/ndx3budCg0cbE4nUn8wsRz82TBeUM2p+hrTtu6845ZavF3p
JixkAJbS7997SrFa4xBFYXe/ytkbdhfkfAlISFebjw5adgGc8OhpsE1Uydj3zs65r8DMODpdW+/q
f6xusSgcqFh1d37puVgdOG8HEH693DvDddXUdbJ8DJHPQ+Gt1+GP38QHP9+20X23SvjqJKBlKmfg
IPyt7rcYUwpElwmlXDS3GG3hKWjnm8zvB2P8gqNaS6uQHK6mzb8oZ4DY7o+h326hY3O+eyFwyxAA
LOIa+02GQUnd9fJ3zvRPJhMHnV9ld/n8Ju6zXjBof8nxW7BmAcqaOpg7IYJbjilOSqJXltGS1+sr
9RBugAzTAf1RIubjK5boLaJ0IRhGrBvT5RaMEf2HIM8p0M/cGfTd6DA+LVfo/1qJ8qQMzrS7KfvE
6ItUBe4Jgt+zthIPSCPcPmp6GBr7BxyLbSLkS6lM+n6kGGjU6PoodEQYz7eF6lY6eeMnKk/wRVnc
By06PWQQIzjmNBoI5GDi2KMZhWv201luQW1JlzMC7YBDlXwQxAe9oW0/J4VC6dOts+0+Zp2+R9Ly
UweAoQlh93m8x57Eftkn59VEmttaj/owMHkPltRxp7FoNtz3GrpbsPXQ1fZE+5Q9PNRlkKXNhsCM
yOxsPjNGN4DFU0KOTT6yHtjlD0jx0VZ5ERM/iCWrVhQFEMomWkWsFTM0P1ZzFeIt0b7i7AKU7taD
kWJzSyaNkyUjZQf6yV3LWG2Pzqc8TXzpXdgYdN8EMzLt8rq8qDQnRZR3+NFPEG43p5XNZ7SPcUtc
edkOiyos8B6ElJIcYle4QPq6L2puRqQb8EJaaUeTKO5UIrMaWzSl8EhTTJ18ZTYWDUKz+WzJbuJh
G6oq3AKNpt+Hxptpht+4ekaPabo7OPC1GvKmCZEOJfiJo01MmdsnIYS2RW7jnB+2MJ5C2kXlauZr
IA3mx3QysvuIavHxGaCrVD5k4wOIl/dt4Z+51JKvmv5kYTu0JTYEtI8B5u7dVfJ7cMIa38wD+vQB
ThrQup+c0AiNFYTZUpgXmLs58PR8g8rKhOg6ESwpwVFQWhLxEXsOVPYUtZoZOzEZZ6vlqnWSBYDP
NoD1FrGKWS+datIgpGEmpiDMH72j1pbNqKG8Bn3KclDf/dHZjb/6iSeuIJECcq043HXqEg9aR8j0
QRkRjVTxH3c//dSFoTZ8F7HSFCN0guXiTAZ0eS71vlncGa39weQi1ZfCfhjvxdXXX+DmmLYtlMDV
CnUbdTckGUdRKY8SgRSyxf9CH4+uTov2wFAvC7NNihhb2FVhTyUurSBkjeTJTTymP0InRYxehisb
J0DLUfwdONGRpaFH1x2/gPuc0laffSePQAGw3aGPl6eW4baa6dJsL1iuz9Li1PUQFEJMN4hwaLTd
ESG5s/NB4d0GJwozej0NrRWl6AucU/ryeQizWSO3wgkGbJevpsAywhrbR9oVf0f2f70OxV7gkmG7
8F2UWbFyoLDk6qP5MbS2aXRPp5BB3pT9w5L9P/fc1ZL4hEwRbPJsVKpEkpvOOzJwCn6Ki/g6W2n/
1ZmJ3KD0nGBJDShm6/DArKrScTdtVunYJwqF9xXeE/dXC8g6OPbcfe8du1oNzq6vdlAVIGAn3zJ8
3luB6ja3ZvTMLPyKLsqyvUZ6Nd+RP8p37EwHLdvIU04UD/JIzzgOVf9wxUZOyk/eHcFW0KVh+qcM
HIsMeIAnPi+JD0AWRH1yu1mRfOBCXM5f/CE9IhZOoyXPiQxXLm9B1k+e12klFo7wHr7qml2sMTNR
QF3qB6FkK8hUFAO+fhWafD4Esfa57ebtrJcacNk1WZv6Kd+Q/TTyKTlEynnYjsXnLzS2V8su4Yo0
x96XPW4X3eTKPHtkjGrB00RHVY/RcNh/zOYRiMyPOs0OriiMh6BF0rTo8JUBROmfyY6/GC+q0IVg
PTgYtHNV2iotvb6/TEEkZAWp21BqJvAEnkPB/BZ9g5Fgz9pOvn/C51Fs1bxTG1kkQTqJRrGwB2+4
FIRZwNdHDsIV3R0BAKkzMuuqF/+v5jlyAU1Zi5Q6MFHw8Kz+vIACgZiS8JY2Ma/xPNosRLzFgYrE
fYPgNNPsDZkHo0MeQ81ODKRIkKDPrklNz+MP9unL6g6Fpb+cccc1Yv9unsjsqSa1eKMCMYv4pzt3
D3PbOwKNXBtin3nwrOXYEPJiYqQq1beDw2y+CQNRJOZ3X1cvwNR/t1X5XLdImpEfLubEucGtnszP
WAFVGZeFy8R+Sf6dzKOfKu5wXPkFeORoITjDT9o/C9eN9H+MwO5wMjBS3QkOVL6Yee70MTKaONEg
3tu4m0sCYJ8Q8QqtNip/3euxSb5/ahFAcCf3cW5m1SDKqsSupc2IR2h6LAvquSx+o7ggaxdrvrQR
H07Jds1tcJ7jY+22i9aDYlon0cCwiWTp/opdKz/gmsrAvGzm/ZhHHdsp5YuXRJo0Av5wJftf164Y
nQ8z5+v+Wi5DOjzkq99fQup6YicvevRKdAALOgCASw2vIsU6Q9FoqrgdtKPYIwVHzpovFGIdRe3a
yFxfNtXxCmIHXrYzQ3kkqLCObE54GWhd4VQFEFLhvvjoeGHY++BxoezsT5E4UXcOtYkZZ+W8rxis
t/MSoouL7VTJgAsFZOAWiSwxw06c91eQRfbeZtKkWIEl3jtM+H1FuNfdvt0KJlQsdsJnH69kP2G8
sWSdOhzOrVUXAJDpwFCZhC8P+dPqbcXqdFGqCiAvyQMIynKfUKINixAyzBas4QLmAlJRnrYJNWEw
ccPu9qFzf7tlYbq12KQboQMiy5ugL1hQVE7qUXYY+bWgIcOyQAmP4cCgQc+c5bM43n1pX9POPIPZ
LlSJ3xzM8QvoBQMNbyqMRUE4mxqYHR243vVmdVnn/ng4b1JH1UXIKGI0lbeQ9fUFtYNcsA7Sv/Mn
GdSgLOTRNWHnEUvm0gbDiM6G2m+UoARgWyAV/H/ysYpJr7GNDh+9KwGSr7I2Dj5JYpQ2F+IG3M9V
wTRKFJ/wNiwD9N8u6mB/uJt2TcTCdrlgSxhe7Q/tabkNd82Kvyml76oerMgzLMB+9vp5GZmR0DEx
h55mLI1j18foHu27fnNXXsl66H5VjNRZuD+xv82/EVztrFTaRzsofYq7DqayheWIQWWm6Cvd+bCq
rfi9LdBaP3THW17hdzOYjXoQvbtFAhxmusMRjUkARTuL2YWcwuy++sjhC4zUB6WB5wU4us6KF/d1
V6+M7ibr/rINVY3UwFgqhPZjY1rZf81svB+aiQCGEyx1D9qNN3BzVhZJPwfOr9RnBU1uCK8mNP14
FwmlcZj3CAAkL9ZwIsJ/YtlJxU18kCoNWWKO62n/6w/NtpmAuNwGeRYDh1orjw1nmim7ND1NMftQ
BP/uwxg7nyLrPW40alPSDHSB6SpZAm31YRf8pwKGMNNeALtVzrjs6LoNjs6sC3RoZ0PYXuXlWynG
QJG81qCkmp4sBKIO3RriJXn6rNa17aw+qupWRWVd1neUYQspD/FP4M5f4vFFay3NnmrqT1BXrK75
W5Ea6mCoOe1OgYybrDMMwWl/41hFE1npvQimUoKDxOr8wSv1MweGYReSHrXt3poEIs5zjeumCBEy
zk82lCCxLUiepNURYE1TvufKByL+G5wDFWIxRnxX7t02iudnC9PaZnbqV44TslmakuLQ62vaT8Ok
3nW38iHTSWOX44/Xbl/ZRBAs86ahtJVvgyCfcwjwaj595zgkytV7vnFvv8+jSgo6sQGQSJ8h/cKZ
vnZjYaJD/mC115CTmePfxBgZHVC9TpJPU6hwB1eplqZK1BMLRC7Q5BMfAp03wWLtJ/I5792NB17M
DpEbHgsXo0IymWNIDCi4M30VVGzAF0rzV9SZMmcp7EHWAKcJAeafoHBzEEaT/+FWfs6FC6QLJ2Mg
RWjjWZ7M3qlALs5JjAuGM++WCqo08M/7WYuzi3BSqw2XB+8l2irjCSSYkjVtxeRz1boUdkKMOdSq
+EcRVtnzEhab9j+GM0sooY6YjRyQpbwpoj7BTicRtdumhOl/DPWMGS5HcDlvD2GkGZ2pQnKQNdtl
rX1xIGXS6q8kXeiDjms+U2wE61Wyl7ANZPCiDcgwno/Y3PD//xkESYuFn+iS43dprIE3lOoBXHvO
ujACCuZETX0rwNKIp7oRHhsXGn4nSA42oW0RJHL36mHvu4VreWUQneCzET+3iScFZhqHjqTzdyGq
47Up0KH2vDswSpgdQYEDHCee1sYw5zuyn7oVEEO4JmM915gtTbNqIXDTmEABaLAC20LdXXzLcecV
DHinrm++j1i36WAUwI3cjGspcrrncsFW7h5woZosXcxxmqMM2Ot4PWv4HaH+8p9HsOSHieVm8MYK
F9umAsQYnia1o1tKmYByeqhSOFJC9XDWJ8CN51nRerzXnMIKXI65ZRihCdmIUsOehA95yEClYTD/
8yaQfIm0NQjiFkASvggOSLh+KI36stH+q0dr8QcoFb4u112t1fLVw+LKvZyRXXl9rkOvgzafc4Ga
RiPYIr3rnBk5zht0Z1jo2ofqV0uC8dZDpZjt1J4cO46/oGgqKq4xkL6XFrPjeHvaNc+KsKSEwbSA
2ihxWoBDOs3iAEjWxhEkw/+ldKLp9i2VyNEzYEO3PpwvKq5DYEGDsJIPO3NzEhEBPOkdHXhSr7jl
L1N9gFIvVotd4LrD27bFdP04H4LvQwluckzIoXH+nIoWeFgLBiBBn24u9s85u1VKDr3HMbj6Q5H+
kUUt7k/80xwYE3vG5EupO0j+V/zCQkSbHjfnQGaXgJt/C0WTfVY96zhRWHhBBGfLgVPnFgAydWx7
dLUNDeQ/9aofTdksBqBgp7oQ7NZ7OpuQj5A4bZHRToOTy83aYdCTVlg5grLOR881vl6LqPb7lWxe
1SdD419TCMQ/e37VHcV+kViWOQL6XbLpb52ofzh5lSJTOGFFJMCQiEgNxP0aRrNikpG9Zvoy2ByJ
9tHRkJICtw293b4XH/FEAKrdxKoSuPuFb9h6VN50Vx3ePaa73hGWnYVKBk/SKTq5wHyKrIQtztfR
5IS2Qb98zzxEZA/8wHRyXKDraZkADnloC6lm30/3kzTPzWMeFfiY52z8t1FbUWxtaWQKaFbmZANN
t30M7EpG6jVkckRg98WFyDHZNfl1u7D/vyv6TvioYr4KOz7TWblm7EziNuKy0I4OdYYZt99Ybwek
hkzuwMTVYhhqVKilkvOMBctzShfGwnxr8c1cSMYxq4g2Wqhf38e76pVPRiSeHZYKAbQzTh7hTl7A
tW+fWOQxhytYMiueompOG3qu8EX5bgXe/Pgu/aHnp7WY1IoU4CHGMGdiYMeDxxDIHEq6vJlJ9liY
emnQq83Ci8mCTfFWwAd10Lb7mtXH8tctvOc9xLcLvwyGpjK/GkBAvsKjUV6Qk223QRkfoYYN55EM
ZqeDph10pBlGxY9c3xyQtIVAJ7qpH/P9DgA7hCG5hpyuSOGaepAQN7AeukTHNvLg8QOOVYrQARqo
R3qogDYb/zCW4NuDfYNcjNxuZOK1StXc7THKPpLljyAWeVaabPpBCVeCFfyecZcPC7KC6gv1ZsXu
veChbM96pdv0tP1u6qBk2RMasVWGG75qRQF6ZoVdZQATT/duPPtQPPXDHPTuAqGhydKqrI/MGPa5
H6Hm2/tX2FQuOwvWKf2q6UD3mDNTD7js/HC9ZFijFnF1NmnwCR6eTWQ5xbddo7M4v+qBapakaMKa
RWi9Q24rTXKtGVOgQdQtNzYxoZLl4biFJjjzk1l0mMNxXKE5BbICESVMxX2eRusLlaz94p5Dt8/f
xbhPRX3mOYUh3fwx7BF+DMIA5k+x0EaR13HfbQqohY6nAVAq2MIauBtLSM/cCaf8yupfc7bc8Z0K
niCLJLl0JJryVLIoB11t+WtexR9Huucen9PHwaWjPHQHgW+EksmNUgHHqL5YfF85WO8HyJjI8GH4
xhIcVJKPKDOvZujLnQigNCdv/Co05vcYbuH8uhnzdXAiO1WrUOBTpEhreLVB4h83lWkgIvgwUQ4q
V+80tOiHlrQxvYZ/N2WBdTJigCszx2QOZamVeXc+CCLjhWKrvhLbwlQ+YB5qtxV3GwCXsbO+pChQ
ShvAAm9wxasRa6HCLnYe2eDNRcspCIeRhko/DgwmmJ2L/uCWp0K4r0OeaYZRJhJFX2VrifOAbtmv
vOg9TsQGZeEip5TFQCGjyl4aWDRVsoHM138Ieshs6i+o+KSFwJVcDMsyhK9PCzaQRAc+TUXdhiOP
XJmVr8r1qkk2SJN87Xhy/x9gfNHpVFKxq5/ICB6rkctiIE7OY5I2+jjS5+SuctgPI9+ZRB/bwlgP
7oycdKI56SY/a28rkmn1Y2/gcN3CNlCbrsWSfUHly5lBPZikPv/Z2srV6odFzgZesWZqEP8em7FC
IqWcXc4KmGDkDK5vfkl02a5+dJpLNsVaeczJKrdnqBlreVIyagKFyvXkpJizoaL+81Itrgc0E7nh
wePWwFuK2n+rxmLrM0tMbeW3u2C4rifHMO/T38btbRBcHcjmiq9KPBRN/bwcOwIF7zaENpn2AeMU
hZ0vYP4UK4goz4JnIF1JOuVkIOFakOJxYY9UGtAB2XVRPBdrG7zYFhFGLXNgtB51ZzDoJfRaQNWJ
S4EDDZ5DyxffbdX5zr3xe3XQ+p6PctRGfhKVaVZe7N3n90azrVN9qSvHsUIwaFij3CxQ81CcI6SA
6yNGSYQ/lCWvZG1tuFhxWvFcFJVCXKN7zt6mZ5NDNG3ffyIKe/AjPUdOw2oTGPrs1r5Ao9T9FKip
XLMMim5izKP67Fq5MeVS1+78ff81CoNjdELQON/j13DazcnAqCTKNA8Z7ZcU+5aNZx14vhO9Wawg
CsBTRMfUCTeMPLdkEO0aW6AgzyUellU7zYsEs7m1fkf9KsfsuDkVcW8sSsVsv+i3pKVd0q2aLKzP
X2+fS8pHzLJs6jeU/c0yAUQIOvDYfsLOfi/WYKlFusrIyjoGooWMmfgxt6II0xbJqEJvZxfB4JsT
WDcIetNJrz0eIL+yDvs9LN+WCNE3MiUmEVcovHcu92qOCLsMEdCIwWIKFoopb+roM+QpTfGIOzMU
i9qc2oB/6YxLlwyPBrRyCEpz+EpQ/UrxG/pBh8URQO0pHNpScBH6AImQrroX5qIfn/UXNUOlCS9L
OPdsYHIjkJ0+YHgyoCDazf3AxReUrxwlrSoHx7G6TQ82iWyxydgXqedscyg5wsmb/C/hIGe1q5fs
VF2MEULicYvl3pdD+Sap0whbL6J58ZC2VDJ32db7bb8Ogl80ppSfrlo+WKnhv3GOIXOK0ilAGoW4
C140GDGx7n7k15ruff6b98bl+HcR8jeW6Il7140ahJ/QugJ54JBUYRiZFvgwT28i2j81LquHA8ej
dYynVj1DiGExawzoaRrShkYy6XB1qNprfA8BQVpRiH5eNZz7khPlUD2alLZSdg2bRZWj5CQ0EKlZ
Oq6UwT2pZHyY2S3bPRW6UleirVCtgjzEy0V0/ohjGCxsydTA2ZIkG2/F3ZNvklWX12S39CQyTSzM
+QT5c66IhRp/TEk16OHbOnDXWZy69nBveT+UpwV0h49Gx3xEsUqa3fhxpX7AMZyaPNi4ropMWo9x
fUWunIFjohRcbuRAWWCJnxN5glrCKcXZAzNbEYXgx3x3g1ffrOqD5kZCn25z3E0izkXqdwnA5G6f
FONqjga+uuBbfIwPPBlGKDDfAfUkSSOoj7ca0w2FGBNm7ErRtgxpKRvt9JmOtdlGWm5zXkRvNSEt
m8J8jDN7yB6lFkvwqfdc0FrD61FRWNLb/+agKE4eUxF7F3npUf4js18L7yNcustXYiRLAShph8Xt
sIlJ/rb9dJljl1FD+Fv9qX3r81s9O4TdJbgKZkSZNosuHa00ngLPO3xzcIyaXOElvXyTAclvFjmE
mYvixxoTSCOnFVKiXifBW15dKB6ikHYsAR26to7uNbwFeWCjM28FAzfvi65d4OlRl4XA9gOKhez7
laMG/aKCTiWj64n1NM4qS7Gv1mNFlj9zOaqOljP/O8T03pXh5ZwO/r9NZQNAmngd6hKsUOgIwExE
mHhxf4DyM146yQgi6CUpZWwNn4u2JpL/e/n91amfIOq5BjqAWEfuomQhn2vFYiX3FP+1V7t7htU9
XfqWp9voRsPZfJRKSVe8YkMCJO0y+gOjPbt15g9nFBI8K+wDGWejruIGg3If6jdLYzATUFwBTHAu
hHuCmhA2uF+tY3t7UMFxnbzjWZbYokBsB/2A+aU6aii0porOs54Jdr6Cj8M/pEIu1P+D33eQiqQ0
hRReJAkI6RSo46WzKiCWz6V8rffPKzmVYd66i82DG5QUnHOmkEaQBaEFO1EvGkf5kZXynKC1p3py
RMIKidEzWQTs54Qb+PkAVzzoWhDg97KZEEWTyPZFn0LR6simbas+cnQu4cXA4tVw09NE45CqfiaV
Af6VkSpnOlHgqe67Jk6r1L/sUMDBA+7fxQx2Bv1dqgmHjP1tub4LbvgTbQIBLkrcsEEbozmZSanL
zDdJjtW4y3CsqRyLex8kzm4J8NmSi10CFuGcpG2PGJ9rr3Cg+bPOK9ZdzVYmmu8neXSGE4iNUY8v
tigNppF4jmoj7R+HOn2SY+yk3qDiSnn84z6GJaGTEaUxD2aInku0F7Fo6mkB9ZEa21XLi+/OZqiS
uCnNvH13I9F/X+Fv1bT9M4EUn/VwcWahkqcQ00SXb2jL8W7K2Qm6dnibq1GtvQNPjMvwSQkAhxRj
bdQp17p/kxRZlOlvY7qWwYJmxpx3V27UpiM82HbnO2Z2Bi+TXZlaLUi154V3RUX/EefMpSSzodKE
OGJtrFkS/U4v5Ib9zaGUsMcIXG2nwYVrDipUeIbf9NvJEL9Aeew/5glmuMjGSVPAObcCNFuPK9cL
HiruZbKDzykLFESZVxvmiLYNoutHGfPPRrLUGpx0rK8vV/kVglmZnKSzl/krKxKPKAocOmby1i3n
RiDivB+v68O7j9wIm2K/Gn8urnxOUU30FbEJmw8WkQ1GG2gHrbV1TiTrgDA78q3Sh/GrubghewzY
kGe9C+23hLjoJxROws1b4XDATb3OKUW9yAlT/ytRVIBEN/GDHG0N66tT2v6Q3NIyMS/l+HxI/VSS
mnfjEYXisVIbVyZVG0+e6shc30i+JepZVY/g+DA39cJ6naLAz4+1XtpYreZNU4pUuwXZ3yV6huPW
M7sXKpQADGtvyEzR1U516facXhk22NSRz1rXmB1fALcmIy6VWASYN/fL5azpWyd1a4jdg3tr+0Wu
ntSrQhY6EqfKYIJZfcy14/10GvhGbRNDdfrOLbZiyjda4Rv97lQKVb0ko8UBsCxwxZC/Ni3USnVV
jdL4W7Tnw5bEXgrtWET2fU67+fTsixlo5elT/peK+TDVkzorIJL4Tyb2TSC5l+Hn4WQJcqNyKlSq
as8DtYjrJBi8B7wc9tLV5xL4/DJWXT+tUrEGOIvAuV4ePMsqqfhlZ6ScBPAyUvpK7UAcfpZYhzd2
bqfLp2ZpJpVtKK7r1rgfxnvLaXIHzYeme9XpklEhgZBHBm6v01N2jYBkMTPwcZR5K28R+l/NjyDh
D/rFzDLPBc54j4w4JB1pl/QYl//AfX+Oz/NVRkKtfNUG3/Cwwt/HbIaogEn6FYrcJLiySWx2/2Bs
MCaIGRxkgqTEduA4/tKRomkyKw2zNc76Y3Xu21qAATDMFA0QumRuMXfDcFrIotfurXtygdOIcHjQ
2bbGRt37/lnHOGhKNCNZMShR5EP25qZiaYTf6wzh665+hKPlJbFUQiMSqnMDly+K0oT7SyA5BoMq
ugyQMKTTIMIVYXUQCTI6TtnmuBt7G8v/p4m8Ubcrss4lGeFP1deEaaHDD/ne0G6raySZd0WhUrtc
3uiPFhdRF5iQJYEhhQoxFTI+Ki8lquXCZk4fMndkHrXK0Di606lN49wmaT1HMEnj1276AebCLFkv
uRJbew7UwqTc994NoJ/1loFnNnmgaOGdAFT1C3M1hPBVMqrL6+QWL0O1XeS2VJkWSKbYPX80Dk3y
OtjQCs5qDmfpP03QJjcsFhwYBOrTWKtE/ZTP8itGi/qnSF12xJ6OHXzocvwKlOW+Z1N/tb46gTXV
vH4sdrbyuaI435Ial5FDI8KzgegZ+SWHyrcegxb7Ec6gLoy0tHAiSgttxdP3V6y1s0UBel8aTOnl
NzABovUUJw3zoweRPqfP1vijyOiY+0zJX1QaN2HDSJ1T3wUvKUZRlVzf33pe9DpSd4OZ1ZdzwjBB
L6/sz7gANZlixbvl3ebo5zyGR2uJZ+eU3DbOuVR032KXj29i4WTkGOYTyH6rkwXJJPkVKr2cMVFu
giQG07WOAKZi41BHkNfKBNeGlRi9wRSFtMKdn8+A8nm1rNDilf9Bwf7O34rbp/dqhUS2Wp8leTro
l4szIP3fSSje/zHRKzq22fRVZ0MI2x3hbelY78hVEmGm1iTJo0WpbBOFHJVBlMuzcNkSpVbZvNqz
NEQAfgDTx7biJAxYcuCicSElByIvE9D7VpGq0zawVIxj5iNaoEtV0obCnH5jaBaYeyorTkTibnBF
kPLA0Yw103wznzzO3Dlf9zr7EeL94v2nDOapE73B4rVLuRPVuuhOWkYonJB83m5vaWY6bKnKfBH8
OdXeiNRlvUISDXnWTg9gkg/zXuf2Fj6kExjmE0Bvgnqwi/w9tiMtZRRA7VIo26fEE7uGtO524ZFP
mAsEKaiyQsUos2VfsWO3z4yDXe8CCHWagG4HYqauG2zPG3dI/2u8V4i/xGCcnrSSp54/DpRvsqpf
RSuiU4YoO1loMZzBKUaRznA4+tic+/lRfbqX5xW4gyzI0z8PFuz/C9Ai7z4v1Fvc4Z+e6vzoTQzd
cEKdZkZnnAxYSRXh+2OLgY3rdv0gMHEFCWz+iNaLlDr6Z8RK6lFqRahfHAGeca1D7DASTMjet4Zz
yJcSF4jeND4557unhhe3LacR2Xb0GP7zLQcu+iGOuKVqCryO7eH4heSZwu31+8we1OXYgfevuFys
dNUPuRG41vbtYg2Cz2pEYmMBvOrBvFcazs/dpg1B6u9DvO1/RzIJ4CdwZ1ncyzxtzWTXLoQniYnN
wi5JSIAHX2DyNW6OuKjW0RjGUuRgfD7GH0nfQITPkPlCr7O7QWATPL3L/mI/2xUNgaatEF2+Sf98
Zuu0zD6hkUtirTYnHLuKC2AMS4Nn57BPcBFakJl/1jFD42hyUMdQX3uyGeC+TpJclvY3WVFrJ95V
Z1n9NZzlOHXEOQwE4lZsKiitEmFRsv0nJI9ophuQOFw21GOSNyC4wl3adqhKy9GBzAKI3nqPRBys
rHkUkH9BObUItxQ1NhCRDoTjC/Gj5vtADvj8eyu9eO1kRIgu4LlHhsmSXn2Luu/W7tiYmNADYdNM
gklpwCKDF3/pxeLNIy0M1Dfa4QihfvmwRLKYEE18Mv4umcis0+or/0jvT88ob0jfSWtUEJC0FirL
Dc5BqpDPcdjV+ykt0kwNoocovhI/dOd3gYDGtOeZ/y1H+LlgggOr/bIETyzcl0IVs26zAX74PQJ2
C/Y8ZhmFWiWCQwt/9hlfbnYohJZRM7XK3Yjqz0IjqDWtsR3DUEqvv5aRSjvfh4ujjfstzp0/Of7I
zrr8dxhQK89yU6KHGHNtPGZL5levXBV5HFc9Hq0rtY5UXrnJWSQEU10C+Kt0VtToLB48ClgiUs7q
y5FqsGo498sX4h28U+ANPRYqfDLUq95KIsZQkvj5fZqSIZYAIZ8cCW6w69s4lXWLJR+u02TfZB3c
2BBn6aIH+wpmHYNYtz4JmPruy4cIiHs4On1IkMAvHo2/ru6rh+YCB7ovYYmf1quUqQbkMnqvHkAR
3JsdgX8g7oveCZEakvk/1e5P4S/WoiPYiUOXZSbG959sVXS2ZHYwRilQnyGy3ntgrs6gc6I5AHrn
zWk0Bb0GzXtEH7s/INWkcYZsuftYRWbHazTNXPNXqmboL+whxzAyVeeAhzSLjy/B7a+SluVqDGJj
jt/rfV43RGi46OMoiiHkYXHooelJd0FiOkaHovqZqSOIDrg3Feijfh29Ytz3WsO+vGOKm6pZFlcF
jxrzpIjdPCteWeS5XfK5UuM6UJdOO6t1v9KNKkrublqyE94Bkjm0IT0SngDhdiW3zHnj+bb7NWXz
2UAddmr5zRmjm7bOhu9MVvyjnrikHz3EObq7mDdJEHjBmwKSpcKh7Zhy3/d5cnYgmUENxg4fl2Wq
wpfCyEK38sZhqd+XH0hrSG1QvFCLTSw+UBxO46JKmVX2FMpgUuV2PTxmNzXSfMrHCh0/WZDxBZik
r9hxk/jINME56XM/Yv327oGCleTnimfbvNLHKQqsvr/phxqu76Haew4QfNgzUvpzGa/MSaL0KTHa
DmgFerAm5XqRZ7JR0Sdqjub9hgB3ImMtOmw8oQhIY9s8mjG2y6FBY6Ml8LV9wyGS9UoC13VLzkC5
7BRXF8aDIi1227FpIBfKK43gBaTxZJsYpNQr8TIWXwvqTUCDjCHGgi3T0jJSdYAstOIgPh6tgYJV
oNv2yHy0PUTnOsRtFfktx4Li0kdNCDFnqCCEG6YumoHvvLN8jvBoKzkGoRiZr3R9QPHbRRadj8ci
B3unRe11CWdQom59tWLc2r4gh4vKEniFmjarkcHrSB4JsZYzcb9KR5yWxy3KkLZuPbB9WVWQ0Idb
huCoJOSRgkhTz0c+jwpBz0/c9+XT1OKyGO558rdzcz5f/Pv8IoIbJnM00McjnKtSqCHL20bpmkYS
wka4RFqCA4hpuNHdRgE7btKRPYlV04D2Gld/YKN9Dqplsn3jPbn89z8MiaqUyR2zQjNjHqQ2r05t
sq6fzyaUUXA7YEzEMcKgFQ/j766fQCp4tz0uOwy/ZYfUW/vFgDRZ72gZd8JMRH8GAL+190+QMIHv
Kq1tmh5dWuu0sxPDQ+fBLzM343yy76sf/6Q4KVm7d+YY0hHynx1zoKFryhpNPATN6rSRpP79dEng
6RQHkT7insZT/65aLJLzcPXB82IsM2Z4JL7JynjQEVlbsZjatDxphcysmRZwiFmhqo9IsBBW0enJ
Why9lVSkPEmfJXSQi7WIO7JRXM3Q718ZSRoGTpS4NwKxl1DUqdkg/klkyO6d2H73fqc+3esK1mJh
V2mARXxhSSKKud55CMdKHjrUsVoCVDQOcoLlyB5esjBxljLh+klwbAq/7a2/vlDG3KHr8S5bcrAQ
iKvXJ4uYvNOLogeq7Xv3akxjL58YbZZkLxNTlH3WwYJ6SZRmN1ulr1MpvSBwQaoWSsSwpSWSfODB
3XXCy/dzPl6ghc9REO6P9FLVgQq8OwB0JvFmDfSk8nD4/sEFn8bYarirrdBRr4Q7kQWeb73r9Tkg
xZSeq7Htc90+Xun3MnyYjWlZ5jxZpvNu37hXQNmHz6IaIT86rULnc4lkPVvC8XJELWbQ6QisOyu+
JNN1rthbXDg5xSUwG80i4rYdI9sOGX3kXcz98VY8CriVL0DcOXH47k92WVqALaHXAm/OGLfmkdTp
bmchEXSGRJY/s92bRm5aUJ94DfB38VbiURAJnsMtxEdJh0ksvya7rJbKNk841BNnSmvYfUR42SPF
x+L83PvFRORuNipDDUqYfQrODlrW5EpfK1VXYJVTyfaKuUUWA5aeVgE9MYOjoaogDSIwUu9om1QS
iX02OR45nm5/voGZuJxsdT8MN2CNbmTDLdDSi4zOS+x3A0OCQdo7YRM883G+08ACtm9+RZ2lXrIf
SgsiJPWheGVKI+RtMW2YGuj+NN1fxSIq+3WhcAdUxyNF1XXQIBc0uwnRZO74zqC7rC0Hq9osvsA+
iyUTZbtmn/Ouy3hMezcSzoPNKUqfi4cOL5Y3S0zV3lXYb6tD/jpqhcEtTC0OIGnWovsu7RGJkMN5
np6kGjxp9k2mkRK/BoZd8cC9lujo7KJzWe8Wnh8Ap8L3Us/e2jezDQx+NYy9IB0Z0i2sN9YndX9/
/m3/umrE2lE6USU6fhnFJZ9yHU4L7y2Goi3Iw6Im6j/enPNo7kd0Z747mujX0NA5JjZtCgQApoUy
t99kO1vkEzc/6xhcJW9dZtQRI7yFYG/Y07jZtbjfdUyhZCdrqD7JkY3L3o5V+4Y3I8R0Fw8iPVtO
RgXcRN7epIoklG7DOfoFx5yqK5VcW15j1OPp5Xn2B4t4dnwtE3ZCyYSEw47ZzRLvvEKX2G2am4rj
NKuRLA6o0Hc+nhgcq047iKk5RUqE0CwPlAhTJ8jaVzS9HFFm73i1/tmVZeFd9wtQ/tLMgAEU4wBB
5EWYGEVMRXALvWN2EfzbhYVBmPVy09yKcBznbsJAsUsorTLTNWqZ8K8OECJlja/jYYl2J8f9HtrB
1xfYiBvg4i5CNywGKbXM7pShoPuGVRJ04TNhk2crmUnXnJ8bI8Ey38G7Kxxi5gnRPCBCkBb9Rx2q
Xnyh97zW4DngNemYyKVtF/2b7u2WDLzN9LoRKI8fzVYBltD5Ej5UoMWGfw7Oh3m3eiZj3DU3paZB
OD6yURGs1WsF5XuQnvR4PjeMXCz0yN1FfZ9GqEn+smlvsL1eOZHSmXomys4OC2pxiIFjyP7sGwOj
4ECdyk2l71n84bb4IQOlwQuwvc6R7DvINQ13QrRUcR8qisLnWt3kdupgSnScOFQpVE4mOduUWLS6
wkCxQK7Z2Bv1P/oz9a6PYt+UPIC8fROdFb0WI7fTGftUJscElc6eXTF78sJ4BMt/Fqo4IZxg7W6z
bXZJP9RYszd6JauCH7Acl/Okml0ZypWiB4qqXTpfH+9UZ2IBrnp4zH+k7DdMQuNQepYyW6nw0yI2
6QTrGZCBWU+kivKvckxQnrURDUuSdpkBzGHiD32ysz1yzOayBYCgUk9upusp0X+zoc3EOPzHCqyB
rIBmZgNT0xZuU505ge0sUSyOhi0Mj5jQmqwx3f3/wCovkmGytLuMK6lLvqVVq+bjzq/3XcMe6gtG
KZcu8SrIeKljr+6xrzltUJ2KJkubMYTyZrysMKG5aHTevpHFhDP+xlhjWpwTyidr5BevnTGBEV+O
N3ZF/5Cz/2XbTOZnaCQ1S1uqGDlwq8cOaeWV2Ev6Tmz1nL7wI4TRquzTKXvqXKeFZL3Yih0rlCx7
voA0WuLc+3hRX/Cu/NNYFxl3HeP9ATbR51Sk0ZeFlZp6cqR9kWtI+iIKm+WTcuA93+UCx4G6JbHs
MzvbV58fqQczCStzn7lQyWHNA6yz6xSuPlA+Kl6qX91JYH4L3tH7KScRRUcDa5usn0AuWJ7F9/ny
0cLpjjBa4Ool73fL34VrzUu3w9wLaq68tQXLECHu5CDNQWLbDo11TNzXwSetoPGo5x/lGF9D6gaE
6flNDsfyKPzzpORRcQM3BFnOZg03v4u4KKEFVrIVN20vmlrpC000kZcPML1lZR0mXky/1ehVY5yC
uqvaWnrBYZSQzI7H0uj+AoH7vhIVMAM9loHjXOgc1ZWcGc58HgWziB5InbuLzMOe6wvY1Zq5TGLk
lF/2wxf7VJpcPv9MIkCCUsyYuZCiaUoNO3Bpsz52JSeIG3Wui0V5xI17LjGgrzlTmEmQr8BBV/s+
nMU01LI3UAfBrhnUy/bledX7llXJxGsgM/AQPu6nYAA/9LDaO2QCslnPGxatncsXE0iLrgSrxL4x
k6fbxK7uk2sVKURLJN8dSfv0J88JThMwf497YvOYZq4EzaToDrh1rRV854MqDROjZ4h7c+eaD/v4
phrJlw/v62JreOurPX56eSOrtSuMQ19tiwO9783ntD0wmfQ9M0hsfmFHaQdoINcGBXMztLBkcLaC
MxKXu+pLBqLiH2hMRulyF8J+DjEEtn+pjIGtTv6ykDBPbjvUzEAmZCyLz2kICefkPinx+K7OQ0id
M0aHBy+rDPUotGS2nyHdgyJ/SjFz8yTZ/BwW5hKNcVt4tf5SwE3dLRvtVdQA9IYge4H+vRrkXijY
FXyUU4FKf8C8XYmfH9daLJCc5pbccuDJGuTCuhqGks2MrNq+jHoHCyyBcTFkF0Y12yTzP8z7X7GB
jASnPklQWW3N7/MzpGlf9qzsftaw6cSpVp6b+quXcaXrM4vUIsxYkTGXSWCdb7PXsZdrJggulojR
bowyf/fK21xALZATM2gtMz4nVNNtBL3XTp0gmHdC3QTf8/3YjzorgF+/UYTovONqIvaCytDbY2g/
91WbPBfW+62DU7SOK7IeiHkq41bp9/Gm0J/l3wxnMqpI13wCe+iVNAbSIYRMmdz2Pf7+kCXI1DnA
zG8ssbD/M3mUcllLcYK22H8Fx6Gn/FTYZ7Fs7Mfk+zoP2kd1aPMUsp/19GGW/obB5/GoqGt6aISc
Dq+JOYaHhmSx+Pt9YijD+LEJDSNdCOghcMg/YI6jd/rz3EXZS+lH6MgJ7vuf0RNTNUKc7+dZTmmS
hc+Qq0kE/VZ1mMPmsoxI7PyfxHBF6PfrhrI20HojIJjpiIWZ4xSzVM2kD6EmYpBgYfAIXxM6JZnE
nUdrCY6uevqUxctsoUXyL2STD1LPfKLS8MgvLRIteLaqfcgNcRAX9qwBsKO6vDY+z/jxr7d4sqD7
72M8Un5jWNyLLFd/lnBDSDZDzGlkLIrd3zv3f1x3QjaMe544DEaL4h5BgNGDKhS84UozHYn/Rjyv
4671tjgbM0VEAZ6sFVDYOKnT9quhUqmOPyrROE36GiP+Z/t7Vhxik9wkzX64tXZtYodgTN8jwj94
5B5tvBCnEL2hdwTanIAcifmXEdycKpgSWTBfC2h9JYFXjtMmRjMxTQeyLudeE8h2VrJLNLMfUPIP
KCQgOe55kehd6caY6osagzgc2Wn+Ol5c1Mow6bhVlkx2aoOa8Z7FU7WXM27rGaeLNztfLwfLkPsH
G23QhAeySm6JcwSNlRJDGIp+Ub5ToIjqYHrCx1MxO6+2zsNk9m+2uWOYK5ziZoL64nXiF8DOSx37
sbVbLxryfdNp+oOjVTX262DTW5ZJYGTTamCqALXYXCbNmNrkyO5/wxr8l625bB1bNoPOxTpRAjan
5ywMnB2rlgX/KKjsFZnM/ttwt+nc1OQF+JOR0EK5nsjTQ+Kh1Ceo2721+Pa3SJqlGZtPfcnZJtZs
PMzVdjpu6jV85tmac5utpMZpPrbSbMivrrCUvL9X1ccEoBA/SKf/Epcgx/zffg7UOwHlzHK0ZR4/
OZZi1NAOzRVMzF6DymAEk7UT7wOOH3mNn9ygjp1Hm5xxuURlJrfWjJFt2nIAM5WtFF1MpnCrPGXP
/aZz/8P3fJ5/H5+Kz6H1/j7O+V9tH3GSU+YH6ne4T9JZX4YeQXuxin0cJbQ/+5CxT0gM5LqTj3So
9zgTWxBWZ6+0wPknQQxmX/shcEqfT0MM8O9ljbfHVop5/QVLiADIclTpWdBXnAQ+0h9qDa6beLZl
r81DlXoC5XitnEkuw0oo7YVjptv1ALbSgylgQAXkUCk4BssNArt8zkgL08GcTY+xN8Lo+IClA5Au
RRLTj+HLCZKwMu0h4tOvnnWEiGYjPSoucvgJNzK7WpEcgvCn0r/CmUVzfMvVl0d2DMfRwu7fEfyH
l1SfSCJSLgNQPi5yamaS60LUw4bun6YLMhxc6TdpPzDZcW3pK7bs6j3SZduAgUFGmhfkKk3CTxzp
TzoHEAxrZI4m1MDHSOFPN5mSm1RKqbCu5jHw2tz+q4SvGqufz0sNfkxkSFNohOyMr+2m/5tpTtrh
fxSuEohHTDJwe6OZ8MojIJh0Td10ZJkQaZFEQCGCE0CSL8fAoSv41U4p5Om7T5WmK0qV4h18v7Vk
A8huku3e3r2TY+Y32OEWjV6tBFHXT880RBvJcCH1doK3KQiMKZCZEsNey7l8V5P7jG1IRvHETphW
Ble3F2H0l2PEIenzvVJpPK1dt5qsyRBO0A5zpES1NndaoY0cLf2hLVaKuIHI8ayeuveGDTMzFTIH
quEywnvs9X/ma4mZNKGh8yrP+7NFhjUJBzbEwkj9Y4BDplmODRrQD8ompQoAXMqBgztJ0o3jyvhe
+k6d3ERDivRNWLyYfn7ml81knmhS3uq1rYJJ0mQ272OLYDKUFuzTZyslRKsis3uCMjBd82NIOHR3
CD5GrZ8Hty75MByFA7uZRadtLjzy2DawM9GAv6REF8Ehbvp2wBlWCz/0LJgJfxq1Y3Be9T3Bu1LF
svqMQVo1TH90xa+B0HVCxizM/CnVIdAx8FYp4DHnD1qOvMrtZVg/PstNtAWS7foGQwkzTDO89wO+
UTE4M6eHWTIk1rlRj5DFUWdVXAmleJl61fQTSCe2jG177VH1o6xdhmnRcrwNjPgQc6gCIkcQ250u
kCmXgZSoflRt+3fGGzUm/FgkmNMsEeQTQ3PuFEXLqgs5EUdIhfMyCsJKL1F9n4s16/7XXkcKDNXk
9U0/5OOo8N++p64cIdFZn0OKCvIntu/u086/15isoPjnbMvoa++bPG2O6fm4uTY+MpXlK8pWcYP6
eukj5mfmLLGDv9KoZM9Y9AJ2WlYwbXNWaIpgnD5hkMp0jt3HNhzEvJFe2BqX0fFyDQw/5iFymadd
fr3Lxob0yC43nM2huJd7NhtCEIxxNIq3fgN0nTRkkizLwDM821+rBHlyxodxq2+Lxxb2ctv11A5m
2iZALswNa+JvzKbiwMdtRzCN6PM/1Mbds46wOzduIMb7jMEb+UaMupAiICOVa6bEJ4Kt+snoLBPn
P5AwvFYRwSb3jwrF2nR+oKhFG+1gWA4d1PBgQ0ZpUKWY5/YHpXx0Yxk5YqdM/bOCr7HP5ANwJFnt
mqCk3XzNmMP1sqfSmnBggkvL3aX8fJ3Fedrc0CQXxp3rC4f/2dl2sy7OqHdQ3OAD5HiC89hFeIYr
lIfO+JiZwhlHrx8m0hgIrU1GW9hpq7IcI2wlo7PNrpCJ8YVdWXQj2lzT+Je9CUOHyjqdWnjJKC+v
ENT8GjWmeGtKn2izlrcFDl8blmxqzODepnV4sfZJKpHYeQunQe9V0BRpyxjMvB7yS19oAGVepuT5
77+TmGwptDslh1QXK+GsQDKrADIAR+oLsRxRp16Tx/pXcyV64cEFrLU1rUdgCBqtJs3DrOIADwo7
RFrIBUp8omPR+IVIUNPaDDjhPlMBkV9qI/LmjX6haHQdhoVRnWvZSHcKIfUEPSRXMMFMbNDH32KB
ngZqWn19eQjK0q9PFZ/OFnGaPqakbply9NK9xrLJVaXOvwOt6xv6nK+feXQflhSN5+gGDc3a4rwE
qhsSt08AzXTNiZMGXlkSefEsO1frx/8Le3KzoPkhOQX0ZONl4QVSH8eGFFhAuLNOsPdwrNXNl8Yl
/nPzXyOCwfy/lQhxe8odpMaz7xB/rs9oelzsRncq4/s0qMu+xtgM/pNHRgL5ofjpWK6eayxupwyS
wlufxdm+vS+XGtG+8We9IY2Sks6PnsCreFX1UTuKHJ8P4FwGMHOZGgKnE5zGKZAq6z4K/R3rl7ax
i61L+pKCnFZbhxAaHFu6MmbI7yz/CXZNz/OwYBYqmSmgh0s+BA+ROS/uc5jUTSmC36m68JHLvJi6
40pgY0WVjbrc2ywTujeL+9lRWszDfQ1YEGNaGPH5oNIUd67kAHNqSjh6TRkR04Ptd8WhZ/HDyPm8
AHOQSPVVywYCodwWP2WqqHI9LoWuAlucqXgt9oKxEIiajNGYHGdtbvc4/rGUq1thm7g7XIecJh47
lGbFjCqR8qG/kaSb/4TDjWymyvfluzI6ha2rrR2cnZEz4QIcNavBxmvvGG/BzMRdVxnCGARIRD1F
PHoRRWqgDKMxp5vttZMNnlcc4dW+9S4QYRvQp6hzsYUXRwOFVSqY1YhXU4Yx4jqhL2hVjWVfgG0U
NcwYEkbs7AdAdBztoqp28pdoKJj0PRmqDx4hY1xzTOdtDhr8w9XZ8b8nC52NmgobngSUr97Gq3FG
LzWNM+dk/+wiRlkmrGtFlb6fa2I2Ww/fjxv+rl3gfM1gBeXRzQJEoTkxtOgz1QTvRAwBYEdXwGpx
2bWnWx/rHx3FABxgEw8D19Mgr1tHlsZSnEoc3j9tcvVaeV7ZUaDW/8iYd8EVj8RSRTMc3ztr20sM
8TC4aji2fYRzTkPZvI4WfLCEfQ60QeeFkiADD37xImFS5uxSsXCMlvVqJ8677OgGIpyBmofPZu/z
INC5ufYm0MeW17c127bw/fAh/ccY8CBSbX/t6+Bx4abg3EcNM7cb8XZEGAM7agLaLVoLyMVeBuwO
4KgSyL0KFKBpRGWJc0r7UttGMcYuETmSeq/jBU74dcHsxNZBLVxNMLlSfwDS/5uLQGCgQoINMUza
h/eJNUGjZgdoG5nkof86Tzg1L7nsBPqZHKKeAWxYq/hYSCeSb/4tunqKuF5Cxe9kOAyQOGZilzKC
YrCyVWruH1J32LQ5IUj7g+rcjWzoXu9Q8JAP790HW2Uu/WjuQnHN6RoL60MoUm9X22eV5PyImj8a
vW4o8WnfOu9caRwD8DfnjjlCtWnHSrAfy+36H/GE25im6B5zrwG5rHTNLF714F52+//OJAAOr2ab
Eu/EStig/C0XkWQB+fDkPgX0DyPyPf3nu5NT+EYvX+oK8Ydext9XJdJwr6O3XMu26ahBe15e63sn
SsRGipH7D6VHfkWc59Xw+usozCgaUXo/71XOCSA6s3AfXpLZSlZrCjwPN/wqjeR6aHZjScjsKxNB
715S46FBdKV8IrLWbyicI33S4/s8b8hGtK/N4UEAVuXypFlD8YS3ZBILY4IADddHMs9gRAWKKu1J
Wg3WDRMl09gvosNVeNNzc5Ak11tNHOTypzz61Q6IS2VQtmUFCd/nY0nnBwZ168nP/nzMP+KUZP1T
bAUfEp1yCen3NgndffMItHZvE3wwn4wd+7Ndv8FDSBdaHQVrIMr6G5ZHJh1LBsemgbZNdz8HyRd1
JX1oI/hB69PVK7Av3xke7bukVlMNY+0xRguh4hqbIeoESLg76fCfYsMk0r89UwlTERLT88M0axyM
KI+ZJOM3RH5y+MvKOCrrDPb7rDt5lKOhdMA1jqQvTwDYG1Mg2+uPXbsGposTMAHPlokXd6qBIm11
Y6CA44t9kHmueGEUq8B9YBTcJ7m4t/T2rKZADM64/2iX687BWWWU6nBajuYo7orNGeOcLJfIFMqa
rVorOhUeGj9zGLIQbHwDdgvPomGhdMvG4R6XE+7qCD7LFgOzmHEAJDhG4cunTR3Ft8/50nJ3bk5/
eAI2UOQA58O8HA9/GajiWoCbxDw/AyQbOPitaDMGmJKMOY54+Ket+5JOo5gtpshJ85ROKU8P4dBG
daPkj4Sw6tXbuHpMCiTCkdaagUbveZF7spmvxpX9pjLjgILK2wDCwRfVuK3KWC1uo5wonPrkRl/y
xILq7qn6T2gE3lRd4j1K5sD0ipOaigZkGEROGp/vtscJ2cU6wHn+xDU+sL4g/+P/AGRuNQ4eU8K9
LJ1IY7mRsv96Nj6JK+YplkATtXPg8WBQPI3+O2D3q5/VlsuPoTEv8QFhJSMxNX3qojOmLxkO1TEG
MfCsx6wVN7YFSqo9Y74q3snWt5Mw6wvxtn8Jn/yo5mwDn067f/mdkudZRs/QVfapnJ4AZ1cpf0MU
DjWzpGidNjLUdo/5vt5nrmwLGBFtigGicKDHdphFl9sHA9Ii6X7L8ptNg+hrBa/z5k5d5B/ylFUS
s5v5em1Ohqi+tXVQccVzxMkarAGEspUeZC7oZ8nvPILKyoQ9xlUou5K82RUIxZAHiedk4GkrvBbw
GPwt062LDOPdoxp6kzJdaLdoTzQ8Gzvk3y0X90KESnf0oYmxPyyRPUSJT88iG55/UJsl8i3spkWX
EwOMASD5XuJtFpfTbP0DUnFCqRElgYiVibfyocL0FX9pQmtC33TPkpivE9lITJCE9jAtNkRSDD6b
xpLwLxEL8ljaWrucFHOoIOX+pGk6LhhyQtIpzWhd+WmkrrUVBYwdueKvTwtaidix0XpnBrjZpu0+
4SrB+sfYWAjLUu/ctvftKKi9UZyJ8IDbH6A2b8ySzCwye9kjAxJNLwZgDiOkOzOmVLt7K8tPiw/+
ryXDtOGQof48u1uMrBRqg5uImlC4chBvzkw8r9HMuJePt77+LMw2G3h/AkBxHYt//Z9ASxX71/Qo
3CrVivClCPawD6nthzirzn7XB2rJ+SnZzWxmtU/NROOH8Djltjivo/Tgnaq3oBZKWo/7AwudOaUx
O+9/UjtjZtKt0ZZRh/Y7ib47ZQVdTD0DQxRvCaE8hW7bR2Ovevsm9bj94zAYtNMtJgRsJDYAo5dB
e++bXtvZ92cwy9tXCcQ6cDnE0TBNmXlc6EVENn9RdWhe37AXFB6NiPeLPVO5RzpwjytCEPZ+vvEu
IrC0GD4hSFw5XixU/R1wMmZO7sTdqYkVg+ipT4/ySFtYyRIbeP66BlEvLZJaL8al3MbGIwJRPzVO
XZKGe03+eK4qehfJe4h1+1qJNtGFZH6hE/4uSc8yuDev8D1JhoPiBcJyx2We2nwFkPnclbKV56qx
ZAyJAoMxCDm6urZGVmUWTDy95FYVuwI99UP6Y+LYyXzYFgviEiLJzOAM55ll3TjePgxcJx+Hjg2v
QIo07qPC0f7BfZBB0EX8CxfLLBFZDfIV2el6SFKjYiBTPrUdBQReoLuryCfSaCy7/HFSedEvR3Ke
pmZwnbpCS3EITavQweb0Vdc3ypgG2FThsVawSmtdR3DBexFzJc4ARNseFc2wbNKU9+vpmRfjDQKt
UYVpOZZj8rt7jxhtWsGO2hOBKnDYuKfW79f/fawM+bUSCr6XXwnL2/3R9bKLwKd31zF5dlzAsd5N
BrJmiG7UeT/CSJexdCLAsDXTfQCR0qm9N9cE7dMkpuvgT5TfXpjOvgdqTP1F7tHRyw4Gp+91VG+P
AFdyWfUrzFEYv9NmtYD1RHqHibqySP2MGz0FD5ioldxig2iIGdYKG3ebq8+K26c1KqCEGzlYFYYe
2n23aWyTDfS+xjMy6zekBblO//5Tu+qC8BGp5MCx0X01jT7M49BeaOtiVBosiCjGedOUshioepCN
iMxVHo/37NOXl9ejcPGgJ1YreTFPDVfOft/sDoA6/zpB8xZ0FREn1/dXwwqngsToxB0KmQOOFBg4
r6XiGUFmWP0sTso+0Y7HXBzBVKJK5iG5Oyt8NFty7Q/cpF/Yir9sPxF+Xt1NFYoS/1OpeqCbAmHn
FcfmJMz16jf6WqNn0inSPJorfsCkqdl2hqwHotWmI7YpTVghERYMZTqKxQ6Gii2oJrRvGPCGY5Sm
OC2f/AvqId/VAhVrAQVeBtN7GpPWMPXp5UjoN+OpXotKXJQLlGegSxh2vxY5vpTt/LMdtFmaZGh0
LRbHJGk9lVMUXhffT1piFNDRPPYnvEs1duBkmhzk9VmKBKX5O5ji5v0bJNA4xTde3jG3/e98EkNr
tCypjegKR7JOmPN0uUY2QMN86lq0Ep8WeEVX0PGCt7BPVw/KpV7SH/UUIbD2RNrfCFz4WRNS9QL4
ScIJaAlyj3N5eX/cRY6V0USqucCQ97ES3KvVqI7X3DMRKHK8jwg8udJEjoqsGUHTImjfcouS/ivM
H9alOQAEbIM0gOJFnxYVzVlg7mKZzStR0OdJCJAc2Cc9EIu77beHC9mD/AhnqWuH8QS/h0m/wSk4
vWhyZj1zzq1ArQ5bm42le80keRwhrQEjRrlvHRxogjyVAwUU0k8TGACq+hnVm378vH8hsAdx/Q5+
w3pax+kqrxG+3b/4VgxBOf6AddEji4BUa2Xqw43WINNtHOcr+nVje8aOZomZ05YVNYys8bKCXShk
Ptjq9sbKBhrylDgOkG6KkYErB5dqj96v8nLws42QF+XkyfXaev9f9KYEKq1CMdcG/naTfYonaTqO
xVWU7v77V0W7Jvx6J4Nql53mUCLGgO1q/Ft4ZJSWRm4EECuRAEwOKmF/Y+8btLwWEOc5eOAKB1GL
p2R0mrXspd6TViHFfg/DeQsE+HmwA5/xuIxgkWprzvBVB/t/UQz6DQON89DQlWpG34crsUMf9l4T
LlVw1KKp1X3ZPQVFii3kOzhO+c+IdDVfWqNrs3fIC8KUcKgXEI75ixYQvvhnet/bQhDvwUNYjFwm
r4XoDsyf1xyh5mj47DqkJjjNcnBU1k7IqORx6JWFqiUJDo6+hP7h57FmwPG1kstGWAQNh+gbyOdc
1rEXjSksGAyWg1WogEjqzqfYFBOfwveNkAO2+GVStc8m8XVDD4ia95UGJnQ+Xd5iBk9AIUYGSzKC
bBqQCP7baycGN6yNal14jx87yaUUeYkESCZ5/1tC+PISNAu/WO84uE66PWcF7m69lMrTpfsawisf
KubsA0HzyS3R0ffkus5NkTsplr9cp+Os3X4IvqVM/HTBQeGnLsyy6qcxuXetmPld4FBED5SqtWmY
JMsbVH+r1dwmUe4Rp7DJFHve3Sxybs7gyJl6xtinPWZ84tG94k6cB41wgZU2O4cy1FedXsOQhTXz
HxYFHga3/plmRGx5nqhFWTVci3Xn3FC/cgqXuYkBJ6YGGltvqag2i40ijINeB1/knsWfeN5Zx5KF
rVez9PFM7E1eFtz/KJ2uZCEv2d6rYLXI5IKBXjyjU/4BjfJCXcSlk58TeBJlNpeh/v8wHRof2WDV
wQeCWj+zUCCYMeRsn0xnQwdfql877KVDbxnDkAlIA2ltxTCDP+4DUg5SMW/FBewINNjFg6wqNyrS
6uY++fYvlL2GQqVgFJgAPqm4EcT2dHf2j7k8/XjONfSk7QqghZQRxkAhYtWFXgMunK4QanQmYfsh
pSf+im0f/8AwVEvto7DUPSXp2piws9Efd0rKwGVtJD/V14T0Ax9d4vzqaaQGdAp3EBdooS7thE+m
mscG2iraAebtfMLwq6tFPTCYt7uZ4+M93n6UJsmKYCs4rouMfhGnU6igplDk2wKj6xW3xzytJXof
Ua+1FIBHDWeMESMaXo4O35oGITO+9AA0/JV1+pHpzecMzjEJxH4Vu9XsudwwiVK1fB7+KrcRy3dg
OHWPdepZbSO7YdB1xs/d5JpgN0Ko3DuyopRKnrMHYwc69FwBIoVBG2+mHftGqQnYRx9Y2otEvZzR
61SACextxhMrZM/7eMFptWv3BxLr6/sQAiKQYLkGQoE4AXWHTRwx8EDNMcyT+YsJFNBAXz8mIL1h
JH7GD8iKH9e1iv0H+uqF4roF9THNXwa9LQFOCEYEsFqJx8B4oJb1GetkrDoh2hlFGDiZgB9gaV/B
RtfO9CbLh6k8h5Z/Qkgr1CpyYi+OikykBiHNXANmJwkfuQM9uYy0SCRpiw0ndYta+Rmlh6GdZF7Z
iTD9QqulTCybX+f/DvJqoIWxy5LoyEh4KMrxoiOwduYPooWqOS7PAQHVCJmfcC7Vit5caY7Ia3Lx
8iWFAZF8TvPqEzBYrFGVUJmCoFW+eXdr0lBknst+KGzUY08Y6dMlDbf4hGXTIdh32DToGdoA4dtc
fKNYCAUleGiGA8tqdkONnx8+ogAA7S4724x4CX1EhRprVyNIYwN8kOf/dp4kSR3Ou8bdolM3TpnW
SH2ndRQxx47AyZxoFGUka2cGDS0/jkjdeQoKMEAFNhRI34pDsWGfL4WdiKPtpGxc8ezQoEKnL0hs
yYl99BxdrLTTtfN/0eLSAZR/HIk9HWBcZ9VFzpqoxpl25rE8QcJy3RLGXwGpyFab5pWG90p5Smox
h3cQdDVKEvc3x14MRhXhbxpiJ5K9xuI3OEgdL/VJHP+q7ubE7i8O3/yPh2OMereQ+uZ9/DEptiC2
WaXOSS90l+wws3iKmyPtpxZeOUT56TV8bIWVEQouPdPCax4UmwKJVR8lZ31VreXdAH4UzDrWqc1m
pP96mZ/5vbAsurt3Ys9/tjBcTjR+r5RtGxkLA3WRhIZqyg5rfAAb1QgdKSMRaK/hhyVWkN99dXE2
g2BK2BqxxVKNOuGKbeA3bN4e9aaH7RAc1Lz9xRzbFd7MwMyhrS7kjPGH6StJH6YeKWyqU9WaDUA0
J3bNsCntWH4Pod2oGYUrGr5ORBLTwff20kqGecnvvDMs/IoqW6EIJXijQRct6uVithgcqF5YFdLU
aRk8XMmz284sC9XH/ZUnEsYXLfCI8sK+OgiB9dq7sT8ml2Ae3E6V1t3n6nNVdXFFs1R6gJQTMx3o
2xrm1CW4dRv/Xp4ZvtliterGg8uoyHp3uHDz5cPJ/hZ8rQpXQ9tbR8NWn62HxrqHX+6qy2W5S4xH
zBU7ZA4X/ubjd9qjEG7+P86kJfI539Dwq0q6LKwSJ7FyEaE1PG2S1RfmJoTjLg3CKsQkSPfHXGSC
JlLY2vSQU96I0PDj1AKWlvkW+43p6jOnwMHcpJgR7vulstaT5iwXJh6vmr6OhZ3MU8R8cI+p49A8
CiUmJ0bP5p9fgWMU754tLM4eUSkGYuBUR8+PNXzuWB2NvF2ZvQamDuYH/Y3jvwoGOEhzKbAwF1ay
0srZYQc/x4xbcvfz64HS2VV26DegkM+SoOhuRv2uLOGsdm5vZaiuh57xLk1Nn01wLbHSma10SaUK
d77q8YSAyF1BshHqDUh6+Sm6HrGuaUQEf4S9dvb6Ixd9C0HUFvAs/D1vh8uKXgs5+dnoE6NNVoKe
jU8hxhUcBASruklu5kieTqmKAPItiZPL0yR3OZjq7s6Q4NJm2GWEeYauyN4sdSS5EkzdWlQfUsW9
ASlIYaDwBdvTLSrgQrRoMMejR1r8cyRZ5OxaILe6qoYhh/iu4ZCEsVnwx+1QajF+MjUIcDmUQSZ3
hfgh41uIN+ufqAjNTeRBkxiRjoF7OjRfp+D++tZPPgdhrK/CxEJQVaS05bG0LIDmoAP7SeJz44Mh
CylfKYfX0oq76B9JfwXTm4f1Iyn/c1Qf+ew5T4FW5iEKGMITLRCCoFvmQiu3IFYpf85DV/ePcgr6
Jpln5ldQ6idrqiNr6ZGjswUXal8jzrytQDfwqab62xSHb9n4DwH5eGoDOqj6Q8ivcNEWQSDHWWQV
P7cW5VVXd2TTpKf6Ky+A1pzyWQBuwssfTOmN6n+6RLyx2G9l5NOnO9H/BNGOXxDSNjGJuv8sIkJS
CI0rmoA5ndfk3i6H+0opI4Nc5f2ozuU41Znvt5+EX9d9mSZ6/bVk0Fezf6fF5k5bVSolPla2+ahz
yfMqRhuoLAj/VJ18T9hTKuVhW+VV4fdHcCEjfd2o6ya3pST/Qvh1o/HdLkcW/gZ1fdJdxcUiPABB
5qf+y80qCf449RXtjSAtXv0VDSnc37wNRkt1Py5+E8VJfzJFyuUUEFJgafbekPWeTzKNped4LmRj
IF/ODe0orh5bQEaJk9P5pq7FvRKdYJwoqpN0b0+OIzbKiZgRE31nSPpnoGB/A/Ii5uMe/o+gUf9N
Tg33kBKnxhZ2RBXKbNA0seS2RKhbvdJyBPcWiW7lsEI31nOqdjYjAVIhWuIOoMjyWgsd1L+HNqIi
a+QH4ks+z1HkxvP1k8Uwj7PkXm5Y5Gwvd+n5VrajHmwtvEki4iEI/kSeDDNk6P/TjeYv3YAyCVnF
wk7mHZhoMZuakja+WwpXKyaAbcr+n9rQmPFZSFYGimWfEBRxGEkya7FzgIju8bAw1tYcrqNxvk3I
ikCUxq8SSCfU2cz8HIyAitdhoNBiC3dp8Pvuym05Fds2hUQc8ipvZgDMAjB8SLkAD7qQbu6bCDX6
aL+KxJdv+98bZApAj3uuhb4OQ9GbWEdAgtDOjY/+0jAVpgEoF635X79fu5Nn/aVAzlvQvdtWxHPU
VEe2y0thrA9Gl0x7CsBhcgmhtU4iW8qX0HKB3fyMHQ+aznm9k7nyEEgRYCBNuvNewnHeYc4z7Ftq
ZB816u6fLenLz0TzVQSKhb0/Ynmpa3gjGjJK9ONweGMNEOKz/2hcBxnfYLc++vSIuv+Fl4l7dZ5/
Unc5bXdR3cMhyyQzlBGXB05FSHtdr/5fbpNC/WPs674n3B3Xv2XixOVMkJPhdpNSHIqMwMYa0V2+
4/5wxq15M9e2WB2ywBIfEF8fvxyW33bPQmzgkk1DkqgHaB/2WGvLgzB7c9oeVx7QUfUq8TQeSN5N
b8uor0g45n0i926H/495jGlJ37SbJqpt3DXWsu6dKNoQSQN++7v6w7EeM94XSJaRQcEYq+/mDCaA
+qstg2ujc3H8jCAeFtH2ybL+XIjhStgh1szU0wUGnIOnXbFNe9kwoiNksWrIJYqIxg+IfWkHyZiH
4Hp0VSwVgMkAMP3gz3Am72lsDKyk0Yunn6DVqUuG4AgYTTNt28HmHB9slNOerrRdbAhe1ShYjeAu
vQ8OSi+TEgp7/WbF2buwMiNr90N1ezjJdBBo04vXhFOWPAKLixYJ7lexFY5uWfRojaZXzj4ULgcG
WNGuiZtgROLpA45vfYwCt3T/htMrjUrYeEXP53/MQNbz12w06BatBolxG/j+HLrjZKuDvl8R5o2H
vY+xHlGINXoUB6brTU6P+MKptgvoNKHTvmoHAkLmugVxeak2mAYS1XQVvBeZ64+i6E+fV/y1RkRt
Z831A/Luz9YTZvxEde6b0puVG6TbwLv2cx9RFEDTaNS07vorHxpnVDRM6UYqnix0T21LesTnrEnx
F6DfEISIWWrzPJxpRlKJ8uPpfSjnuDTEvsg4BlRw00K8Sja1ba7kslS2JE1oB7yx/2JL5v+tSrYc
Hms2AtEXlYf1CW7prp6mH2Vb0e/gwlpsxVYCZbEopAiVIuKqmP5fLneuQNKGXIZC1THkt4d7bHPY
ilbdzs15j/ZiUWZemNm5abZekcqxhW/JZwL6iIrEU7lZTG/b6od/ZIXhn7tpMWNivUo3XGk4BZ88
NqRY0Uieq5RaNJe6/Y5ajeXugd2t9fAIUv6W3T5arZnxV88IUaTY0kWOUcq9eWdMVNLJFTVmgD8Q
NXky+/aDkPtlp1Clk0a69X5M6iybmxRrdrXz7vntAEBPAziBTZGwRE/okrhtbnYIx8mkXvOBDcQt
Nufmi2oSB6JbFWotkPE8rKLAkbbUdxcO9VGdIOHnKtbHw7wpNugwF9dxlj0NspMBjGxyEzyFnfIe
v881ufnwdxEJwk3Ex2ZPFI/sX+iACh2ln+HXe1n47znuuVyvLYUb6hWVLRnqKl0awxwxhgKkeA8F
1gTqq9VmNHXBZ4RXwPH5CMpLGAWUIsSacwFv4tGLM2Kx/HAfAajBUYOJcaD3nQZvi4ls52VL9AHm
84dIDMMnZwrKZWJnIRFpD91xn/qB+SLX6G7pq/IZdmwn7Vhz8MfTSpVOWHIodkw98a/b+lm5zt80
QLc5w/76qX78xggNuAJdIsNLENAmXk3FRmqQheT9qDVMKKkTESLDcaSAQAZgSarWsyz5BKSKUljz
HwANqdIpjnEfG6U6yN3hcaHKa/n2Vm4igJAL8vhip1DbFDmQqlJd6Sq6yh+VHfDU4gsNh4jYZOxf
oh6nBZ4sOegbTt04IUBWfRyhemaEgMKa35vLRDAWK6eDZnYP9YnofiY41ZtgHInXA2rmO24D7hI2
mxVqedqyzJ3rLtwDe9NUKXUPGLKF+CGtCRhMLxVIM/EgNtL/FzRerjSOopxZ5uNli/4nwcdYvkHw
lm0AFIwzzzaZY0CRFNz7fp2iUVkp7YeVXOxUZoDxBOya7F1tEduEFHnlFc4rfJ8jQYJSQH/yuxZu
Dmx2vL0mqsz2tuf8XA0F72xrC73AT9RObV/MfwVBpZrsKdzQKlVJwe0pchR/bQSskjaFZFS3NAaL
dOfrDzXVGq4QI5ANotI4xP5oS6rj3x+wproqokThY2ejsvsmhe288nQG7gN3ywILgza7hTTbB0EX
9jH7Z3vEmuf92zozwhMyO/++gEQsQT77rqrxLKK0nl0Q6HpvkyDAn40eT7JSALMQSDs6iAGe1aC6
JBNkjhygogSMxWiqfpLfvvP+ONNwbjvu33Hf1Lx/9VP42yPZLTUf0IjDriDkwjrk3b/QH3YQaopD
+tf6r6AoTg4bqCH866gvJ+P1/Dbap0f+/vkcf8Qm61RxH5jJ8//L24SlByg7//n2EZaRrptkeGC2
Emdkm6vPLqxF3ZWXS/5aujQAqVZVV+ByUon5nLGuHz6iskdvMy+WtxHlPMNJjQuHo8yZi0SJwHxy
i4KzUzGUEbVSAWo3n+q8kml9aiHjvTJJLLdZnInf0yzkM+B6MMhG9nX1KtXZVmqch9MaoPlhoNYY
09OYP2ett2N+nLiTTUgc/xLc3bdalhtW3I0AzqGsmt6fXhRkA22qcKyjbCLpRlQvirHMRLaTt9bt
a3vMMqlofZbcf3kSbwaw+QbKHfS2fPccIDlTwjuJY9jaDZkvZZoktUBVxRhO0dKAJ6p8MN+n0F2V
If2zPZHZmydyaVPhEqsHsBT65UU+VXy2Ifx1BEYHk6srfAumwj875XK5mBPmihyQX/cBneyZb/hm
gBjNyEvcBmVKw+W1OVtOGwse4AklpkAsJjc7l42+MTKiMccSldYAoWUjw7f9hffZ5oCv0vdBb2Ed
nhHafeaYIfdY5bKSq9b9Iul6R/3roHq7cTUmTC+BuAo/IEnR5k8RYCJfAV1R1FjOs632exkx6WhV
+eJur+vqpwXFfD/0Dx4YZWN5z6WGT/Fje/qoqXwc5fBGJfax4ddOFV3X4Nhq05OmvNhuFFQdEz9p
awFgPnpngbxGJVowtfHEgjxaLiIIr8NzcfVV8DI6we3XEOe5OMrMMTDr9jx+ehAGQYF3Wx/U8KLI
sSUjNRxfdQItr7Lj6d8houNXVbDYGb/8B8/lmTxJ1RNXYhb9/SZAQO9wgsIthzOpzV4aige0Qsod
XV2pgCYw/yigagNFNSITsZs2ONxKG2SuiLo556+RGWq2LgS6w7zAqCY/Ao9Tfh1amTkBTki9PM8h
+RxSBqGYkDm+nZIu2lYACSmoF3QTM15SEhvGXJr5V6UsJ1Kqv23DYQNtZ65EXj2tFrI2ukkTifQV
pZYgI4n3P9c9NkkkxRDd+1a5DueJpNvzUol1ENMv77+1GH95ZoCemnWLGHhcNqz4j9y4CGTN0X6d
qNG8RDl1X+dqHkuheXne1tjhpHG5nqsk/atiArljolvKOPrxCIgUBHxrM7Z25UXtg1JWYpG3UdmS
f00kIDW4GmJT13V3JGDsQTpg+BS2ie1mw53PvKa0My8BHTeATPR9wv61bC4xF0BmrxMYC+2qalzU
zEwSgua6HCgGIfm0mZ0/goHQM41oU5/TAg7oF8rnFQRVST4/qklbNS8fcmec05kN6BHnBzXCNG5c
t+6sfJteIVqi0A3HGdJQ3hrJbNwmjn1lfmE7eYWijZkhkUCOi2pOcAFsW6HxwtoGm4sOlC1oR4ct
lKNPJFUV/Gq26ksnLEfphtTtOThMoDO+544S/87GrcS7/pWeJpRya/UTH/pEbabrGj9his6lV/tg
oJ1C4BOQofV4vTiAsYjep5lkLny247I9kqL9IRBiS0rK91zDBvp3Ds4KYCVxe6OGeFIQkJg4U6dO
7E47TzIuxvhEt9jtzJcwSXBelrXZZo2x7qNHeZGZXouDP99CgNzZLw+FaKV1kQgO1K4D+o1ZB7Iz
IzrHD0VGfGhkkb2PLThIUN74QnhWMxNQ81FBX2BBPqG8CykqW+iOzxsvRN9IDLKUsvi1cQqZi4hr
pRP8LDiDatO7Uo2oEKIMzfwlgzM6u65YlRrLXuD3uPZs5xZjCe5+Maa5TsNE8DTtGyiowNALx4uP
FqMyy6jo1M3BIvOLVyDy0cStuTeRfzKJf8yNmApGQrx5pdt4RPgFGrOpuQlQg+7OaP+eSRNhXWeY
DVFoUY9madeuSwfnCTGHlfqfuzNppJWaGHyMkPyE5h2sIShLfi8KJo6VpIfrtkrdOwa6TJ03Pjwa
eSGGQ72eOoekhr3cMmiMreZGbdA7aXgKCu0U+tDWRRdTLFhKmH75z/8zbFsHEoF0RCiaRpYwITGy
W9n/xXWVzO6Q70bdQB4dHqElqb0z7NgdJPhbb7uVX/4i2nUShjrm0i9WCnYVe38FLKV3vkF4qlZb
BidyrKY6AUugqv8w0g52FuV4wGgD5QAzJ8Vt90fsx18p5zGOwkCHYvrnnPGdHBEm5qx+B+8jvDwf
FKHLL8pyOsC9Mw3TFpx2kh/Ju96JnC/ws0URC7u7bIad8VQ5i7hp2jCmCOhkCVTJAx0Uy0/eQkY6
b+4ZPzEHYf9gu9OKoY6wOBGwimsG7A9RNVLbUfgo/unTYHqllaRIrymZSHRw8o1nuurIQ9Uzk7uq
WYEo7qvV4z/JgOUXoyPnIRQferJ32X8rP5Q/KOJ9mukINMDhNcvR2gLKAqG7Bea3KPOl15DSKsvD
ZBHvrXAsCJIHOddms5KJKVUupXg+z5kxhhw6gyFoBteT+IviLIb566TyPBZJ9yAn36pXY1VsI4Fs
ZjJV56FsSJP4VZl3AuZF5e+Zk48Z5AreKkZiWDkEW6lFu3QNjvrrRcBEsx6OA8DJzlHgULJq16bP
GTpbAIQlCH7p+OK4ipV8ovXEVV2uDkMOZjYBS4GJN7rLHTenAIPmw05WQyDSz/FoNMzu0vZZqtHf
XUojhZ6CgtXk0En+qnm3ee1Met7MeMC1ffxTjpZlPn56yKawVcBPA/G1H15ojZ1+4KZNRvrljbcF
VRnfGc6W3K4HKAZAKqGPTd5hvX8ro5oFCJ9hQNMALtTlYXayAOPFpfFM2syDF3JNkh0BY7/TYgQL
3Od+1OysIksytYtPEr/Mvy7e5tKGvuExQbeO/7id/JAnRfKvM1h9qRU2DFzyUk84DiEhlxTtafpj
6Ij26VPG9t6QlwnZZSOBVcBdzeMPulPsCItJQZPniTwcEXFHnZcmUZXSyFQb25E0ZMX30DxHMOiu
KkFHFhLGccK7h4lm3rPQmcfb4qLs5WzF+wBygO277KoqNLnOESXfMq6p6a5nJFAW+n9CnyXErhOV
9A2d4Yb+p95xz93hqDpERgvY7G1xpbKNfa2nSjV8eHAj3Xqyi9TqCfyhW1CUkfQYX2D4GxNMEW9j
0lnkGknyg2cHkIX7NW9mp7/Be4aLcsJL5kX7D2/88TsOPEFB/q9dfricVbqaMLMEK01tDqRb6aq0
IaTCYTT4Gqwj1BTean0RfLAlTqM2U2h7V9vQh/NYaEzVbMm0yCtGljpARsa6ErKOzrQdVxKK8L17
IpW8WF9jKU1ZZ3vJZ3KuD2w1YtcIEHkhm4YdzMRx9xHXR5OzpUJO+csWz0bGbWtvF0xp7dh/rkqr
PfYhCyP12WOLaN+UTv4bZRHGkpBalPb2pznARmHbBOv5UEZzylw7rs4PKa4Rv/D81RMSGnllsehO
GBcvnJkYTqcgFRk+a45AlIW86vgcs77uOZl0PNkoZY3NcW4bEE3jampTPE5/eMj1aj9IczyGvMZr
dt067kKYPYE43fhvfDOJlsG1GyDG/ibl1cGSX9Bve+HS0PkofGV8f9QLodJzNVx1D9fV2ujjVbWz
k3a/W8YsJIRLdfkmtp5g8tn3Pob2YtE7pPvEwqeC3E5cY2IuIIu7S4DGWli9+5O2QDa4Oug8UTL/
usDJELsf/SUv2ZcQ0zut7N/VAfG3zqWWC7Yx6trUJChdGri5oLKTq9r9pf565E9S7EKwo6qimXCE
jP0hoLmUpUhxM4admjzB7AO2WcFBbLaScI/Ho7jmzILSgD6qqoVml98FuAvL+jcNWufZ/6jvwdSA
g/jMth7aItAvRBDS2fIjNUGdNONIRt3GsfF7+34ydYurgnLUUPrTSfMLATpHpi2e4J16HvwMJ9Mv
0OnSB9Y891ARVvMBlUa8TgKCwPtbHx6F72nyKd1WDd2Jzrl8VHs5R6SiHyh+1cjDAga5YFwpmf2J
bbdLr/GB0ywOxQ8ADUkU71L7MQLRT/0iNEK/9uGoLMCvE6H/zLZ02F2PkVtwyWwL4fpZ2j9xTWtw
Hv1xpm4pkQhj7zfjzooKHLuQFh1x5O6a9L2w4heUD4qkorfhJtBV51b30mMOVpazpIDIMnbHSL7t
42pCZPPGjpbsG193MAonFtzziUe7xidVbs0DssVRYnwaPyzrtdVKDFjES3rg3DFGj4LYLbAhqSDd
FT+/GwC49xDz0s/0BGxyZ8kLr5pIBtqGISxGEFjMN1KoPRCXF8RXdNepqgmHWFthub23x3I8LD/g
1qYEO+xGsrDs95T0sMcBjaHlRtZ1QE9jJjBglzJMX+2a1NI+7UXY4kf1wMRXL+N3sempcZl1dEA4
5+pVlBsMTapbWGnGr72zq4gAhEehLTlgUoj+e7cLgwswLCCS+gJgVlyxid0L0B6MHxzEmAEgLlUw
w6bQXl2KBaEzRGKEJAt1ISoyFlWfpfrl3ZhxbrkKN5aGS6uWy0IYBKeoAegn6XOGV3b0E0vAov4o
eS155tgDkGttL6XUzPiKLRd0X/7tD3cBKE18j9moKR0qIeSJTNcT5VRc7aZWT/SXJHjDkIxxBWQm
vNo7pZ0X+v/6orWBUuIdToN6NxKPJ0wzkAA1ZcojP6XSdixAyT6vfpvlAcJRkAEQuGbrjTIFG7fi
jqdIxUhGMYIJzoU3EODBUbqagXyoewbhS4QSQWtcgIIU9fKDZGPAOmABL51nL115K6as8eWRfAgi
Mtk45DdEMgmH7XuldFBBtT8mguzfmdYM+cJFClc0OoacoKT9L630KeWK9agjA6VHNIA/+wlsgyxb
h3duhebTWNQbmuR8CgazEn/7OMnw/XbslaQnju2oJFaEZfwNOlNmSriZmC0anHIBysdNE3EhOpBw
q7RIOW4+m1JOHuP+ZDRWdOgygMlmwoHby8ne+I4YyAKezBkkieVF0Cf+fZcpEb4qKDSBFzA/oejd
ojgTgHf8tdT/6hozoG3+KYjD5AISbe0m4fLu2rW4zc+XL6Td2CcRHWFuWRX9y94k+rxLfowonvZA
dJkOFTmq1GjmByfLC3OOci8f2OAKVSLqza2E26iV9Ibx2urkDUFNcGfedep8STKVGrf8oDGkI9Mo
iw68eEzLBeYJCtpO/hUMFFlyImMYklw8Jl9SxaVNbTUS4sPTOyR/g4f/gCyNxfnCuKzHbrtGF5yB
1dl05tGDZGmyHTJ5ecWjC8GSriILAjmbsH4DSnKvBRMjOpMqoM98LZqq6fk8UDkkd4Bd902V4xeN
BWT3OqvCIXzhBLfH1QgwMqNG36N/Ni7JCyYE8Ur4uqO/NSqLFvI9jcG2Aa+JQniDPhf3BcxzgU6K
PuLXeC9QiF1eDAh3b+APj2VwZe5QMJLg1XKqmKLs50sAuW37PtbNS/M/M+6LLAz3V5mxZJR0Z14C
KzH24N23kD/h/C41Q2Cz3Sv8FXPWw4piCez2sSamuMCzJod5ubkHHbnSRlMZ3rhsflAcR23wsLEo
0d8Jzqr682JiRtT3yjp4PsZLRm6US7CW2g7+PwYVHFOxHkhKOFDEc6AeLOV1BLbq1D2luHn1kSPA
At986VTYrQ8XzbFFx5uQ4OvJJF171nYayemASzXtYz//dXtq9iHnilEZb8+66Uxv05GyxMsxSzH2
KEdqwe6YNj8wZ6M70YoY9fiBXaKxAKTgu3wPOxx4i6MCojUt0D42wgt+JAzoY2TuzEZDSQ6Ro/rD
/QcUpofcz9BaQV4gOwNCF+1jQsbqShqdCvHzQehTMa6bRG9+iyD7I9GBj0qt0g9t6x6iqMgyfHr0
6hjq+Fi0APSE+DaZPkQeUM3UWutE4cXAufd0IjG07+vx2Js7C//ZPOhD2S9cfMPeRqHUaJpfAXsf
ecJh4ZWtoQWyzlsDybZ5O56AMK3IynoZna3fBEaT7bGE6MB7ww6RZSm+h+VNTBPxYbtIxfBKWxL1
UC23XIO7wx2e8r+EJQ+sCCKbYxttX5qbkt9+dgHUhGGIGHxyX0Zb4zFlWOE/oHsvv5tG9jJ1cMFI
+I7hZOApC8sdde5wgG1UcZIwpasa0keMoAdf0y/hWQQgb2+h7ZOFV0sgZD56xbYgDN9bFI9FLffd
NuRyvYQX0+YcxcO7ViBSyGoUi15NnVNYLVEEckF71ZpiKvdUqsTGB3LNY9QFCIetwYrap1/DOo86
6Z3tG/HkacDkUXLnknbKIKUcxiIWDmwTb3M51t/y2SRuFArRicWw2MEAcFPgX4oCx4Xx0uCCYIzD
GrBckS56w+utxqUlkmHuIv5qu8jQn+jcg53ocEY9tLkvXq7e7zgtWh+4Zm5OZO86ioSPPpJ2+eWc
XKW4zWdJz+hGgw4LUYd3RoprH/qPbGElW9sfYDUsZHfAaBS+ovuSmj69uLgGaaM8tIj0zUCUNzIP
eCZ0BJWAtCF6pEUPExLNTNrl0yMVljajnJEgH7KrsvLfHumEcQ+YRDDcCVFSoOiWFvPPuyUoBez+
SXmv24RwJFcqoBCuyk7Ls5LZpfIQvXBmPipLT5iIRGmxsJi0JXDQ8DfAWdXaFfkwvisuRz1wtDdq
4Bza1qp5icHv5XrWkdabNZo48L6mBFLzU/sRh3e/MsBmbIL3bqRsSHlzCb0EvwLPKtNpe265fxPh
WZxW0CR9QWOVVtKbGKDupF7yu7ftJ/kKafBMaX99o1euq994hMR3LnIZ08okK+hjGSfOAfoEG7Kh
fupJjEBhngDNcPs7wATWsBwD8ccPdYqpQvo9/XMVQ8W1WJ6QN4+pzwKeyMMs0rpo1zNHWCe+6Tju
zuos7kWfCrY+JmQS9z2a7KCz6sd5g/ZlV1+ahmSeGPEPI6PDLka2jMPsklWgaDVzbNH0IkNTzDBC
Z392GNO32+sucVO/f1oH0D1YiGRGvmufumNtUVmVDk6J/umgCefehK7KDATMPqKKstC/HcKuC2zI
XHXGfaASFLQvOHVMTA7WVwXilkV/ybRFKYm2qsXz7xl6AflkGD6yMS3Uk9z2CP4UXYzCBVrF7dW4
2VCFfdxrZuJvbjIhTZ9MWjdKWKHsDziI3Aeo6nPCTg9rUz0Qcx5TSFRfcNu7iDx6cbXjHAXI0vO6
DHpHsFj5yo1dwCKpHBVzKXHUbLs+vyLQqL32aLz2zTQIhojqs41o39Rq2n7WGaqxUxKk19Y2d/0b
1BEMFh86T2Wgi1yMPKy6rcpmKEBD6QX6lSDs+jWQ/zASyRieaD9P1KM1C12QDh6dp7TmCBtI6qTw
r6bBSZMHts15rYbTqgoIwfnKNRHWsaSAMPNWW0HGsGPb57YUOJVjB889F+PfRHTLSzBYB7W7GY4H
JEaYiiKs04p1hQvdJbUVGcnnzb+XrjIeksJUYJnmZbO+F/RQY/qtU2XJmmGUx54LGX/85MeiA78A
VEVFM+TGLopyVNeB6IjMtV3Doo/GQsrKYhu9Dg+zRWIXeshT2mThZhpYYh1QtFUd1UACzrYvzIEc
quAsNUEM2bJO87M/JHnL8UieNvWxQAW6Wpyfziwpvj7LWd62CXeSuGEIvMf5o8zvS/9peEBexxmt
kpyO4nBJAMmOI9zacNg9oLjjA3S+a6OGyQHe2E8vNeIumlfreEngI9sIj92TLJVp81lpSY7GnEo1
khKUMz0CbzCEhdQSwdh5eJNJFFPxvjwyTMiJMcE5RLALIDFzHK9NB4WCjphAePrW4hD5MEK7ezyc
eLvBXI7ozNHGPPfLgHCSYXpP7qDuo4yUlRjXk35bqTXECZO7ysr0vZ8XVjlH1SuGfyZU2R08AHGr
EADQMin+1+CbX1azhQp/csvSfCuIJv7VpVQKmoLwKvMK2Z4ugoNaPCtIzDPKKAv2s8LHbUBpkDyY
pv1+Dl0d/qEMF+3bhuS6cc57Hb3Cfpj5faVrKQQNhDMl4r5RsnOa/5FuezDAs/6LOyFc5M0Tt7M3
1mW9I0RCm+0Nzhs8/YAEWs0wX+2ry2wc/TPo8wc2X5tsc3bqJ73TqDwxUcpq0ipudTmOc2lZajmX
xVkhunq+r11yTyylNUllYSJxwS4wsDUdisYyVGthpP7q3N9JeG6NZ7XfeDsue/6683MpLImTExf2
nDx5H+zlhayrhfIcfRlyV0lS5/9ZwK1EInB+s5XtM/LDYoJfruCmMMWZJQdwo6bPg01zxBpw06+R
/cmj1YVqUdmSEj25PYm3dqdYgawzHmcB/9cJOjtq6gHCNPk5JzFX3D5LIxQbmBWbUp6wOl5Axa+C
MOwSHlkX40dn5gHO430p8jg4tuWEls2i7WODLKslOJne0Oac9PTK358UXHZz4vWIxDtXBUwMRyjX
IDd8NRfOr2VQhs293XgfWlwfZEbK7ARzJtRG2TfoZ27EWsOoDJtFvaY/MB89ngC7tJU+hDV9TGg5
IxTO1K45kTuEmi+R+jbX3MA0vNCk0lxi+BpYRSQL2Y/dvlI724HaOz9EbZxFxXFvkIygLQ/0VyeN
6pDq+zc525ibFsiyqyyftLbNts7fo0yG7ulc7EYKRUhU5GzbaMLTXhM4i2znUVJSZri/5t7cyBv7
yxddrp0ooHAwyLnpMngA/5Fd/sCsmvf07Chkfk8MGxhwu3xMGtg4Jxx0VgFOApRJH6/VuwCvYn8v
2EBfQgacaC4K9tN7gjxcs6nDT1Effc6Ydmc08h3nIegA1jyQ6Q08jYpgR9ilGEtpg8H+byL+xjBs
y+BOwoz3FzWTFcajsC0Uu7Jfqpzn3aGXoABVpbfeCiwNkuf7qILtARUj1spB1inwoWhR7EaXu87m
+utiUjbSsiu6+BPKl7uq0F1eB8Hn9o2ai9IJ7M21MUqDDSSEXpj2f9CXW7ru6wp89ennCTs04oXb
dzCyG2SgvnnhEXS7BqFlGXr/bRWaqe/TAOydmUsZEQEjZn5ZP83mmjjRFdib1KhLAn8FeRaV726a
sQedbbmZVyXbPUPhEJq8uYXQxp+Ry6387ZBFmSnFwNmx3C8jM3ySBEkYF2GdX9B5v0l+YXwcSIon
yETdpnzvlbsNYBXiY3h+S/UDTPcV3e2V7QAJHKTMjjcox7NYaCPgY3kuBx4CTCA1huN/NEJS/3G1
12isZSgtRVeZgzptWyBV9Jzn0PELANtKjIiZRTAV/c/vZiSWwxFO/0D5RMtXT4rSMvEMgJdiRvxD
5ApRpHGShjMuIi33Z7dTbbWX1bEvz96BXkJJfpTsoLYCxZ5n9GLJinuaJMsyZac/0gJr/M8dYz3L
CJIgSiuduUD83uutELfsycgUcADH/AVhqTeSXSYe7258m1WMdIqb2DJBl/pqs3JqNzpgxJ1sy+T5
fbACyjvdoUkaweMk9PT/DNaJcfCKvi9RuwM6AUubdy2XOD4Z6KAKCUTFoPXxNG7EwV3Yv0oCJ1ke
2LX+kKQS+bm2f8HVYu3YAWGWSRHlbDIYObn09frNxXBdHAJgJWbvC712WRnW4uiVMUP5Ftdmy/XY
Lmc6NWVeQXBOnSUyzxq4k/tWFda9sZ9dsxncq5qxS2b9fJi7TwR8C+x8X7inJMByxpyAeP1zBETD
gprAzBParig1lr7AbxD+JSLowQhVkkm4DCDnn7O9C5gAKXwpsBw1Vf795qTpdk7ZLKc5Ng3/Cw6m
bIMpQE8zDkzLLsWSxACfRmDGMZbxBcVqjg0Y0bF7p1zIPTtT5THvE9sTIsFx82y1vfGA0ebjCwwp
0zuqChpT1XEdWBTAHSS1Oo4h/rMptQs24Cr158tEQIsqk5G/SYTCl5aop7ipGd0Qg7qfFbLYyo1U
dC3J/dyXdZ1yPEcFY4ngSQTh2u+8btBNKrpSEM2aAVaXriYEKw/V9doTAPGRMQDCx0WDXj/ukouE
TMdwibvvq59Wi67ZZoiprOD5tbks3hnxJrkLNCCM081f+DpzdH1ItajVZFKjvWaPVnkzHejtbgGd
nPfMwszT0+Y8L+NNruPeUBH0BOVk3BS7jXDjyr8luOe9xtQmUJqlHpVps+72tJHnMsoOVKOWLzBD
HbOl7FbDkynoWoTiLQrE3UGBsjJgIR6TcBau5u5oNJkIbbkAECM6x78MY9OVJPkLE661Xa3TC8lG
wv+stiopr8xZvLAOchpejgls1ieQ35+sSKVSOvI8Qb7pk7uLRtqkBaRQDib1r+6stCMyO/22OmUu
MJuhmn8SDUYq4yVH591iJstwPHSTsUH5O+WitVBM34K2iv+05kGdTribxBZrMiMt2P+chjw4T93F
FiK/eFXI1QgdCoH4A1vaDrD0+8mGrrBLFWq2IPzxjj3UTUPl0B5VHrK2biIYl6swPx7nz+CHxGcc
krU0UtpltNxgw8sOEdy2rGJnJ1ToFF7JTR0IhPa0pEdmstoK4oK0/LcY4yYc+IjryshsIDdvuqtq
jqFptnutM45oXPT7bgPw9Fhvt2KXBUkcTNm++s7hrE29lExmalJAWEgkIcHc0Vy9mQOZMSQMIXRU
rMIntyrqvKYKa0KhHlxJ2S+hFwGHfiUgeq5Y8by+EeRoUbUzngcmgiqZ0YOVGkRMLR2TYp9zV0ab
DM4iQATS685lmoCzj4M6g0eydX88DF5d9B4lnavJDgwU3VBQn0Jd/1qWlAA3cJXiyehrJkVhH19B
KyACtQn6UAfGZc/AHEC+qY/YPxHFl2GeLbC3amTSZTRMzR5oDr0U1u1Lh31LwOHmlQopMoJx5SBu
G1isSzhhdzhPGM6XfoBDah1DVJxMgP0PqobVUe9IDi0pg5vk1jR2uABN7PS7w5nx0MH9Xn9oAjAL
0TORmDYAu9KbiRSEQaqmkxNYQuWSeeddDGioHgBXNVkfmBCI+VLJ7lSPpr6U7xPXkAiQjWNBXUSz
QjytrdmzRp0Ss+RIHjxOVXGvoNcV3GYaCzcqrY02WUfOa7C+6mAiaY4G/DHy1SkkidOlU25s8pAE
qYoNPHhv1ou3NGRXdt4JRudTFisLoS+3QlQVeEWPO0FwuWq6QRfQoc/Kp7jWIsCgNzuxrPdXm+TT
NUzyW8gxMmikRYiJ9EZXTu1CUHuLEBL1FhKfsH+9298wIaYG96AdyKi2FAzo0MakXaeioIxO0P6K
L+4JA3MxbApyB3YEd3sHMf10hTZDFvkNym/VW7IqVq/Cc6f2QDArRJ81vKS9BUDJ6IsEf0funGzh
3HGRZSeM/vFZ8g8xosc1fMS4hvPyoUgAFjy+WWwM/g2ghsdg7uLiP3Db4L2BxnnkDAJYujAG6BFb
hc3/hwnwJSKbNLcsR2Kuixr6gvH4q0hgZt2iTri4sF68jGUWzRq4rfghYbak30uCinaaQlq4v8W1
oTQ01euHTZCMIIzixRcHn0zlkWLXEbweXxs3doSiDKgpGXBtwIIW7rDLDOALYZL1eJbgL8v4YHzS
lPQAcA0h1ceHucNKTECJIRZPyBQ4d7uC+02nLDpAaJPddMf6/uoCdqkWtWJWeuOy8U13tNMAzhub
0KSKgyV6Hz9avioPlZ2khNAJQQKurfjGS1tXWRQJ4E2BI9wPVeuAR2ajry1nGzIHKHCh83xvKDSv
0d32rRo47iq7UJcuSKsr0xQGjJgWBoxFkbN5LXVSiL/ZCc7c0Wch2VoCSG4E0DJflIrSMtN+/Wjt
nPbZ3/99vUyzEi0uH3oqLK4Ik8AuNbws6UD62fSndWcD7IJbWvpfNYQmkFI7i79XAEQ7yC2exIRW
2xCkXUCiprg+7k7TBOUHZiHjhWR9Ydq+PZk836OnE6QtHs7lV10yZQ+JbY3W3/6ab1uT0QhC6jgX
yrBbvRWGoNymUlwBXpx6Kitp+oNLX0fpn6sp5uDuKx3hxulx2UyaGB0oifhjl/mveWkvyGZdg4WR
fLB4uzoKtQ0+JFvIE5AHkGFWWIDTrqzs+4zmWpy5FcldrHraXka8jFDzM3O0eKnKcqa0RKFB65vN
DxRtOSjpjOE5/5ewrlEiyw/PDYw+PkjnRbgbRqbmuu+OpCx2MhCdTf9P+n+0xjJwdmfnZRRcxTQ9
I7Uem8oKNVbXdMe8mcni5afVvFMcLKMhgM1Gkwv2OwQfTsVcuJWrkdpg5GI5g2dZ+VZsJZyf4JeK
3tMFX7EOWdWTs/pv9TsSdc3Xs7dIL7roP0L03oRCRiYTntUYZDe7G4qUuGxi2mCMJUT5HmUIWEIN
MJ7Chpg5+i7Q3WSjGEbcAlIdGFG0xA9Sjm7/pqS7GL1IXJ1RoRMbsXnYJh2A7MI2ciAdrm9eBSxT
O6+8YIwQiITwPeGR05OdrKgKI8iqibuagCxXTezC6omHV5q92zaCkBt+ekjQI7uNAXHBkQQJdT4P
QNObMrJiDpyCGcl0Ik+pmDnJCuOPIKtWEDDBz6dWvPREmLHubdp/AD/cfLWk3v7H/oTXMjA5j9jo
BFCr/nDj2KRRnWaorYlCRsy3pTc9ksle81WTOWmMVf2xQ+r87MZ+gXO+E4Q+WwCCQve1TpCNWHee
UcSsoLJqFUcIgQvM3v1tr1uu8usRPXI8N41T803rR6qFFrsFbULl2Bj0kOHXDxxNt/eszlkswHi9
oyDcbGq5cKvfGd9G338J4fVYw6o24yryhLPkkD1vnc2tRX4Yv9OEgwQLBH1fF8CUzl7E9fMHAaNX
EiCCduSIlpFnarDpgZ6v22bA8SGAdM64Uq+0RzfsYLcWJzJjzy3308QM5i1aMs/U2DrLojKKx9dQ
VD2FQES1/T5V+0pAicPlXwIDVwSrwsSoyNsPCxGbdrsDH6z59bLl5aAHiF1YFJPDNVRJOPJKgqOH
PobLSXiYbMJr55UmQeGpAiUXQ9NUKCIO1Up+mzWAkrJnqMZRyyw/JsZSQO+rxwKnDyzmVDU6OQyM
6Q8hOIYqlAE8otruO8kMHT4GysG4JhSQxBg/LvyAO4JvfxS4t9Zn+UDCpn7436eyDTORE8J77OYT
BOTfZTkUSSjCmFUUBkglmO/y9gMgE+eFPh8oLb+LtmM8BXANOFe8H4A1xfEXnVStdcEoEdVDg3xV
4gcftQgdT+R5C3g1heeix0Zrr0UZqxGdp1kOH/YNF9wfgFj6XfkVlVIQX1Nir6hNLLtLbBNJ9hKR
YBqAUuestqpjE8b8ywz8tC3Ezm5O9MtsA82kDhckFa+Db1a40kLmSWu4LxAeNcNhWZYebhFDKG6z
JyriDFeSrCJdwdvDYtZChtLd0fhn23VjRGtjkBoOAC4dHzbBpyT/Kx2NfLIqT3iUWAthZ7UoVSMF
fMC5KfvO1gLcO/GbBP5egvWpolRbflB4tAf2T5VoQ8QUy3gRsJExkNOSvXdLzVal+MBDHYwHg7OB
3gohvrwVEOLSVIriHv5PSxqn475MCv+KsRzp0SEOxH4v9GyG6w+tVu9nVXEdeNfgg1vl668D5JKQ
JnDFUi4571kJyUSubeRhblnfVCKXRwBgMWY3UvDLVM/wtm3bfDV9Md2VZ+u/ocl+tgOpqD5O4YzM
cFSXy3Z41QlxURihaB8BeGVlQoezec4gyf7TM7VMnNo2TlQX5Adj3VuFWTgzVxxdg0H25F9gUj9y
3zwxpsYfqTQX0u/IDhmzPNjrJBYUuSbJYW4GCncaor3fnOAms2m4UVgB3/Jnwu2XLs8bRwb5cfkm
QUjgLMR9xAh0woe90wjLC/U9VScKpFSLicz3m1Or6DQUiXl7pSxvvTg1GVNi1138eXQXJ0LJnxss
84yZKD5uAUOugztoFkey/k9+/Cdn/9PVwQ60qC5zI2dKnJXjx0rONCXWq2QG9DWFak0ifuv/Zaur
+ZXeMmyu4vg/voODmpE2n7bWtUIM1+Wkzj91NNvJPLEMtywQRkUMJ+BKVHF8KX0OlHsNNaiwRYvZ
I1IoV1LiI536ZAfzAA3Miw37c6murqJYR74ZzJe0vw1RkaSIBxul8tVssLgRVb70VhU4huf2p+OD
Ff3RCavvmFYlku54+4WmtInx3rLsgfLzX9htSYj1L2lpdYG66bSQphrPNDeO6Jz/RCZk00W1S6q/
Zy1oWXXOZDU/D3nAjESKJiVJmzng54xcdFcFw4MVYLTccB/gxB4BwbG4eL6dVg/oo60xIXoJL+wK
bYCFKQE/8TZyVg3udS7+UEF9xADSt4nxkt70TlpiGaHRyQuXNoMnXoSZKcdyu2nv/dkjdspB8v9u
cwRE5NPx+l/CM16MTYUXl3K8YfXXjmDQVnx1iISwFqvGWa6Y1MhjmU1eB84Nin+UUYrwV8rIyGVB
VmJPlW4npaN28VcTUnDVU6/Ugdrb/egrsxrCRgLDDILnuEyNBed8RNVnoA7MnHksNbD8SM4yXzCJ
S0x6mCMuI2Wi27t3U/9WJ76JyHWi9binkc+mVvmKY765xOaVgSwWIg3bfMpyomjRpXha7ap0HdRO
/UCtGi2mfRDyYmmjnKtOsRbjincdhN3LK6gTHOmTXAZvLphloMEF0tKZRSXW4doiEvJ5X4RIr4Kn
lxLBQzY9Xuz8No5acRH4T0dMNR+ouWETi4gWN1h2oUVnIG/huoj1/PQ5GGsNhBveZn73GT2e6LmJ
FQkcwt4lphyEcqfTecUgIZBsH7XK75HQyfUfJWAQ1DQmJRUVPc4urkNhx1+Z2k+k8AQFolYHGKkW
uoByCmDUKDy8CgI/Fq9XykfriF4lwy92E2MG61hJse9+4iruRPscaMo4coHo2QjZIkQ2AvZGJ4GT
ij2JlnPhMpJwQKbJqA7jUn3Yxtz+9O8UfOVo++Ns5FIyd0HCOmPxPaQ7buEBwLJ9sa6ItBLdkzPg
b69x+BtzhlfFXuxg1gOURDg7oLghNIGkgEiETQEziEb6EDqdIbHJNGbkoEMfH61lzxldEXZPXv8g
hcGOdEsR46UB1owAv6K9OHD5wW+jlFqVEQN1HbmRqAJJmTUixFMT0M4GtSfcAGxhzb6rR34XvhIt
FS8wRU7Wn+JaJeJhcO1DzhQYaQ4ep9Wk+tm767AN/u4brsRhAcEWY+ZYEY3baMQf5J+OKC60nSxs
DOTeJxPg73Qy3+N/r1psshRxQBygnDSbMjMpXSVyOPLXSBuL/rT+tG4+COyuzHf5pDTAkIFKL3KB
k9VPSL7n2DJafnmO0ki/+6J3noMtz3/ee5QO6khkOyNirhAPmOv2FxhvolRs54utB3qJ7n0tBLXY
jPPCYG47O8R7OOOJI1JVe5pzTNBtmopzaaj2b/8taHQsG5qrsF4qxJ6RJaRK2uXOKNU9sH/YDsSH
fzDpzQC794fnwoxep1aJhEi6ayuXN27EFicburRrL8yCGCJlka+HLvUxRYMLwCj0iEzXf2+1eYWI
4ZuKRGCoEH9Za6O/7gykGds6otaG/mTeJwBQ6O1n6m2MbW+g29YmY8U8OuEfPrD9A0IGyZ475IT1
yFk639RWjZzmZoKa/jjOeT1Nm8Xh9jIvhJ7jLt7Jp+Sm0woar88mxueW7agqfJygTDB5tMnbq2Xh
E/TzeCfLT9R3ksmAukJZgqcgD1FNcLB8y1GtAu38QUBG/GSkJP3F1cikmzf+5xIRWbxtWEWUumJu
osTCqp6nTip8dNz40vsuLpk2S1yV658UxvcQF8SYBdCLmh6xJVO5ibnsUa46JOcOL1nvveyIIJ0K
IxCuZSHvu5JE9o2KgGACE5AEK+1PV5CX29cVJkrUymTOG6Eu1sIxME1og4tWVRY8gssBVpjM9+0j
XQx2w35InMzgYAPw/yzEQjCvfMS0d88btKlq7dD8UJ7fJdDk5LSx6uafx0+valgkAl3LffpZFlXk
NnJPP3g5+zAIHdtcBM28fvW757GoJAQuxf8UGkQhJsefplARxo82FH9BS5xXZH8UbaiazWMMsU3Y
iPnY/JlIYHYTUcWbPg+p5cRn+SUTUQu7YzL7aG7xClfMPjyx6414JTUfYYif+gxF12kHYSuDg0/v
sVW8RYD4GpG8i5WA8kD2UZ+RY7N0S6iQ/sGmeWpDP39ESpwk8W3p1qlHWc1lHpmPYCbpnie5nkUq
v9JPv9uLNQUDxMXKkYt41Ed0TKGOOqR049X5JV6yj4bgv5YXWSehKi33A1Dvf9SI5KdP+YKSyOjb
1ozb8AQAvLUvXntTb8+2axK9mYTJ6Xohsa/AfrmfOlBT6nfgrpoN6AF38QbqB7xWs+KIDAYRSKMG
yGetenyAoa+sppI0+bLZ1zOrwVWZRWzkeuyM6JiRqdKS0VQiWpfT65/M7g++lZ/gSSqK3fQjzwYe
0HfxPtLeNJ0TfM7UoolCO+rAgcxuTyfAMBmiJ2uOBDlQuEHxYIXgMhfYX+QZDTrHpXkIyqp9aypE
cRdhAG74pvTBfea9fVvcHAVrSpbhXF0Y3yB0SPqqDy3/pddDfUfUWzJ3i1Qbep+7ZMwZ1keDrOmN
PA906R3MNK7lH5Adt8wS7f+dm+nFhSyfaJOxaOaLrym/3bdx9P+XSzw9P/NS9QZoFgtoyU4iwMxT
deZVu2LAPPjuEi/RY+EXmJy8/PdT09wAyQx+FdFTMVsbMP7cTao2+1eZpDS+0gom09KjW1VRgDKx
JsZG/ZfGnRd9Hhdk2RC/1xa/N5csyx5LTPALKSho/GYwOA+WVpg0uQXToTbLnSsgjKPtjqUUTUbc
M2sr27Lr0cT7yQCv+0MysehW8uq9grA76IYCZdGGO9XORjdfE+LImYaICZquwWHufzEYFTEvCnZJ
KoWE7+jkQzPd0ypGStBbT/C6RhfLV1jmboeCn28wDK87h3fj0VuSmmpUmbuYmriK6d7B1MX4Gj3O
ivQYUdwZq0kwrJ9hwRMZvL7fHQcQDqRS+MbgA6NQNKHOPCC+U40b/u6Z6cJ8IQDdUcaFVoN0nb9v
4n+VScwK/4sFyzUolfodMirjM1Q452lUGaz/jnfaEZVrdPlBmCkwufNJX69f3rKVnTk/RfkRGb3H
bI8oq5X8trxJtVuWZzrE31EfIvwaZ8r/+/EGL4j5L4fUUD8WpJa47G0Z5soykBbCkAVgyZ6BCfFh
UAJo4zd+2LID1PXigj7HRMqQXVpBAG/dea0ROPXGs8xyWFqz9oYYyDBh3Bg1SR/bQX0VurTLHILP
8dMuJAwdSMqwFHJ+s/SWnnhWqEr34YQLD73Dh1CnqDNo0fiPY93MsqbUS1lpMX34KsSRR3uFRbWl
MAXSBxmDBJAP9veb1s7T6DXrDeoDzZiAWW4gHwTCeFGSNhXSRXu25LKikmTM9Mf8krpd4hpAaUSa
rgVQRAop5urQ1Iw+3PDGnX4+t/f5+pIpU29rY6S6kT9tW0/YPFl5pitn+IC1kLKQVq3d989kp6g0
p+NAYToX7IqsoQt9EccB0RKPJSf07aJPcR6O2YRWEpD+q37Piuaaz5/aba07z2wBlG4TIy33Ma8M
eGchueJdBo7C576xaawEKhmSf1xysVyjiOHW59LTgq+C/jYfduGjWSMs+ARQzDoIbwNnIj0h0/1U
NQ2yjN1Tbkz8FhdxhF9bX3+GSrtVo5KWvlE21s96Q8ePahsTisAXxeHPcWT/cOV4V/iFDu6G/UqY
IQ1YXfVEPdNxDq7JEwk9d1IYouUpwvkwqfzR6FGlonrPrDFKoZB+GrIsWhSTh70mcdb5h2yPysuP
P1SdkxLXq1Yz/8rTPpkwlhgXn+oBrlnSHrJAQzF0aO7hPHE9M0yboomdz4h+pH/hRsDrKnPE2NIS
wdNOGA7VkyXRtJEnDtWMH4wJ86aOJXdOCnUzntIS/3etOg972C62Qv4QrLZJ4jHRYhk9DTUwd/OT
Oe2t97CHeoDVTmqBkltmE/wrM4Z8FCGsx075Fnwu40hcuQnb9cVAtp9eAREUsVtkosFY3soaExPg
hds0MTP0Jz/RmQ5F3zIAzta0y7bgPzuNAuKmMz2XDSPo2nOsIcSTL4mwM7GNMXgevZ+wgZzlerrn
3YnmOLD984WZsHHTpswi6KV1i8iBNflmd38DVU4CLADKh55L77skf8eYZhtr2kfKT13okVJtRhe+
JyatqSjeL9+L9aJwfds1vLPolBD/tqR27yvrKLK741TQ0/KQUcEx76uCQ31GSzugfeOL69VyZhhy
GTvP87jGLAHMIaia9qe6mZW34SQHQ53F1sYxaA+GYm2XrTxvhzVK5Ltuinwl3Wk+fD6MGa2+kKZt
5aftitG1ow/4HJRvLvNU9O31cYCj1FQp2+3KlWciCZpvWRpYth8aTDvzmnm480yFnblBL/Y/HEUS
lm3tCtYNSnpX+S0IPN0kXWUDdlBgYYv8zO5P2L64nPfI7q25dt2Gcwrb8shKfCaBCOOwaaiNdiqX
NvSuAKGd9GVUCdW96tgeNvjTJHNxXyYLFw07LSK2BapsF1rqjhiBvv8A/LMU1Y19l65jWrUQG/HP
Q47GySshL2McNNOiRf9HnOZB8R2ejfJv2+ACMfTXJ8YIfPHb+f4yftFWIenV5180FijnX6NxsTd9
g18rsK90fvc+dZ+iPP1sFWd8zNKNbG0M72xPak+cMQFVTG2P+NBv+lJVe5q7a0NnNwQsWWzL9Vcf
AmzEidPWU2ST82MGxbUNRe9ULVuL34EA9UQNNBoDDPL/DZK4d3/72folTTgE+3Bmdac7w5Rsx812
NEYPzQcgpSuYhv9K4KorXqPVOhC+D196o9YQwoIJr1HOaR/zDiZlLdM3DKWGVFLlpa8sQ46VMNg8
4sEHx0tzPwn3/W2GjMGLRKH9/fZ23dVDgpJURC82okUQN5E0vi4ndE2ClgzQzhIQ3DOxolb2LjBG
X9xA6e/duXKNdHhlZXQFspE979WYj1UnoFuyMoLwS5j84HRPdYmlJMqToyXBdp+ObEEtgK5Bgyju
oF8ROtdk91csTRtkAl2SiWbtea/kJycnaJKAvmsS+7d+vykyZxPAv3CsQTE10b0pAP/hVAUFytIu
/WoBlPV409pabypliBacpW5IQ+WAL73m+I8g2TNfinjeTRtHn8jwcUWdaMx0zuWlVHw4rgamI9LM
dd6Ox8i4a8fED+qKil9/Zdj88/2Y31SGNbpCoBqg6gMb+zYH6dnyQ4+CZ+Xqj5LQs2+9IthZOjC0
h88MDdzDuQ1/j0xfN1xkzYPU9r9UsOSQx9oinRMEIhSdwzLeKvXJd/8Ev8OpYZPIOoh8JUNQIrm+
hvt1p0IeqkcRXUw9UuTNjIdUOWBt4BODGwoTuwqT529AwmdCjPX8bwss5rxEgmrvNtQBjYk7oi4Z
wNOM1D3Obyim22esVZhuZ6kOdQVIZBV9t5VZBIouT+WrZfj0zPnxZqw6bChPyJpoDtUMvV1mrYzM
yY5jaD/1SdVE9Seh7ilf6TOqrTDckIBRZYn7fbqOJ2E5KSpAFL8w/cqIJuwF92FIOmJvoG/QUfln
tvGoYHJ7p6plh05PaXNvnu82oblevBV4ftFWNJaEoXQ8QRcl4OS76jkbZmEWm+dvNWMU1wuiZI48
rZ1CdKXIEUDdJIezbqQXKS2qnjT4eeZ6XCXpwXhfk5fI3m1ZKapj6ff+/T+b02gtAl2Rd0ltyDlg
yIgxq/0PovHsGuBgt03UmmEYbJDLMMoghPDu6gJwzFkSHFOXofvaco828S11UoTvc2F1uHSTceez
lIhJddIllTpneUsEtzIVMfARkK60sN68579qnx64b7dZJqsgl+jqfUdEV8zmwDXE1On7CEZKm8qK
sxbxrKFPwLT+R8QhDr707ZYAvSw90PzakeGFWE6GIydrnIlvVqd17dOyKuDnuPXC09GvYm0rIEUl
P5Q3ba6S0Y5VIamsaqLY961n+p86chBtmEtlAEg6U9h+wy3JXe5pVUVfb6hFWMLS5zuoBEgWdTBB
LyS1ahPHSWMLiQzwBgMjPINL1VjKF282MKrTq3U1W0cgosWCNyNi++zQxpy1L1buU8c7X6kUjhBm
oDT6jXzZucUN5k2rzMzPbmXBbOiM+s30TLUbR4dgpJkzjC081w9cw48LObSIfzb1jO0pSO6GJLZU
4hGJtpdGMA92qFCsjlTOzZ5h/Pcdm3em9L4wKVEB4JWMoQAc6RxR5L4pcja08o0y83MdMwFU5Y78
dv6CnfAcTBA9/itvfzKJsOr4KPbVHPyWy2ZsVTcB86gq0CP1P0wR610husybG8ShDgm2GFVZ5eVR
oFQSaXR0Rc5lgGc2bIMHNEmMV+4+EUMfCUFM85eRymyJ+yx3yxbuBpQANOj1VnfZWdnJ88pDDh2K
QzS7fkKdeEM3RRruQxWBC6Quv7U71H0ezeLn80/EjGSDag7YBfjXIp+yqBZuypW201APebyWQKl0
FuaKkktn5KgaCJyGXZTwt6rg8D1vg7FilatNZVmWAkSjTNYrvElNo49IWgDM4xN0Dkk+eDX7qqAv
1ckuX7pBPLt9tq44hPyI/txO9D0yeDIIFCAjCpfXyzuOxTlyx3Jp/gymncAu7MIfixUgOilfguAj
24+iOWAqmnbkrGqQynqDx++mLhCy9D0uE2GjOcboK8hvFY01RnuAHQOj1c4o+SGKKc6dbIZ5Z2YL
MEuD5BD3tIjwEAK95Sa2V5krmmax7sK+0IcC3E1O+YCY6fJ9Y3W45+JpfdyNB9A5Awp6kItAGgF8
JzJnzEvtvxvXbHjyqBTzKJo6mOoO8up2oe5AIuTzZvm0adnrjBZ6Z+9Mjbz6HUhrvt+mbW0W2WKL
b+toecseOs+rGaL6t8J5e4nAVlySJxragoPz6s9+kf42JMFIAfTG2UmBIxf3BNubzt2Q3kcv3U67
TEcXdGKzDb/nbZD6ppa9HbwJIfIGsjIZ9lQrQUCHOy/JwLLqKMimg3HSJSfU9a70QjZxrphEPqqR
2ibkjVvgEhOX9a+X6LQW7Sc+/GLrP2PEyyEyveTEvPZ4KrJqr3tB1kx46PgStV24gWpHA+sXPLRI
MHe/f69eWJ7CtS8kqYtmwTfXZFq888xN+iLFGq2xZskyG0wKwV+cgrjgEDrIoQtaboV2KXzB5LQc
Id/yyoVku6IrIi7H50ayfYTZLhKmCySvUqD4yzA6AjZTfb6W3GzOUEbd5ppsw7K//X7vloIDjXxn
f4P4J50LXYrx0gF1Z4JrEN6NGgaOUvhXsEQmEr/thgZNqNWmxQ1mLR873bISfwuUdKN6W4jnZKrS
t5qiwQVdxl5z3I1gtCKLFmdshSXfwg2o18U3Erv+9Op1i6iWL87nLr3xxQyErZ0JAjFndJyvoHJc
AOusWuY6zNexO7nR5OekU7lQH87qIMMu474XIua4XPWprbdPl6UcFc9R6iGs7N3T09oj9Ql0n/VY
KOapFBpaC1vx2T5/wDaLeWQqIi1gcbW345/DRMmr57dKyaZNDlhAYrHkyVdJx6DKo3xPTnXwI5D4
Uu74btuUS4Xcn4juyWiWK/+5xESJuqa9r0fAca+EQ5sShGUFbLcbk0SolLFvyS0FJ+rKuwnxdB9Y
caqcQSW0LfvomQXINCiSRATNRR+eTdq+fc5NOBSxsR7A5JFtoR2zsIWLNpHLm6NkUbfZx+vHs1D3
dnuyNzWzhvI6yaz9+i8QcbGT+zQvpn7+v22RSHM2Sf20eEfXJQ6hFjgl52gmMK+0VfdjytPD1jR0
BB3KTDq5tpiM/HsKwr4cKu7rf6cfklS3Afir0Fb3Gayb5Ixi1DgzKWSq66TqV58IemALZRhuc1Br
eQPUBQRMlF2hBI7WqaGjirIa+IUfZ3Upk7QpvMK04zSe+GvNZUfiC1EYHqvh5fNxZOLiTaOtBgGc
t0XX196ideAT4kAAGQzkMgEkmFfMXIaCj3BD8/nlgfdy9JRKzZ3AnAodxd33YREdB6R1WFJqlUWX
D2DrA319rLaV9K3r3iq1au++ObPp4E5dgJRzh68jXAZcOJrDmpKY0maCMv06YlKzMAKlnNd9h1G0
1EsEMb4vilbBHoMg4ohEWlIreOa72n3y9TcIoXV1CgjVxOQ5LwtetGDCIfQR/P9zocx9xZSrdjaM
PT6KX3pDV8YZQF9W2RIORhw5xtmA+170aateSthQJSEERMnbFNc5TTu+Sl4cJjcuxRUjFv5oHNPi
oDA9zVBo5AB+Rr5n5DkxmT+4TFA/+WNjmuqfVu3DfMP8vi4eMm/htxZ20yHIWfa7UOzffJeH5xK6
CFFBzSvgkBFeyoQIIOAh2u61WUc8eBJ8EnARWUnkB8YkoCajcvtTVIsEIYOPJqXhAS2Oaneq4K/U
HbLvoQQpWLuVhxOSr/m1548X6uimFg7A8qOOK/Iq6bADEOlX/1TKmAGoJZ1MRgrHgnHFLUGbcWJc
9K/K4smOrL55MstACnYFpPV8ZJVbNrTfaHdkqMylJ9NODez40hNfcuiNggw2UCC+4MVuOKeA9ZKN
iqm4PTO2VCVCd46fE1BlZ5wyExlSI8M3WjIoewhL14Oo3Is8qKlnvcxPNF1KjZCE7PMCu6l+Am7a
WSCNPxn8tJLv8fP3ad2gfrfbSteyfGCJ0E1JlW9SBNcBEkuGkhdOUJ7zOi9N8wmCVIvLRbZh5I93
QcLykG5JrPv7ErUbFuHUnOnIp7Kgypqy06fAob+FzOgSLykDbmW7joLQAptN/lJvD9ssPnGCKPdq
sq4xKcZ7iamA3mVp9ZUG8Kz4JVLXqmF8eSSR7eV21MBlDjvwwBFzBwAxNowyRlOvb610k38c2bpJ
VJ2qv34TDKhXJMR8D9eakrjr4JuDLafYpqqCLgEmI5BgYLuQ+HjMk1cUjzGS5bMXz3y2TMHMr0Nr
6hArbJpI1NaNUkJfvG+nNhl2FoG6l/+XyJbw6I2aRaz3P+XlP5ElIirXeAeWPlgVczuO4fhZ8ICd
W6vNBGcAXpJ5nDjVrYWKksd72pKKzgBp4+wK5TnrCG1AZg549ZuPQlBpu28el1Y2dxZ7eSTIF4Kq
RaThaIMeo3j7sG08gtTgMQCaIAy7bop805oFhiWZaOU9bGu1+JwhREGigyXXQcTkuwewyLGZcO3s
aRRFGB4zR2vPqMHXeMrozATvHZCRMtJpRhJ6lGQv1wNuDwXTdLx7UvonUhi0Zs9b4ZyMgJsMOFYo
7MsgKrmSsIkAXZvITx6hBZkeLTaNuLwQLUv9tzlXCxCTiM9b7r1kvHVxC+BH7VEIVYTMBuQ8X/Aq
HuTHIGbQmk1QNchix0X84H82XddEAoEhbB1ZXNLDFzbUlBeVK0W27W5LpkwYPD3331sV/EJYBP2j
QKfWXOovd3xfh50oAImLaiVUUfDaHs7KQfoKV83iD7/vU5wKhOYvRJRRo66qoWLW5VfdEZ3NmmlI
/6FwfMNRYxIvhJpFd1Lj8BMi0OM51+DnrvurHPaFQNiEEQ6yrkHWdbakQfFAP5Q6nFSNCWtyVEvc
0Iv4DKTyHCKyINE4GAfAX7QGuD0X3I8gRg3WX2CK/kkXwb2PEbG+UVP7VO8a0ouNgjv1Ir0IpNFM
zmTxy1bTKmlHZBEbq8J/OYn5fydolaZ2cmc60N75REtQRKpcs4vmZcd88Kwc+DtJSH2OMPqj2VEY
Tg2J3oSGba9ZZ1e387ns7xj50GrpipB+3mVSIM9jejG0WyyqhYgah5kYyDJ5eUgmxa9cHYFwJiT+
2OOehvcI27ZHhLmozw4Hw6f0zIBOcZv7jJK9U5BAsycsM3C+qMxHyS4YGS6md2h3ISR7qDhSM9JK
qUUFVOujKw4JuUaKwIBO4eGVoqmyzC5WYA5F/ewhG4xF6ddUhCOn3M2vcpwNKYzPa14+XSb0Dq13
Hf78qp95bjo83ApxWShwSI840aKAj5HWcWdDrG7UqNQqzZQljhc2Q1qdFux64hrG31fsUsGE7xfo
dwbqDXDkLf0wSHb1Jm/znq8Gg5SOL31iy80cTk9eyvoB/qYUXthCQmEDrQJCo6r1c3CbQ0AIW4r9
eOBbOt2P+vYntwiwNH9p0xc3aB12OrcSJAfyF6T5zj2/av8Uo5fhjvL/MSozYZT4opp/zo1RYM9e
KOM4f9Kk1oZQ5cMRzzUxOZ4jI0OrTWJjCnA32dBL2vcpXtYjbTUF/JGRV08ylIGTgTKnYsLKYR5a
p/eJKdNEha4Nh86qzHMtAhqQf7tgGY0aGmXCZa4nu2ZFlPMrxV8fEk5Iji21bO1SQkF8doqoPLZY
e1uWdYy7qh81C7Y7VihXowMnYmNUHMQnrYVuFQkVLlwpTcEBmloGohx4hNtu93Ldozs9ZwkdlLph
H4jZYqzZZOrY6BaRDTvHegCWM9n3npYEzeDZeBwumwYRlJYNdcNo0sEX/K8M6i0o2PvsixCMATZ3
JsInDiuF1GcKVg1xo+Nq5v8VKIUef2dy1XPAL8vb91o7lRJUc6ysv9q6/re6taBY5AdRSL9VKaty
4c6LCTSrgT1M9D2vsAjG2eOEiO7lFXepu2ndSVAQESCLi+TEWNmlL09yXLHL/T6gQWOdFl5WRXjC
4Dm1G2pHQGlthiUSnsyolPO7PXAXHma5lPFRwNUsyuA07xhyXfx6igWxfZmeP/mZxZhvcTXvFMO8
C6bjbmkRLqpvYuNCKWe5srsPrOSoj13IcUHZapQftASUc6aeZV2XIdOSHEWTjSJnD9cmqqrSKFGl
xsSi+y9IBl/VxIdOg9bha+fJ8bH4S8YUdJRX2cofBK8vCSzpumeZojA447IZkaTLeJH08NhKOiBe
LtudtC6GqV9Uxn7jRdkMhliZnTDlL0Q1wtByBvpgZ6/RaBavDIfAL1r7SW6DYTN+DhF9sY46hs1I
Nh+/wnjT0zR+G1lm8qUWvSBbwNBDiiX7dpxqhUiDX2E3yTLonw/RBy3cvbHvLxo9eS775AC8V/9E
qNOgkCXKbXRF7LjOhY8XFyj2CmpVeAhGAMmzX/TinZOrY803m4ZfW0ack84d1GRqj6ubcFaKrHz6
dk1S7JG210dhWrZjQlmoisCAhUUpG4O85pduBvKRD4Xc3Eku4qGjVN6g5uQIsiYoUNDMJX+zNr+Q
Z/7PHTA2BXPGdNRV1EH29L0FV08IQ0oGzKfYbzaZZzrEWpdwR2I/IelKC5KijKq86RaOhrwinVcz
q6iHLJ+8+vvoGnovQq7AB5ylDuekXv/mGyh7sLfOXCEGNwIPGwH4j29fwRsQVF9TB5hoGKdDG/u9
MwXfER5dd1B4bN+0t9nga46MOzbvaVXkJS3PUPF+lYlby1Yl7P0uTtqzVBn9XR2RFE6I+Rg4TUqx
bvjjNWCAsZuUCv5Dx1V5q3rw3g43c4nJLbjPmTSKKwDQKacfNAP4LCXfyMRePX8x2ozuNzRexY/W
Ult8ufqFBZYKrlrZQRjhlbERPjRhLv4JpHpa9T2U5w4FZenEEUNZyItIhOeqUbw4VJGcJ12+ab0o
osG4GHPKPOOMu+gpxS5+QInQuUl/joCMwH2afnmc2C5HB3B/FdT4gUZc0Ax87pN9JxWToflvyHru
GEKjI2N1+rJRhq0nh6gbGFUkTx9qR8IQpWa8QtytJKJ8Bf2j2EmNoDtpoGLWbBMvmMFpWSJDNUY9
egEXS/s/+QV5G0ECyP7Ewp4yFp0/Zof3mwm3wgfHLO5SUVYQxPYLpvna6+COpy0s4mFXrbwahEgB
XYly4IVmf0VbsF/M2Jpe3zUx+Qpvxjd7OKzkNznRIxXtbXAKUNWzorHFi6tjhb8wYeVHX0IuO3pj
w5Gkd+Jds2ohqRDRvj7PgIFlZ8A+R4RgLpc9acU3qcqHS0RATpkgQ3zXNh02xkEa0JtKf5SjFyH3
XL1qS7Oxr4O8wsIUaAD8RaLHIg3hlcI7YvnyHyi4T/8/Ovf6ZMzV6GsG7jD3h3+4qF6pVkBeCudj
i3ixbrRq9/SxZTW0IyiaArbGR6tACLsF8HMxKS44JxXNbLSqd8dHCgtWKt/SHVWk+DpUci666sTd
N3dEU1xHSRPEdEwLpUmv9d4T3aoSBakFfup23GPzKgyRKJM084tHmROm2jvWkhfTSV3teNLwEECr
2dAcjQ+3y0AghQrcwtj/+B+FXxZGcZ7zOoi7twQ0acAWRvgbZsN6tbvq7gcVLR4yWBYBqupnRDAD
d713NR0C8bU6Y8iBn3D9oOf/qcohFxIQ1bJw9cv+1JAJWUj4o7wM7tQa+nVwUYcdDWJx8H7pFyS/
dkJ1y1gbkoOWp5WPT03YldbuEMZxuEG+Ga/wOheMz1iOvXDnIWh7ET4w6ne+7DrxzB7bHWtke9rA
DXsmfnTRh8YMsnOisqLQ4azmdpG75vRkiJEJxKHYx0XySbd83yqziLX4nwSe+gykdImLmTrNK5TR
W0bMOMTTuOyl/+vuoxSVfhODzKuPpf+gJaxq4lqcwbMyE9Yw93cGabGhcmVmRZxdGtx1/FJZ8/CI
2L0fA/GXOEFLIrLW3KaYeOSNNXUMDfu3fN4tgLwyxdRJxOt+iuWYkvAyGmAzdLY5ySGM4rGeLYp/
MFbhoti9w9d+w10Wb5QfCbjTPfsVOA8DXi/z3k9AeUvp/CwsIz1NiYCi883KHvcvxcy56guhGKeH
G9t0/6kQ5aspruY77oB8/8Yj3s5Y89V6N6Fc7xTlWFnyCgDppUweZHHTSFtCkYypwCuiDrIB3t9I
333lzbt0brUxMf20HbnXh7CgSIfdtW9Ps9xyd8W0nShR4iEl7heBbL36/2K3m5WB10FZZniJtP28
pR0eOSqQTkuNqBOSp3HfLiZ5+le28KXCnpkGaLrsaSl4XXX/Jd7Q1r55UXMLoia6PnmW5LjcwUh1
6gi2rcy0rkMOWg4Z2wT3Yyf8tDI5FhaonoHz0nVPI01QodTqNVisF2o2DB3lq/tBpd52ivAXnRQv
9dItJcH74vkpRo7YFq6kmb17dmr3dNhvUfqZMQWu82kY5Nw8SLXbZfx7nVfEo0+CfdhGF6jWB9ny
R378oV8hl+UTgbFu2QJBIDDxSqZhSzpF1Rsi9MQgLmZHd/eUmQblH7WcfrF5yceO6GnYg51spIS2
alloYUKTPbIJLnXNKtYN7PYTLVwrpwrC3eYK3xTilnnywj9rcIP4jzEcdIg5uzKvB9WEKWACJJt7
/qBx5oSsaLQeOAFkfqlt0FWzSn3/UR1YNbH48D2tijVo8FOPyRgwTBw74afgiZf4HvWASZrSAvWz
tx/593yadOt/sDYCZrHJfhUDaURQfn57WyMYdUes27ZkHIDf7f28QtbSrsw8/TeJn0+YwCCSEBer
sA3Pj2CGiaraH7ySZzyO9znf+JFXb+1jVxJ7xku6Gd9xZKnDaydxVVYWE+hYDdWb6H+Rlu59pQhv
x7W1NrT9NK2vo5Z9gu2golFUv+gq0QTsE536l5c4IJE4cmqB2dyk4YERp1EIlLg3EaSCi2o1WVzP
we9SoU8b7uQsqRcdV7Pu7avgNx0ffItLGZ6eL9pGS3qEh0ycRf1iVIUnGSUEHMsyh13q1PIXPPy+
gN3fFL+o9sLDIL5AU6OCAJ1wJwhF2YflU4Vv4bwC5Z8RYMBFlckFy7AYpD0JO3lBd0EnNtuytpdV
WC6IybVDT+i+SVNUoeMyrPBGkTzXCiN/HPVnI3iBO4MguR9XAuYgFQtX3ohMroDCCWB8fCB6Xshk
4kgU01GPlxMNVb7vHtUXtrRxNAi9X3rCgYhYCIxC02J3Y+lhjwz6LpEeF47Gn4B9uGUduC7DQiCI
78O/DTk+ne7y14rYrF36WYIYLLLjzelMGVki5+TFL3D33HJJT3AEH99FFFUKEjI75FzDY+pcK8D3
uSL3h8N0TcaMlMCwUzrF/5Qo2v6Hw9iXvCs39GH7Er4inhppge7OODvcOyvED3O2zVDSrI27De/q
r89EYjUIkujsdlxxg0QVZ8gXbAUMRA/Vv+LNYdVn9sTEpdWqbKs0zWE+Rcq463gJr7QgLG+6Si9C
IfV8y9dAGPYscpOhYTfJoaZkW2ZVAxTn8TZpCjYYat4V/NU8xf4mTe+M1LddPdtyiNsvrG7SqiqS
Yyi4o5iVaYC2BkU1KO5Z/rOB7KZLkb+kOACos7reanU3p1YK5GtugSfjridBsSVztDiw9ug6nMiJ
xPcCcfU0QFsjSf6m/pgXJE6v94K7yp1seqQNV6i0ONuX+kWe+JuAPRbNn/MtzsQRUvmA6HECAKLi
sRJwLa6tBwjIR99Rp9uusmUb+SOJf6+bq5CdAOeU38gOL2U7jTGuLRpQxH3UCrgE32rN91uPfiLv
a0HiiFczh8iKyiZrIppT6Cai5n3U5HQ5W+Gn3rLhR8fuqm5Xho0sGWBcOe/8U1gvU8JerRq0tfwU
rtYhAy9nwfjc45oUldFZJgN9W0+HvPt2wi3ZZ6hJPike1ZM7jOY86IsnetdrGaI5bAu3NRKQoG6W
nBslIp0Njy1g/DcB2egc/vgjP0NyN60FCFO0ymTM6Ia/XyFqc8S7iWPxlYWrisovR/vE/3YYdQoD
R9Cs3miTGdxXgadb33xLSnvjyw3UGqq6RDMPP0Q95nhrjP3o5BBnZjxdTJkYuhPudXAdwQwoGMCL
6YPCK4yY1ZmpiPX7D2T8+jTbrW9FvBztFH40W8rWbpzzzml1gfvDqAORcgNF5pXIL0s2lcl6bzUy
w9xddoO6ql8R0E6kRUGAhAKWFxUI2JKHcoyWFyGytpZmBuugrHbXsvIo8Lcz14ayjhdYWpaJ3FWX
pHrf+scdoPC+kND26x8tq9mqO16SojM8oAexmWIXkkNWIzrRFsYX6z7SiiPPv29b4ez4UA7yPMVW
ndChMa43v6l5zq9r2sqVGYSs3SptBs2jAboEwIGcKdF4RgO9oMLfuuSFXNkOApfO1Hdx8Xic/H6+
Rrg0vS3Mprb9EO/70vk3IRIivwdADSYDOD1noj90yS/fv4oTQrndrukwUYqHVeG2+N17+ZUD+gq+
9fSNPeqid8wXKKYFR+ov5ej6z1Sieixd2FhkQbSKFuUpq5Ej13ELN5BykHsbi2K1pB6qUHd7cM4j
Nl0E200hjtWlxmlCk1ta6LwvemP/OKD6S/rymfeN+SP3tNQtHYKN9cMA9WBPDG2+CTB/JyD5cq+r
cFPDRp7NIg8n+Xtv5QEm/avymYHkO7nGducJNf2YYHHIX3kJlIqE7x/xlGdS05XJLvfcZHTKDzsJ
EiCzYifUEfwlVKxVXpL88RiQqk0i+yuACv5vqzBS2JtfTqYWt6rtQALXiCOZ8UBu16eKHiRwSiN1
ppMCcdnfDAaixm40nUs9CETtGBeRB84G0462TRYcC5D/gvBq/k/LqvSY65w3X5YgQtq7km+AnLRe
LLCnQP7aB1uTQxPIJkPPYR3LzEQqhS+0LaoJP0LH1JLhq3JRnvuaQ9fKkuYX4xcflNRVOnT8ZZb3
SxiI0WhMQ0Dm5smB/XoiAoVHdeyUiOj/mEPBlFOgmv9yL4QL0bAJPZvjvmLFLlSIglDk8Yp4WVvc
ATR7aNOR7E6N5vFADi6UcT8YKYM3ZZ36eC3kWUvFSs1d/CUkWg4VxA8uLxyQJQPOVQpPNqIhUyIo
aP13aLZGYqWC58CULP6164jk0vqadkuby4m4ZURiPS0mOzTLERfxSuZqaEF31OoBcAfz5XcfFlvh
cCTW6Jw7qpRFXwirsEzBLyBZj82Xsjo1e/AeMpFy87+jDPweq/1h1NI8WJieL/rNyForgbA4npfS
eVoSYp6vk6FdckNpM3qKSV1FWST3kmr/RXN5kK9sudPLlvn5Pit0PWnsXN3ceePDeEMbC2P2V0LT
5Uh1Fe+OqMm6zexYCiOUZyPxCm56KuG6m6HOVmkmru29PzAcyjVmkbONhR0plKNrpgLQlRXkYjrq
O7w6LhnQsS1H1qggusR9WDv0xE5jJ/J+62f3sAFM1CCDAuF8x0ytUPnvNt9Hs+Z1349WOa/Zs6f+
SCO5qEkv4ZhVwFLORKveUbymvAYpt6qTL5DESG+70yVW6e6dbtApgDhMfM6ahK/KmXf5B+m0UgLe
M81v4q2O0Fc+6Y/BClJtYGbq/cS0qGxFpwvKOLNanU6FSMkR352+92DMeeltvSocUE/oA8adbcda
5ssuYqwWzZWdsAIPxnnc5dbH2ws+PO4l8afJW9gDfRdHd4c/uHQQd5V2JS/A7QHjF5LsNEQkv4+S
j2tGX0TAybIZgaYN1hIMU98lUKBvjVm+NV3ncpll0k4kRd4pL5Zy//jYDYAN2VfYGFXMtKBI9SJY
LTLO8Um9g99IKo4m0YdqUqx68wLRzcsHNuY+hIjCTSnkDxLko4d7Rvg+dSibUD4HN08ht4NWUQ/+
WTSqQ5MSwSbanMNfiDj/vm1KKF1Ilrgv8mGRm6X2P4V8QvVsNEO8duh1NVf5+lx/t3uOfiu41dHx
1bg2Llpjey2R+UIeDc19x0o9XBhte+eKCkqM5tjgxGfMYJ8RUEHZknUrBneiKMASTT5e++EgU+zf
66+G4Emrt2av7FxajYbSBumuVAa5BwwppKH30R88DTCPzatgRKgg5RMlR8wnUaBw004I8tA9XBsD
jrCdz6M/ERh8kAOiJXziH6NEsxb38s3oUKPhz6VlC/5UcTFHAAqHTDFBV0GLM1qVLCkqMwzot2TE
mCIhdP6n0Dv7899bo2e+eds9Z57dd5mykrmqFnNBXZWl/+i0p01Ct+Kl7sUo945wHfvWvQE1OB1J
kwvf5ztOOPcB6T9zpQXRvk8DLeBFM39mlWt1BLzIG0wTnY8dnAAHkwLxGeGgTBlAr4HgF/8aZCbP
VNv7ex/hT5mHZ01xGKsbbw43ewXzdstEShT+88XgtGUawq6/DAxXn9UGmW8ZcqEIk3h9Gru6LzGh
vXMtZcYDnCWzxnpwMplheZ+g9O0ELmfPQxvWc317GtGAerlAPyn2c9BKtmiS07XAZT8VqtBlRLkv
ztPp/fVcF0h6kzmw/9lm3hqmPmve2M6bNUZBz9WtWrwJJfxJFNJXazX5oPXqkbWCtlG3SIXnjMb1
evJnP/WeJI3WtQ4WKsbiIxX9lBypYL+tHkmPQdbnS2Sprr2T/6bv5+n90NCvCU3yLBILvZLk2jQW
U1U7TC9dvhRvJd/C/C5f0whxhNBQlERgBoZNEmIAbBA0ZDKu6T0byzsnG/pRtbBTOvKR8UlF6bZB
D9s4/qe9RcVhepvmrS4uWkKMakGU2krzOUZvyvgmRtU40qVKAyxBL6EKXrneBUh8DbcyK92c57PS
DvOCzO7vLicEp94lOVYKOQ2QvCpoF0uehZKqLVErmc2GuYtLLdNpzHTjJYEAmEarY2MMQ9aAcI+q
mYwH9YhAs3mHT3P+G0MiLKgiP7Yakf14x9Qp+RYe+lcyzz6Mop4rLhIjxzsu0EVD3NdwgjyxfJlb
o5JBk8TVnLDfuCfFcUKSVESrRNBwhAvKu8Vg93mJiQ2yv/obUvFijhauokcAhSAIy+kucMOLm/Kx
aIQme/zY9MFH6lXyHjUltHanTjpydhlApcy0awi37IX3O7l97utQ/uW4TM9KcR8HgQbelwA91Uz9
827qJBDQzpyhzItko+vSswfNd/7o+/Wf4ayaxSldtsSTVRmNVpizgJiIWQ4A+QuUDHB233gRalZI
PA8tGC7lM2duM83qn5rjrsyK48/+jDFpTuP7uaVnL174C8t7E1DH5Qd5w4niUG1bdKbcF/oEEMEY
xBPn94pLA/GlgkuBDdvUxEk0Jeq2rLNiCI+mZIRDxm2uUe6eKJa+4EjhS+qV1KkxwXCaJIe+M6X2
H4OfunAHzdCvkahglqCPJa0tp+l6Qfb/KxQGnAZRKTSgAZGeqnaYWLXfiBQ9lCkK3jU1wHvgXr9n
/fN0cDK1zjLrRmcctgb0n9ph7hx7lvRF2XxSk6h2gjyMuXcu5d+cpdtjC/ddFfqwbasA0b0Gko9s
eWLEED67Qq+ruvhTv10eEY+pIQlbPwcffORn9u6II4pwJ9hkbJO7PkD9vlzLAxPTku6/cL/yJtxB
Fmuk+bBpVKz8PYVzkJvVAWlVaCpubxsIfHRsnsPKwsch+ZOX3GEYQku+UzWU2u+6qIRr6dYIcIYU
B4+z7+04IzDlvgRizEORGtXcLeAU0GrauGAAkKw8uYbJ3uZ7EaA/Wc1RG4CceSW7Xj8Edja6vTm4
a6GAJf6x+d201WSI5p/xWEgi9qt3VYnDezXosX00nSO9Vvf8NcWB8nNabVVfQwPOwqj3r5/K6OYi
ZWOF5LAbIUOylzmnyYEvMezIarWdUfUYhzgvmv/GW2xztNy01WkJmJjvIiDV9vxSx7pIfsoKlv39
TS7Fk5OlVyB5nz3ZNFUzOzs6xrkOufA1XRJD0kroZchPgZEe8Dwnz5S6iZ4dLMveO1Ma9MjWnS5h
YEtvsxQ6EiTx61h1vIHvJ4+Hg4A7NGYjhlYblNO874YLobX4JiR8LJ8StYh3sH48ZuZ2/ul0jaI7
uDFiVqUkKUPV97/mS/KOUKs4YveN+oJK3fGyC80vdF2hoe1UUqm/+eI8Eq3WhGBT2q0pXgooT6Xv
yySTXDv1mwCMB/PWwMzjeHL11TQ/9kvrsu89/sqoz155ZrCtF4cXNfu1Mg5XN8PW+d4wVIHa+ZWl
5NUP2KoT6QGioh0YCdvoDW2jMad99U/stlh5VUVVX0TgCOVQUwlYz87vlnXIj3WtGfJADKJNaxkL
YjCGDXdAb7faftO1x+bSIIP1EgSMNxD7/Sx3IEyQ52IF0pliMUFc24t+/Ptbi8ldFdhZ1JS9QksP
g0Msg/QXXoyecch2h/Xr/ciK5MpzhYmcdnCkTI56xD0szoZjB+0SosSfYa3C98Po0NKQGEfw6BPA
O8pLGQVum3Ao6xHgJynlkJ56K5qw3yo6zljrmycFMngZcBDQ+mxGtgTtoLiDzd4HDRXaiVt5JFFs
yjwOelgojPhbk2CnIZ1Nz0VXvrkHJ4WZoh2CnCEs+hiNOzlLPQsWvwwcFx11Up5ppTeh9FgW9wMs
UnXJm6zUOSRBGV5/mXLj7hBwVuBpdra9ZgNTUCaGBvnYS1hTUOQKnnVd4f1G+qt+wTraaNIqEFoS
d6ZTeN/vJelH4ZTCpDR53FbEf+I3W3Y+5wrXkxP2rZJStMANVg42yGtBbhkQILoZF5qweuJPwI0X
Z6WATKpJco+U3RMds1cMsxxI958dm9Yuy57SdZHOq2SGscNKnK9KmuP1FLG2XhOwr0jqeighG5FT
BreIy/g6yWvkwY+CKW6UGMG5iBnR5gbBX0FBRTeuQgkMFsT+vXUm7iaJdtX90CEnWNviybAGgHtl
GQx/aEBpdROCU4UqCpl3xuvqYJshdvoCzDRE0TznEI4DW0WjBaY/No0Z5VrgFm9D/YxLN4pnTgqu
5E6m/jQp9xmCAxczD/cyp0X3JCO8898iV8A3BTieKR5eeteUjNSv3lqhT+LjbLrAqrCryjj+KQ/L
yVFWBXpdyyLWCiaPsDRgF0mJgXAJNQ1oNd+bOW4+oI0LBxy3eqfn05/89eotN1qCWxP2XYTynH5d
eBgoGs9xOoKUgXsO/A4eHNtR01qTdKtbm4QGDc8s3fkWY3o5gyolpdJVafuRY9smrOxpXD8TE82D
ijkv4UKBjGbW/EH+TpnMkCXJVnCyNIb/tNpzpz1O0XZcngCtTWMYY0jaDQi6cY+wavMn6mCPaVTh
+RlSrye8V774UiEBl2nxlNsiErI8wytPJk+omzyAiypevKGTKhb4uMEXwjVqGcXYhAWiHIsjG/Hf
hXjAkX6b9a0QOCw3vCdSDRprBrd5XVss9hl818hcJAA0+RwddisUkXzRg5bTlVyEcA1+78gNRpqf
Jv+QuLp2mlgBEOmQgF1tSE2Z5GwKTjxCJhyrV0d+G9DZq3pZbIAVOen5Mk47QJ8X9jFLq2xHJpFR
ee4vXR4FCqAK7/yFTu3OorzEn3HaEiklbrkjDdEGz2DkBc4IIeHQX4GnXpEFyTwrc/RCdQblgUw1
+Ov19IXT+RC3JLH8Ke8QKR6UBNnVPiShIlS5vpzdyqOkjzghiL7nNYELZ4hJb+KZifxRacEaQ4tn
z6xDMQ1xd7AkqTs9O+X3REOyri9nXJF1fwaDKnfP9RW7NvQvC6nl82y1RYVg++Hal9EV0xN06+lc
RQx6Ga8453S9BtHca6+rJ8b85PVS37mp9+S91VbvlpgOSrui4bstQsLqxfS3QA40ahb5jNJ/BioD
6JdAKP1IP7aSTky+zflo8HQDBGwzpFHeXD8iBsaHHO+IIJlb4ROewjQnOrSq1DdtEk7DHMoNvEBn
lVMKRbwfvZQSu0sDC13+X0R1FrFiKZT0my+ZoxRmA1LiC26kwZWPUcoKqfTSe9hbQad1MzuSik39
DXfuxZIxDvwLACFduhqVRNCiUjYHnvDOIrUgXSUCQHleRycowT+c3qGEpJAbOT20l4sh3Ag7CCbp
EucxZLlYkuq68qCS6p8R6tj1UrB1KKeESATds9I7+RTFXsNQWX6Lm/gx3N29v0CjhJLNBA1X+LBy
s6AVgCMtXvcQBZ0Oz7Ng8BhbS3anr2Rt48wX6YNO+w1WvvH3ZyVeKZHj9Bm/4ts0HDblp82S4z8x
dCZC8Ud7zKM1pmFhd+ru8lL3i89JbkH5nxUSMM9LmflhLVqHUtq7ySQqDs6POPsR0LAL6LlJiMIq
rELG+1sU5pe1faXPBWEL/XPBEMleD+m6sOgOw6HvBRcmQv1gkEWf/lFLMF26lt+8YuBUFgKVQEQa
sqNPZMNnUgKAEM/7hOs7d/69AQgoEsxkxWVYVVn0pSiXBW6o8PWJm4oEH3AxlinbgsRppDahookj
X24Cfnywyl1yfUsCmw+DFc/GAFloZUObdv4v5KtIvDQF4yxdvFxRJUkHQFZW0tFEKncj7W7CCL9Y
ZYHJr/E6HxFSKI9MID4VG/LicH/6rvkteENAauekMbEpYQHNNTYQKhoQUdjyUq7+j+QFS53jpdh0
2T46XNgPOkoL57XWML6jJVO8/dSFIlbR3ARSCuSWvr6BIEdqIrLrqJs+s3DJJfQ8++A96Jop5UIV
cj2tM5/UAE9L77/Aw8ffOFnqApwD9HhWt4VbzRkj2e1QI4skTUsSf+dqVMraFj1hz2MwHUhIzqUR
FdJiPTe2Ngev98MFCEMMHxvuRbrn75dv4eaEE1knYOWfO8vh5ojoI7CaFyeMD9qhsFQWeHlRr2Yc
85CxmQ4wk/QpItyyiVdM48QSyKTzXT93FrZHHd+MyEwyEcSt6CNH+FA/pqihktEkjnEZ/t9XaVR6
yJZnosLXbQ/xuOQtNx5mDKZvRexlxMn7h96v5V5OWGG8Zv6NJVZpB3wXD6AHsFaBofg5HnucEzZB
R+C7HOjK+75gpvLzq16yB7DJTYtYqANiZFmXYwo8yvJxcErQBo+IilmyAt0gYUacWFp2Dln7z7PH
iqLn/vij/h/4UKBa45xOfjpzfEHHqJ0TuPmdXrYFzXc/0RzgZoTUeNgZtC/EA5eqfZQAhlBKup0d
sOXQ3MGorivs19sOo1TgDe8h2nuYEhW4vOfY/bP1JSMXKVMTFOugyCqZX5VOrCYCjfX086R5Ycht
DI9xph+TgK4yb13VVYF/caFThASoY/Y45yB0gHLHivzXtka5vlMOryz17Xr1IxuXJhBDU4ND15hW
+CbmRIJ8uKRK2+A3iq4X9V7Zq69OkhcLATw40lilL3fvLvli+ByuQy02bZu7djnFlKa4bPuUE1OZ
6gVquXzE9l98hA3BcgpEDrNQ8u9hJ0NEB1ld+czhKUfV6fjd1VcFnKpy1ajvjMC8ugJgqsgLb7vy
cO3ul1zLlOBQT4iUHJfxjKkNRArnT7pXgs2HwO8vvb1LDDk3vrPx1MJFVjUAyL6aXq9d+Ub9/iky
bqDSFGM2DKt57VB2071UI5jIz+R3mZCsgj8JIlTZVnDgdXVNhA4X2UCbljlvUnoBHuBLU7J+lmM0
EtLPu9GsDXVh2Sg1K+k84oyX0kJjpsqSRS4tCfkETLO5DR52R9iWkWhua9UPtuQLBH+PwaO8gccr
wLKCDKfFoxNzwR66kKHBTnNbLNfoQm2zEtDkZSppeX4KzGFW5V0NTatwnYtlKfDMQ9kLHahkyJmz
UxkUX6PTGBi8cI0dr4MJd+LlR6WjyDG73D8Q/A1OJW2Efbk4Nwnahoojwf40gkh2VnMQa+DCySTo
M+soX22/9tiTOWT7H6nqf4oJ++LfO+axvnm1V6BBMtx1qwHlFAx1hpFBy7103x8K+/qeU8rIzwpw
G9sFiI9Kd7s3AC2xrUpUMlPI5qhzJZXYFPROw9sIrPWNnPlRfUVhgF7eXl8AiUx4DcWlL1BVTodf
KfeBnFn8ERwDpoD/CDUvtKr8ZFLv5hNHhayUHitrmKhtCfDn634Kp+7RVi4fXoH2q5Uk89911qXB
AIDecsgEkFo/nwClKBI16A4C5Wu9NAUBwOuh0MQbccFPC1oRWfJmfCaKTFTK9EpFthivqrwvMNiE
LCeuBY7/Bq/2XMd7O+Gt1qFU7G9Llkd95QFWdu47A1yOnzEOY7G4fUdJnCqkjgZVQnsKgDASnnG9
Psu70pH0l390WIWAqsHBnlDaE6vj5l2uv84xnnTc4vmgREd2SOpAWTcLqGJewG+I8pbCdWKnuTu9
iD/JZcDJudy889dnefYnfvv73Td7krMxHXH7m9l2yH/zfKk0CxCZszCCKfXFhkktyjCyDWjjkU+F
BOP9abDPHgGsG4tBQcfwvaFVNqvSpoB9m9GN1uazSu7WVZjw+XkRjf7Lt0IMWZpsKoml9CzJ0rFx
3Vryfv51Y8u37rnhzmFUCEZlqw4ANWGQd6pAG5Rov0ecDdqnGwdsrj2FgN1tkBShzMsof6rWGS1e
jfff2iR9d+PyLa4zRQID04IThNZTIXlxaXsjSGfVs7FY5c0VBbSdG2O+y71mjy37aIGvvSLi9zUW
GhkTEMiWlmC4LgVHg7D7yQbfPtXlFa9LWB+8NIx6VJCvmp0HPeJSD/ic3iohezOGx+CP5ecL3t+M
rNHD3zdRKx5spaFugdl4TJnDDgGm6RJWi1q8MSN7/YPnjPEEyWOqwI27fRsg6PUCKRB2qGfARluP
ZN6ATiJqOsuGh/S3jCAigRwB3DftMBx8KqrXXNKizVxB1TLvc3qD9oDlx1IlU08nc7gjjaI0GOXN
bcIgqDnJQ1PTT/esdXm91GIfUPvZjDG0iU2N4mBZaNCTJ8+H9tYQBh/5STY1lnO6A324QJxNHdNa
9sGdLtVJl9aZqW9HkVxzTGzy+jd2OexeukQPEnXHjN2mcec3VS3kNiQOiXpfo0S1HEDTecy2d31B
fl/qW6iTAwzDJZr2MJ/sf2geWaT3WKNCXDS8jFKs5jsaSMND+G/9IsPlYBkspqWuoAkgQfhnecv7
pbGC11vx6HJlpZrWBgmsqS3iPKkQcToTrdZr25XV0s5IXbaigiD8DiLjI/WpNRbiCiDDxfl0IiuR
qVwsMHVoVJizK5/5B5qnhwZ6AnmvBhf0ESSign1j2FHf5+0bdAArujh3iEVM14TQY0RoWLBavDw7
9nDGplIaZN6mY0Fh3SMeSwCiov3QYUh9MTQ2UGAlK34T68gvVy82fXsl2DBcRz05IEs+ukNOPHjP
/RG2ivH5oBDqnBYpmnFaZbTvN8QMSnCs0YFUo32pIKqk7JUS/Mu6zrrSxjJKwIb/q3z47wmZJszN
IHKvgfK0oBYQYONyPChInjVw/jK1Wxm8jqQvPjv1yi2H0+RxFaEJKZxxkzEuHmAIwk48VrYEPnmt
tyidKKEO7su9U5VihtQF2VDV6F9p8vpGBO3PA8hzz1EaIWPIrTwhDQlAFiYK+z+fxutdFWNRTXqZ
6m1RjFQVdHo+5i6fggV4aZb8DeYDnmQ9/Q6jgA/7r+czlTtGA4g7rY5ogVXK6wVRmak1MU74V8BD
qyUxZ2VPOem2IVdLHuZOHK3CPFtc700H8ddYIuN422eLp+xf2zeA5h5pIVE0GUn1fCpa5x6s1Y5V
csimh2EYUrmgQyh/Fwlp5OHFl/eS+RNfXVPup9WLlSlK95MQhJv2w6rYsuFELm40PAbBxuqoAseX
kZLmgfriygO4uDmTPLPrW9IkN/SZ8l0Mu6vkVIPZFx2oQM8OcFrp3FVy6rIFgkxKxbkDCcwDLO81
xn57gx/gCr+OR9kfkoylzz/ZO8uLMGNnUzQSRXnPUG7tknSQhygSUqkbr8EDb/3+UNCqqRyaBGBx
aQA5Nf4ubJFWc9wYYJwpl+voRUiYR0aab6Uxftr7S3IIYXGXz/qjVr93UghPQqSeT3cOdbcIg5Yb
Fm+YysXRFU0wNhqvKuxYrQL5j2qsIe3Twoz0Dp7s1RYbsRBN2Ophj+bzTDo6G7bwGpTWF+BQX0Cy
d0N06YbgMaonAB8VLecClBeuB7ITbhwtI3q/6YL49aRWXQKvo+sxrnuy/yFBQxRfH0Z5DSrvbhhG
aT3jwUBcBFNOxWLjIx+WdGKGnG3EThoOcfdbymy4rsz7szMawOa11Lu9PSZXQMSZ5uN8eOx217z8
LHvgNRLejl5TkJPgX3KUzLVYIQLWZDyM2EeQdKRZeRwSGz6c3xgl4mOHNgEb2trjw5idbGCX2cRY
tpNyXNWJi8wgRhUYNlazQdefg6LMX5dVNm0TSNm1AWItNBPN+kRF09y7JyzWhnizUyv5WGq6kLcS
YbfUmxNLGUBe4c7QrrFW5OsfPtH4Yu5QnA+s1CyFqcE+fHZIBmB6WPkpQ+wEL+f/VE7Es85pxcIC
lJi93s1N1MN4pTV/C46x1K4SEaGOl5XDhDa5vxvW4JSPpFhFu8X2Z2ETyqE8zVALvYRp2SaOnnf1
B85MbmwUaF3FcDsGX/75rANZ5nqe/04M2HyHJPMCHA4GccgpPdgVOFLd4DIuLqxvtFcLK9RFisTR
nDg1t52sBPasr9jWeeQ1v4Z/wHDTnB+aUVXWE6yL+UVsnFgR/OWr5keoRHJeKDs0eQsrndQJlTg9
YwVrxb342cSPhwxIGJPe/wEI2z+NSA3URbEQEP/3kNM1WSsoSW5If/ADSkcxSGMOfZhysY/IQUnL
1YL2aZYBX8JZ1KS9iRK5ao+szHtmNBMHnrsY26dNkdM14r0hF0QmGfMzMMEKtjuLeJkV/QbPR0Xy
htxjHCOKAvkhg2FxZGFGw4CTXXSZnIX7HAwSSUrPDAsoFGvDbg8sE14Fskbyg08rf+vqdXHPnvw2
YogqX2md97BUFvrGkCey2CU4YgHsXBAbCzbVXC5sysdr/U3p+W65Mi34AYlAnbuLPKj+NfqNC6Jb
KzlT/DCnoOvOX+7pu5dRk6iyG/nMf8iNpZWnc+3O5bHbMvEmPX9hRXtcU8f/1KnehV6RcS4C5v6o
YmL3uvKkmgGF0Qr9sy7b4M1XDhGpV2NntiGgZ0gqlPz1qk2gOpLiv3bx6rAiBQ6KNVrTNzw+rMS1
MupmTrVX/A7Y5QQRrjLlv4kbcuyF+Il9aTtXMfHUsiLQjR2kLNQOhDy0K06LUh7nM3ntrWn+I77Y
WAKJdaFX0FAedxqZR8dJ0kq+2DptluQIIegLew8b0G9oM643kPPtDOnF2QYBIODfNjox52FyjWaL
16xyKu8pSunDWahQ3NONdxPoyWDCxjHtu2tcWOaWuhUURuhTR0QclO23BrXLXpT+TX5k/wjMJUYd
g4UMla+mDBWBqmSMN4uyOVgkFljLPb5YXSIkGcvRfHcmSIvjyXvZjh6N2Rd8v5gBNqdOfT9RCr6Y
l/YP9rdKOGKpz3Q5c1DkWdLyWrOghFQDxXMtKB8vrOJ9svGKIkUkYcU0xuey0S+d8N/06kskpDHp
cPQNR+IWRCUodIR7qKVSfPhH6OOtHVESWSlU59VbL6UQeeFVRkyeS1OHxXy02/yi3lIZEPeZc4Y+
zYRR4xv+rvStul3/2zzfdyH8WCMJXmC6yStwXaXYCrAWkimVkMhJSdNQWwm1qBsg4q9YAgn1dBpP
sb0phPQz28fF5F6+0GwnnqyrGH8twS0yM6HbB9cZ7NhyfSxthlVvhja4bqRrSdJxj51Gya2iGLVj
FLFehNuea5n39QmtdZ7ULKEWfnln6km3GlyjWmhr1A6Q2IBZPFsMA6zIpkisjLUXkfj3/Rgd1Rm9
VGwp2Tjhl51Y2L76brd2FwF8GoqbngA/eHFo+Nx5zi8+6RO67E420oELItoylXpio/QUjDIFTOPJ
ImoyGgg9B9LxxTxbT+qETLyrZA9U111+eJxTGNw7U0MxaPQNVYgqlih/V34B5OLU88N6waonW+jH
+P3gCOTFob99FB68iGUefCuEZzhB3DzpMNXN55tk8/YnHYY2DFyK0lfIdnAlqatqqL3sPKWbGCRu
rBb0qdDfgvKezqOBCCgxK2e95hg7iLB6KNpuBJyB2qbU3SJ2QNdDq5cPgyNJ3X7EsKczPyND2R6D
zH7phizYakslOdKKEUBKvq6LnrKTYaNiaKVfqlzZAecoaJ9OHEKI/DzONilzm7mUebLUukakJzHD
5oBeJ891xrUhEfAA85yt9VNCfC6EBnlHWGZ7UBHQh12g0ZNxurQXnns4b8ROKLk+IrONa5Jj1yD5
f7w5h9fXB1wZCMg7ziLzDcqBFdF/3UfmeUi8qUe++5XB3hHfJSgqMwet4hEU3kWVVF5P951YA7aw
iey7AQ3FNLm0ChckIRFDGT7cPZKMOdaGg9FjHR8g12tAn6A3S44qpAI5bLg8vGZUIPJU6d4qUb7d
uRgdF1q0cKhuvzNrPGphrk8SUbaNKvMYvnfRCOtp+MQjyZoDS6bhoso6Pv4fS91ECy5zIzvByq4u
9Yw8ZKi5+Q67OfejAtlMrXB8bBfNYHsTcPU5DTf1p0tG4saH3jhYGd5SrPNYvCVMwa4BLpZQ7nxl
tG93o324m2rIUwtaCSUyjbBnmxHCR5KDuZ0MuV0vtvHs1WmB4ldcqer8V+bMpChtGcunT0Z2muka
qRMcexLYdTOYGK6RyxZgJrnDzrNpLqQFgeAWQTsfDCs7Z+zSRkQEOTXQo0Vu1lLKE2gvFKZ4Bq2/
3LeQwWWIT4HxnNPMzSywm++UMNlXzr2BMFJzJuujCaR7V5PDpRu5juAMKaH5tajGdqKn6SytpEre
uEw2DuMsoXcFJC39ABnIR4pAl3hppEI2oOZSxUf1BVjxDW/SW3nJm3mYcvC7z8M6M8Bsaj6P1zj+
+bQ3cGOHhc4bmsqbFd+nwuMoYj2Q1UnBOjDWWbmJjWF48PId+kK2V03Gd26KGyZLYQlaiK1WOhee
8NFjrdmDltgkUtRWe5+CTZeTSXS1GQBPkEdkCT2p/r4rFr0lV9PbSNVQADvrDZ04YwTtqEb7FV6T
y7Oa3WxOJ883fM4eMlq6nEgqxMSn0X+P0dT8iS3UwcSECf3OB70Kmsz/HtD1EsDpfwfbFAzGdrUu
nIcmxw6iV6S0iYGP0xE2uPANPJ2tCXvrvBXUiNwKYf6Qzet6O1PrQJnZ5IXTFJe3FnXvg8HBe0IF
HU43JNC4yiYo1ypJZ2L9v/t0cHnzdv9ni8kw94XMZadnN563ZE2U/DYZSFsysb4sQzzrvskN0+Cu
bqfgIxIVJ+zUsnzf7BxkjX67HDdOrHbZK0oiFmb+ZD22WWy40eIcxH5/4kP4zPLExMz1Av9CjDPM
BrJ3NPBhDrfj72UCZ9oy0IomEq6FZBwYCNDw2Q3YYtEtQ19zVr6ISdBOYimWuHpeUdT97y2uoBlh
vWcwDmPmt0bnCtjuDGQhqSq97Asdim5x2r0M9dGRd8nGHPKUwIttFzzmmo5tXPFwKTlDIeAGtdy8
Xp9rxJ5egXgqvV7TMAX54VrLww0Pk1COyIs5/6gkmgEtMZ9NI4mW48wSFYK6GCPgHihhdKxynQtH
cBW1Tv5//zzgrG/G9M1vUbMPsE3R9IPHW7nncLV2efnnmSDa9pX43nnu4qN/p1ySkJDiHAbqsUEK
AR42/0D9ngfDXuwpwMxwYUHOZsMh9lARAechLsMiss1gXZLD6ONpzTZ0fEb326/0S/Kl8A/sm0CD
2j7IN6MPlweciWGCz2hl+pQtNav10kcaHJ4G+4FrkBDngd/w0X1DhPN8X8q9kazv3K7iHWFK1qpG
gS7Oi8H539/D2UgIgv89Wr7ucCuT7TYQ/1dkTSLrxByka6vXUFe5kqrXE89gAnzwhN4dO1P9SeCw
QNeNEpDlh54fDlkFNqLPWk+wmwi7HEsW3qB1uys+nHWDu/k0goMMjXI5ZjqDOZ3URU1XRUAtOpmb
ynXqfkvgCKi3rRs7qma3TvM0pGv/gdflHIPLJdpd2S97nwrdLD4UePcqEJeCwDbLYs47PtlvLa4I
yDU6b3DWL+/rBWyYC4Sput3q1LEECTsMkkwtRZ6Cw9B7oK2AzazVkoYHVBLq1S3dWNyVUN3T9dtE
1NonJiIcTEHC71X14af8s1gpz4YRqHUNzVltpmuXUlv3njYZMZ6chcQSESXu/ePW1D/0I9S6zA58
AxO4Q6HpjINTGO8GHSY5lTKzgYpYF/OMJXKlp7bktC/KXvJ96jdCVaS6JJ7LSO8FoN4OphPmza+o
9jYEUPlmeb/mtX/OQ6yT+8qevos5jCPJUc3ge+ncn6EjKe5GYYHzYmQuIA/S1aJsW3qvVmT5WwF5
DzWRe+uSfRBinO01m5al5uXM6ZcHUFGeg7WjAqBi7r1a5+uc+lvcc5/GwU8pmBsx+mEN5tyq62zV
8gw7zQx7dMu99KZ6cD+KzldcHpvUG+Mbz8iTC+LygpMW4WxQfvdBfLR779SPjx0RZzdnIweMWZt3
RXj7tw9mpVqdXBqtb/ZBuSMisJ3QOwUQtpWRgV5jRMpmchwqgD7Iq9+1umYxuoLPtqpt+wc7ErKU
MCIiZo+zj4D4GHOaHHhW/nTJD77ENHsFiQTP8EjQTe9IYISLnSdjtyUjqS1jfjtxmYk3J7v+a+bd
ED9nKqgSfbK3y94nRjPW5WXsn2BoE8xku4kchZf5rI76tmFtiY8EV1CrphKgOGdGdTpwbpzuyBNH
2xot1EmzkJI1ss6Oz04HwPwHE+OhTf6VKpMqdZ1Hxbq+MrDjTlKsqxSPPRQWFX4WhmEmTzPUhjtZ
j/Ah+iCDs+iYQOqmY51vtNH3DFtExc2ndejP25YQbv+SI+ZPEcUVpR7HzDShU+SYW2fz9oFZKce7
+pXkIgeOhUQEY4EALITFpi7oWaiox9ZL/ryrWrHjswUgiaq+GOI9/jdnL0DfxtUbJSutxaEIno7P
Vm38MRnAwGFTGV8JAbGNI8euzVIbWBOZOzoXTiw7NuW/tgAzGmsHrTivCZfqExIW6arHq1ozmIk2
rGFg94QfTBebX7C5DLDrmw7qNaC4wL+1QxISI2GDlA2EOOykcMliYQl41GNNFAGR1etqAuu6sXoQ
iRLGgkcwxLkiAq0IRp/DJATlDrzdD+0WRPJR46cRrWwnb+gIQJ1IKGaudY3m+40YOkH481p2Cp/p
z7l2ncVFekwM6aLCCVCWPvamA0rIzVOJAw6Qv1dZQZneKNEFeQhtie369WxXfuEOoh8+Vpn6JRNk
rtF6O1k4TPXHgQZ1hnRIhmHgbdGSQwzvqebMIAimpWB+bRdeAwiItNX1GA0sbT+S11/dBATbIRLB
LDb8eMikdPBAvRIOwks0gVYLnCjvCBEELv37Gv9hAsjb9PTgNiZvD48YDOongTYaH41QYz9gLg7r
KGu9AasgOmiOm3a7SqDdAt9/HOVxGRYxfJ/3xgpq1M7+5AleLl3XdvKU3Z7InGwtOR4R038B5cgA
0aMFrYtMFzRSbQAGnSmNonFXUvx5fuIuH9ibZB1C0Uzi+PuaSZSEL/olU7IMH6Gf2pPf+3IBAmtb
n0WskpXaGyU9q4nWpT/LT4Z5Wu/8lHTQ2CMB4wsmZn5x/nvEnACA/1p2eYQKtadYJSdYAQ6TAwyU
RRgEXXU9sKhuM2YFRivytyh503NX3QPX2PwFW/UJSsrjzMGtXD660S18EfreLGHSGD/K3SCP/kB0
n5czFJBf7v/8AIHMYXRnJTQGU6dzWBhc9mfel4uiAXEuCcKkSE/UJ9oP1mzS8ZHvgdbveX8S0Ol5
WXMDx3ZfDwEjkCBNIddJVUjVp1Psjf16Z+w5MCIlV27hCXqmQ4Cul1SKRDkC3j6LLf6M+3bDe5Qw
vHrY2uM89AYxGBE6jwVrVFw4vqBxAkv7rp/rG8j5CaTRbfhHM/8jOkGR997ncd/XVZti/Q2Cw9Ow
xKpbeGopcOKKp51ZO82k/IyOoFHp67aRR3qGGLg1RgT6Chf/lvEAsVjdxFAW+05HvDjD+kvsvQsb
iZ8rDCFpSuUWybR2Zt3uDIeI54gHofP212XE1BPx6Kb8//je4Yam2cir6QLivSObxRgUVu+10w2S
KJEvkgD1c8WkV24OSzQSj43KcM/IJ8v93ZEMi9+xBDLr1zcjB2cWO9xTG4hPnPsyVgR6l2bF/JxE
h2SioXKJkVMFk3kMGVpzBw1YxsUCGohcm1zSrvKKxmzOxngNpzPZjXeI0a1pffN9POGowh6yqgrH
2LT0izG+nsH6mekLNbr62sYZRcrFwKESLBl9EjUmjp6LNFXMkfdgZv8Pl31goojUR7FGu9bNF68E
DYU9shFzO97tLWrdtobieYhYW+4eP83ptXPMuN1iquAKphW0h9g1pTOPkndfvShiykJY7oyMGi5q
REJUwa6XNfyEBgR4Z/i2WbqwJ4SYfbkUvlaqvHKX2aPlV1pIOnRw19ynakxqC6Ar/QQFKjb4Ujri
2EKoxLaIyULxBAYYrrrYkNuqmx37yaFmPFMpV2wBtIQGzxfqmrKADwWLjX6A5xDoaKzPK9mgubob
tQNsMKLrZ0DRiG3U4xZTn5ZoYfabsRJBLGoaZLa5Fa3fuxuqE54LdSRBS14igcNm6meu4/kGqgap
oT9FG0tXASCeRdTFmlP/IaiDBAUfRP1ogrr8uW8OWgJCrPSoB6SjRJOj+ETr3drmW7bCeazPNXlA
iAYvcVkB2ZBWLQGq+qaq+k8s8coIcLpjoN4Nmkf0aHDaPE29vOuROEy3XionE+BcO5mt2XohPxuy
vAapsoyN3KgpTR228r5fyaO3auYDBt+hbCWUniKTSOV1aHcrRn//VGO3rqQpAQ8HSjMe3thRecVf
PvCNfPV2RPQsqcpM4KqoHURGzHDuFJa7zQWNMtqosqiQ0/Z+OLaM+x6QDenbEY6yKc3T1EucVKxv
RFjy6Mam0vbcZ0WuhNhVuPWoY3EaDmp8iWC+uY+lkp4K70ktjiZhY8m4x5LU4yQbXufxHPGYrE2W
kzNFJUmjlnPhgqeLCJJ+kDCp6nO4xBrzq0HNw26iY8hVYE/TQ3rUP9LuFU+vc8U3ujV7CQdWOOYs
fIChO+KdMwisya3pq9dzGtpRmX0OJVRgunkGEQxbanMfqUCy8GAsxqnn6cGzRFiAi1lgl54pQNEw
6iB4WmHnDFBC1BC3IfY1l+clm5SlRT582qeRljDhkIOVEGFIp2S9fbwwftm690Kfhl9bzDLSFsUG
gKIFLgFQkf9yb1zBhoOIZTCTD24cmZJbz6XFimTe85bxsItqhQPEffEGqULsXgI7/s0WASV2Eezq
y2nUVav6pLlqQVfhu01Iy4yhUQCQJGNBanQtn38WKRDXV25vWVAvEdAJa/PE46BKb/rCPARaE+jm
nL1Kq6Cf5yMEK4/dx0seBrNX93e7HX2fe2SxIVFw/fsmPOZzVOsfcYLrBWftCpjteqjr2qxah5KT
CxJFqUPhHkHrax3PCvZ+Mn1HzeB2KbW7sR/MhSSUhoZW/AMmDDApWkKM2fGAhI8S6PyTfnbSW68E
+3WYFI7If7tFE2o3P9zf1YYNVip3PeK7xD27LBI+sSuRxOQMTb+5yzkyVRQaVXHRONfljVgwr0AN
4xjOxzu+iIj7PDT3rZyV90ELMQ8Fc646koeuwUcYIghFzcp2qhpMfx1rAZgbUROr9/54B3CyfIPP
y8e8/5BmkNm0FsUPO7P0NvTZd2Wm43QjE5L4VifPfG/hbBPqn+hNBgMDSZ+88WkMiYqwvFI7RhBJ
XhQhOb6yOPAukYrWupQkOI+3hptUyNO6VbEBlQP9KAP5gZP3CwqfXwtGY66+LLJy47VVsCjlZorg
lh4RBKj1fLenJO7/owCcnqxA8L+v3mxq87dB7gUM2wG3/QoYq7sMzrzPRiaXDDmAG3wZSihHhZ1R
2Vdp7lM6VYNOo6yk/jaT6ZilddMEJcxx8I2AuVU9kB/df5XfH7Y2wniIibhnu+0Fyfh99yHwN+51
zUWQF7pW65fDUYt19fKol3T2E3R6S3uIHB/DkzRfEH2fp4kzffL4HX68xo/3H7ezZogL59Q8NSdO
ZZk2J+37szrsl2eLa7rjg6gCzgIEmmwFgj4/EQtP9W9vmvHsFf9aL72hedmdwhmvXrg4lRrnfVWh
ReXYXTJLNV+ZJvNfIBjLRBV1LCGAsGsUHGYvzxJUkxcW6461ztP+diiny/HtvbxQDqoWJkjenaO4
sBAcYN/70ISgq/Y/z1Vdww/78KAIX8he1Gi9EYLe1RPYhny/PLzCaKVO/SNi3Rj4uAl3sDNx7VDt
6OGIEpFrMZ6B48SsGEg3SO6jkB2jViE3mK6ZdDpwKc34egnwbXzys5h/j81dRv72ZHRdC0kjtq1f
iLAwpAIwaAaR9SF3B5PS3ljgO6E1NYTKbOEJdW0pNHcOMsb1DRXpLKYWLsipUBxAQ2y6KQnu6J/O
kk4Na7AhrG8Zdmm1yArwQg8HJs8S5Q0nfNZuUkQqZaN0UlHx5sTwLuOSaP5hzptRc71rDmlG+Nxs
BNcoPd0V/XQh4MogqQiHfDD4tR9rY/hkQE+6ine2/2w+JlDcSDwVUWE9kQGvbYjxq8xMM0s8XU7Y
+sn8YC1JCqSHr0HBh+C/R0jPSy0U+FRQ5nwC2wFmV4pqzpzAS3UQC4qnd12lag2fx4fw1hhh3MXr
JldQ6G+oofyCk8YSiVO0JlhymJsgT9u8fA+Eh2Uk6+oTJ6fiVjRmk2LbVDZJC67UicFb9RwJEb6h
SCLkEsA/Tq8Zr0qI6NPtza7jvoF9g8mD8sD5KGgvu8XqfY2sQ0qNAZDKAOOHa1kpxFA4PNZiupr8
NrTWWfygz+2ATcC0bgPElkEyIfUJHXGpjL4dw/qtE9C0gG3wB1mDXikhUWmaLqSPxKLGE227yeQ2
JbI/RXkRpk6FzGjjrMoTZkpd9rKHWQ1I9K7ZLNM3B7IsUo92Sp1EFYNcPOucJ9qiUT3xbGT2qV5n
2oZIoojGPhru+YHrUjGdXGBduOFtLQxpNxdT6wVgODuRvF9jLI+9G92L+iqzXTxHT7g9KTDeW5Mt
sH9O4Gw+lOw80WWe+n2QGXRBh5Fl5LZ+JfoclaAZuG+/a+w47Zic4j/1BuJmfHHHb6Sefx57UQ5S
KonmGYljtaggkFOXuBDy46g8NVDNufHcf0MCZiD+WLyP2TqjLD5T1XJ8ylQJvIhmX08NuCKSh9wl
vTgqfPxH7Q9aCHF+HxyELTIk9wWsd934ncy1rOTk/GlEeH6ISzK9S6VIvrdHn32zVB3RueZRKD7w
qVCQCvlbFdGWxBTVYkc+IJKcFF6qeNht1dYnGkVPRi4ITEpeEsN0uQVz13KMGaVcMyD87of/RF9o
4TEIfboRQm4fhv1mfHomEkL4WsbEmN+CQgYxVZYHV3aeYeZJTdpoHHIQxexno2FvE1GCE929lQfl
ux74jue52+T0Ys6LuqiU670INCKekx76PaVElkDNDkP7fGXSyTaqr0EB+EEeCA53lUJCtW1aA6WI
9jJWgdRL9kNXRWCx9nBPBI/s6QzLenX264aPEBDQ0xn0Y7eeti0NAJdpOgtpV9r84F7e+veNEv0o
SY6X5cVFqbrEKd7W5J6oeddLxvSJ4hOFRf6rMDq1vR5yl52bcWqaQnoa0ppM0QpvzG4GaG1rEKG4
6p3QtrOELTcqcZ5UPHFzawNNNG8SBxTU8dV0NPysDuFo9TxA9ilBzhlXKOznhtAtEHjbMuTRi/Af
WT5Rt/Bc7TfiZaOJLgo/fwuybljWQRuWV8yiDMUaPCy4PpGDvPF/bIlN4vaCRNiyvvpFS2EYorcg
rz7BCR6/zdUaJcCOe49GrDjrc2s/K7wNrZIwOm5xKSKvciTFza+V7F7Tyfpn+Lo5m4ii7LrYuKl6
Ri0C6Asvupr6aa/v5XVbvQAHyIaB8xdxMGGD5z5WWyDClWscjEcRBqMEpoEq0FelvbiH0G0aNNUz
QnIW+T1/EwgR/9NfV/Yy890YAWS+O1oBTKIursPAScJoPs7rksrnesMHLZQijKfqPm46TL9NhBb0
GLGra6WeNgjCAJLXaCJ3DHXI8MLn3rYXzlNpMkIb9jX2+3G97mXED8IOzR7457ntIPGfeF43ne6E
bDC4vgHv5hP/AHDyiBCQ/gbpDYp32qtH4t2qmwc6bzg5LMtLGUulcMjgzk45TP5USYC8V135AkwF
Nv/arauBtkjoLky751yozf1aIpDaFja+9f+dAFhQP4WGrCe+rBt9vHayk8iSK/vJIJd43qHQPGVq
DCz0pPlPJpBy6cW0fEYPfp6VeTl9sEFh9bLqDJUshFeBIGdTT1aswfzBwIq1feb/D8SXDgrlpQbV
zT2gY4l9Jjz9khDmK+IcDHlq8eBW4f9Axq5IhXxjjo8QKYJrLiGlktFoeYKkDGQZ2IKjnIVEE9MZ
7OF+m307Nh8QMkqNJ7/+1mbup2uBSKmvaomW39hj+HjEp9bwKMIDPkSXuvOQWA+SMYXoBWD4kJhr
E/72M6oG+K4PmMIAl8NSe8ZxHmtV1ES8cYhJVXbWgyYk8Gd3Fec0MihZy4L9qprtwm16R1Va1216
LJjjI7YJfsPQZ4kuNO3iuvvUkd6mQs4vf5kO0d3xMPo7oSltil+G/90IXSjwAXQLeayy5SFSyycl
Zh4PzbjKmFeS+SQDz4iwNz1HPYoXbWfeHqpGxYBk6YdXZprXs8icUJmEpcC3ez+h8GxrUDzw0oyC
0xunT//wtp2C6+z6kV1gvGF6XWqsjtlbTi0kmHspytWKTne8HEZ7qt9XMVzILNmx0j2pepkIc40u
9Ti4XX315r4A0yD/mvV258vcR+lyEfK5XLVbBVDyCDCY9KssW9QlR3x5eU2d0v8DmoOVF3T8wMRg
8WF+DdbV3KgCXnNumiFArXu1djbg5N34/iZdxk5KwuJvpe2thjyVsZ+vY/Q81SiRg1fTbVfX+rMM
uBjwxDO9Jv/1twGX6sYlXtOqj9eJhHTaJeUXWjAp7Rs/5bJY9g3m2fU6MVdY22nu1oJmfouun0q1
Drs8M8VsYocOVlQP7a0A8TiCuTGscVJ/gREc+7r1N5uqzCU/2j8sjiydZRiQvbja+eCaB+UD7/xU
WedF7ADrPNBNxTy+0RX9n4CNajugmfXspl8eB8LVMmZ/fWbeG3UZ/PXwW7GfWg41rnQrVV/IfYma
jqgqDaiH7iylujWPN3+7hAZWMAVFEYlG3eg3PmmwqfytYSt/ss+ziZnYO/MMlMaX1y5JJuj0JlTQ
SWBdIe2x/7+drLaW8dbcHQcETHW5YtuENtTtwqJAdSIG6yHmQQE0kgCcnkyH1yhKYro94bf7JPPc
7Sz9CRGCA/YoJvBAiHFqtz9AtGE0O++T87O0eu/KJxF1ChFquf8eTpcD32aJHIEyT9cAMasqtRXz
LLMzSh+KKdqFjODlZqrVveTuJslyenxalA0x68OcJt4SQedc9l8ahV1T4JT+88mepEs1L+vj5Pqc
n1YLbiDi7QO8gNiyB9RKoA7IRfJHrm2zwFWLgiNuDEalSPI9WidJ3/w0lLllUoi1aCThgQ5gGyik
Qy3xBW9glcKVY8DQKVnLEoHQHiGqZog9mYVGl+pl7utvq7Jxlaho4jWVBcFr/WFPBC9FJ0R5Oop9
nhx3rOgZUhjOSel7d43pjqsR+W+RzdE8u0qUSULVD3W66HapQNQ7SYB4clG+0qWuvYSjfVDXkluk
K/ROG5ldTSy/MVQmn4DTsyZFrxo7gjMjMTscd4TYnPTXO4tYAJFFb1KXIR8RTfwUqzTHw1Z36OTf
E9dZx1ynpSiC/4Dh852/XP6r/1Gk6YcxbmtixxpZpK+hsyF8nfqS5FX96aHGlBua3zmHWwuccUaL
FJn14VLGmi8NfH5wm8fYEETxMIWebcT8OWxV64M0CdtVIVzwGAiwOdpHBfHKp8D7pgxxobbP488M
D5KVPwZNa4Xw15fZHWGX48NEP77KRaE2OOmCE4qMIwy5veDgWODgPZeHmpLNLRJfbj9od46Ogfmk
hqsy+nLnFF/DBNbZeLUcOGX2J4Hnh7msUvTKj0wEjmB2UVsvdSaLuP9yyTzQibgxj19M/GIp+nr9
ICH1carS/5xLTtmIGQpqWYVgL4MQcQheT2T53py1Df9UAvGmJBD1yJuXLwhpP27HmmC8FzTXRFVQ
w55ppv0wLveZ2zbh+JUnXcbTVBOmIWk0dGGnTTUfrc0e49Fo8AT3Tz7Y5OJ+xu1uoIHh3jxxrMW4
rNhjWHH3rTdN438Akpx8hEf+8vtQ0zVY+NzO8IHJQ1a4bQuwIUgjo2Y/SJtbS21ov3lrq46EJSbT
ZD1HqSxrdJYdSW0BmzIPF+U8tUOHsauDMw+AYqRKjAwdKYP2i2al+rOQra1oyWeW6Ut94K2g+Wz7
PpQgnkwYF5+iCJXn/KBKKSG1h6Fze16q/ZBnQZgVv8q4tgOnpzLSQ72jc3F2XHl0DYHEC5Kf2xUm
dgHzLUIffOMtEtWly2wzk2ph6Y/4uhOorPj9KUrxTkoXwPIrEdReZ0GUbVzSH7pTiut3d+D93Mtb
bW+0yQTa+XRW1ekSXxGL1KElgyDlpZgksUQHlG1gB/Nk8b6FdDO1hfR9Ct2OFqwvfVUEYf6hGvz3
JvF5ydzqJgPj+U8lHmRdMKH7be1BE4WIrcL06WuFN+u5Dap9eJE23ikp1m8jsZUgBpB+7kXhN7pG
xt5VDTyKZFJXNCaZ1JHyyk49yBBmm+m+STqm6yw6pSRtmPrnyMxLO77/TTSMa7JcZYMlohc1GlD6
HIcFQVVucWrHadz8sEunsd/NQdguDpsF1iP2lZlO/zE++ucryvndhaa4NAF96impTP8ZZKElYZGH
3tF67pnTkLCbxr+eMY92UAPYxJtw0IoJBpwkbpfaMJ6nWrL1wAc8GIt1x4A6cu1aO76dUSTMxCZT
BIwiPvW4rXoeej3mOC6Gkn4BCrhuEnfGdZO2No5ILT4UqVaoEyh41fW9VyBFf1Ndd0nTR+MVGQwB
xapkuFOn84MES2lrpca4GLhPROY4apwByYJ3gwr2x3gtWlumEtGdFM7TqdeE+HF9+WBnPORrZSjE
hWGk/RKjeFWgFJclCekZ+OU5/AekBQXSh1lIbYjdhts6zqqQPm/M28fau05ZBv9BsZyI0bqUXkPG
5CxHKSZBrKAuBz5hvFqWaMDrITczYB5sW1CRW0gNIXU7H8GCMumbx04NiXvWwgOzv/ot6/FrvboB
1Evi4uZYp9QaLFfavk7RfwoMpAZjxXIrLIVwL1OVFkhLEzXu5FlENm9H/RGBn3FwOhSCyNd9d/L3
/etmBsOmMX5wBIZzdlOsb8cUqw3c60rnkJla1TPfa79W9VZpIORjFOsGVrdzuq4O9J4v3lJ4qX+1
Gfmhv8cInpQxxxkQC295G0OlCaZXSMwORybwmDfRJuCKDqgPqY6V9nVvHu9UBGrlMPwJ/C2cGbwe
ufwofDNvq/UkTQt9tJV85BYovDafxAFYnKc0JHw6eVf6Bg9upMnGhz4060mx7/OjnulNxcmDsXnV
6ettyIabraeLpBMsuqwiF6LzeaH89hOdK2PmoPz+EJX0NXtcQBR6ASYS6Vbi6Z1yyTgNgK/dT7rr
21tz96NczhgmPb/Cwz29NXWtyqWPRBw089VpYTppwwiELjcTLD9CS7M0McTCGrXU5qY6Fa6OCnCK
aJ8vc/vd8BjayRhZQqTCS2HV+0MJVQTYPghAYJDzSagoDUjuruVzo+8617dlqU99cvhX8kUiqE7a
9u3Z8mf40Dn/YCOv65F+OTmUjbN7XCOhBMrRqnOHLQczuNUq/feHluK/UPCyC6MVGfnxjZDBgmqI
SjlovwNfWYoXAGT2v65fjN7Oc8jIfWMG8/xqNCrg813Tt0hoUVmbiBCk+gJyM9xm20HapDote2yq
J8g0GSgumiJD+m3vuu80BMcHJ8IeHV7wSe0vm5MWyaedCcDE6QUneX4I9FyCfgVK/iQvBL3WNIZe
aU0WJXBmCcXCv/JvFmhxnloSLGJe3wf0LfEMGHbOUB7aVq2MPRORlFu2m9a7JoWkukxKh/YLg7To
YAwvi9LfFXNOpqBp91NFoYkw6Dh7RC22YRr7L707Mc09mXGlHsJu/lEicR6Eo8kfbFWnhmdgaPMl
XUKYbz+nSZ0j+MjJ8NZHIgsopvWkmttgo4tb8EYz0UCwXkXRew/lVFxADVucSeBYrjCmdWq3QJRa
f6YQITNj+B4WJm9k3zSNr8CszcsfPgTFvU4t/KJ/2v4qtBy5b5Epd04rEwYxQc+DASqqrSLeKr2H
+L5EvdorFP9R1CxYasUMzw8MuqQP5XuWF6YhweD151mI2yY/Qz77nvD3ugjUrO6XKeOfpc7wE55n
oX2ybA9VFx/2LPHaT+Gnyfi9TTVfrQEMmO/iWjGvrHwD5Y/deKJWeSriq9LyFchFXPKrHyW5VOEQ
qfVqiEwJpNy5NvnjDy6qhudJwunicn+idH7oXRoLqxw7SgJEUPOAtHk3VROMBnK/jZgAtHfSO5YZ
QVNQEWEKuBbihFWU0ctmudFNiFKBT2CSEH6On1ILgLQvGx7iz3bAb05TMSGi7taNazAtJR1Rok+u
BV6Bsxk0KPDxLZmA8yPChnopmszcRc6wp+7sjMR65r2LL9d+Hmn2V/WgeuJADDUduTyH4agkommk
Y35m5VMEs6hk+XEH588CfLpiCWZU3mwUHeEOb82v98HNAiYbbNHg3/Tl9//1g5pPLogGLZbW2XqF
r0lVRgEzK0S3qhU4g0G0OB/WzP+Ro4iE5cV4glnlB1I2zUO/xuPpie7eYJOdiITQ/kzMKcBWMfCP
tTfAUclaH25lrojp7Y3D48givaQz/A1IjmqbOyDMTSS2X0jlvauN8SI8hByEErrDHez/BCNGuXwp
2p82BNXdaJYuuwaO/fKf9fSZxTGXJm6Ryj6tQuGaFYx7bs/p8zfKoF3Gczy5Yeh4k5x2uA/dA7g+
ogQOpD6bhswbWrXWU/sHEaFOoL5S5lUTQqEVI8Lz0VtpJ0PPYsQlRwLBNwKrQSgAsc+Bwc2d7Eeh
ipVzOxk5KB37LjGSFitPHX5EBCOwZDK/M0mwwZVjFMuwRHT0Bd8l8XKoK7oLVQYBa7xD4zRnMbc8
LpY10XKlIODQvOQjTvXEGIgaelVtxvM1dEUSomHLksO6UQ+P2sI0olFHK4XGNpdU5x6YXT5uXzQO
d8tq+exzjZ10P2t8TW5qCfpbjTIiIovOh70DMR0/qvyhnOVICjtuxqAKFadPjU30eNCsqJWNtROJ
h4kj2KAfD2Ax4LCnr+vfK9iv3IJ7RhmFed7s0L0Hdy7SUJ5XYbtfd9jC/szGGhhCQTqCQMefASOm
kc6woOAtsHW4/DCq6ykbxMYSO2r71P90CusVWCFhQn9fIWOE0kQxJUJnPceyrRWbVYE84/UvEWRy
2DjWwJ9NyJjHy7Qi3SHBRHDCZS+S6HkX02EsmCiQehyO1FvugCQEOQ00gYMSEkvUrCDeRGh+OtnK
zY5Ux5RAYAk7+l3XYrqLD3tyNc9sP0YoAaxnQSETTmK5RD6KBPVuqG2w+3hig5qFLLmDixnfhNTu
53wbNuqYSCu1+99xKYRnI8Oo/EVWuIEEIa9oF8ZIYrqMmU8GIpcw6bAsPgEaB+/xBJTa7Kkf7q+g
7WcRQjEfvKcGR+YtYQdoBcXZVFU2f6PHQosgX+/cKgKNy3PtjedqGYZGkdNwjFzbH8wI8WLWJycE
mh9hk8yBrXO4i/96JNpUcbwBC9CXQyYopmy0qTEG6EGwTptJdWG5Cj+qXFcBGt3wFoqtZvnm8hW2
gI8rE1lJ1Ckvz7LOYTF/mnDx2k41WaOOkudsskVfVegFCp+ceTep1rghtp3Jaam+Wvt6k62P9BJU
2n5wivdW8ezeLfeUNY7nDtM+oQvX2dZ5JkF5zJnNiOVXIiF36p/wRPFT1NON0G9qNjteBbyhs9nz
t/OBUxSgp+OcbTIN9xph8E8/a+eDA/XzKyVoGE80s94fe6R06Ze8s8jnJ6k0bX8B5c3chzQuwUL6
/8yrJGBlsfjBbDY9OFPdFpDgGOEU1yh6kvisMEmx37vTFFsnCiTl3WhO0BJDRUJQECmgBoFyNCYI
3UsNuqZFxRhMt+myEzVek+fzC58JuPcaq4SLeiVnc/2+e8u6QVehgRftqCu9r/5KrbqHkDtYP6wt
dhsdAsZF8857WtwA4EHg0sL9lhhESqfpcEF/iMSOil3fYAN+nsMd4g3CtvHjF6Q2AkPO6Ce2npc5
0robf9hJLlKPtujphdbt83xc32t8BmchXy/Aur46xkTIcqD6fOnFtPp2nVZSjeh1VWvgjpYVp35f
F4KK7p3R3NogUmkiuGxgGbrrQOV5LGsifVy9GU8o1AxIQRY9mUY3f5O8oQ3NFdAMUxz808+VBNfG
Noig6Q0U1cCD1qpk4YdRB9Bkd4wg3Jqv4e9nhivYKtZC/Q7IG5N3Mgb0RfYH7E0g68p78A2Hk+mu
mudJevytIGhLmf/KmDZ+pcRXhkezWAqVuIXBqJPepWCWsQRZSUGQI7b3et8n/GapW/zplMWE7R6E
Lqo3SpBM/e2sq32Drduy182IUXg36cIxkA2dkR+qrqTJuwTYbYHMJjD9iqGVNP+29rF1nQOZGoYN
TwSpE7eChcGtXL8Z8KJlRJqVCzi/Dw7pqGyLli+yNJYoqh6VmXqTy4lCxi/FKvV+ReZfokllh6ox
b7MoXyzvYXz2+STmiTUOJEkfyGrnwuaF4LwxqsSV0xIqIRyXmrNVFnLlMXpzE8i93B2FWEs8SRhf
RmqrfQF9K8pbnoGeRZt/uswqjIxi4CVHlw3FTjRkLwZSsqOaytK38KgVnfT0NlP0ODSvV5NTAY88
OaxbBi8rDjyxdelIuV0yrU9MvupzdgTfcC7M0cjeBe9jp9X+HuXSaMcYHhIcNEEaaD4hwrEuGMo8
xQBbAw62Vzkvkf7jKf0JaPdVP7gcUXmAhpqqPvLUEwQyxy929Kidqi7QVGoA1DpdSFj7ey+Tmje3
I3AKiNX1CslrfiRBJ8yype60U2krRbDmUVMVD9TJUvQEWVXE4W1Hm/aTFqDMeAbYFlNYQKASRzr9
gKJhdNrP2uCzUvIlH+ppmWFKwnwNsn4PmNaRBQlgUmEMDe4mxUFqC7EkgqGv5umcyIaHIk6iILgm
3DG2t9nqs+zF4zRml5lGqt68ThWnVvAyyF0wY35Y6RfN3jUbC9cbjBup6yJMJr1hPmzVvru1TjRQ
6DsYq9UBcvOYUy9jRAtFmiLvvCOkNCWEsvFw+jB/qbexZdxdv7bEg+FpyDvueZryFI20CXzySotq
13INqZBgepuXoxZG/8rsS3sDdoNRdaT+xedyt12h1PinAsIy364lN6zWZI2Sn7oivOPtUoJW0bBk
4oTJTFh7s95qAzisjoCkE+MaZff4SSiVI66Xc92JhrxvVee+G07oa0T1nxH4WkpwIJymCaKdFmfa
gXHcmlZL/k29NcJfZHNAZEwg5Q9CbXptbSnT4tyL57wRHn3gifQ0N8CZAA3almQksKq7lq8Pp6rY
PbHFCQK81ZSpUoeciancghNaeTqpDt45dayqqEZJBR/hGB2ZQRpeZcAS7WNkn04Rnqhj4zvWWGuB
nt0gwDNfrjYr653NS3rqNi/wl8O17MKUSxBZqMH4o2XuDwRNSfT+1L9fbMk9yaeGCgoXA+xUUeXT
iN0MGUj1f6TmFQAXwHrtITtRAmLfMRpcG5NUUW0xy3quqAYUg7+KeqXUVzDd52lW0GC4gs91hYhr
rhZ4kJgF4tVlVLfuApgYj/zC7/ruU3VHMRpaDP52oktLKFgSI4fdya7gB4aUcrv+3/asPHQBIxGx
+jo+CL6RjtYim2nrZ/t2jXDgspmD1lwe2JW5cBc9lEY0Y7q9VAfqJuGJW+FxvALcku2MK8Z3F+Fd
ayVSV0VlFMXEzPlD8XYJH3ukxerQgTSAjxInaX2yw6rZDozQpX2IglRbYaQFu4owdzV9qhNxvNw+
fLCJZmteE4mOFb1q61ZFd3f0hrZwx4KkfUDXqqJhw6xDqj3IDhKMl6KPU9GX+QHYytJRx+CtJ90h
Vc1DsWKD3Kqd83gh1hGVDT03UThoKCvlFzdL+kTHtk6ir+FdwTvqGtxuKXdTZIQp4/f1zjzCaDKH
a7qQI8qXjuveXnALf6Az+BzQjdYWKSw9vPvcNQST2beQTJ2/5vLPpiwu49+VHn/irW8vuHcpMYlN
xyAGWVU2/MK5AkVrXyFOMniwy5+3L7jwtHq4vCDDZY01oPakg3Z/4PKDvT0/gRGfZLR/tbUvtLOo
sdjIr903LYeWSpWreA5AFxSeVyz/iC7ZAM1ydtKa9xP/Nt3bVf4gu7mIV53Fbnm+OXQ61CoMrnCd
QKW/sVEPXlx8CUIPJNng5xv0c8AKUpTdZv+xlJhz1S01IOi5V0zvf2QonnQge104Iklyy72OgOGG
hjZInUMObGPcq0S8mKkgQtjcRgzJZAZPZdvFQX4GIrlSkwYuQVlxHm5HGySDb0Uw3g9rlRtvANa2
pkOtM+CeMjFz6K0bwMx+P64Qs0z+HIL6Qex31nmOzQius7KzlevJyxWD+2syrHzCf+7Kr5VqbxSZ
dJ9KdgHwBwAuh1/M8IbVYPUDShnQ52eR1RFZxfxnO1r9dAL9lYsAbYT658uZI7AemUZJ1p/qp2fQ
U9KS28wqBJ3c5U7+1Q27YDMsvudS8/OOB2Ki7m0tXZEbogVNiXtO2+Sc4yeHgfIgV1sFmZ6f5aHG
XBWfmJoU4UDoy87sRYBRQ4fcK4wfxiZx830ryp+zUjxk/aqGcfKl3KcEFjdTEm3cuNoLC6vbcJrd
zSmJt+gMipSPf31fKg2H0D793IMZ7gKkmrpwzg8o+GPtBTafd7guih6qgU4w2oTjMU11PXZzbVvP
2cyZvssVJNAM/CwPtnsyuBbT4esC/nR1+8hyqQ2GtZEnr6gbdw8rr/hfy1QvlmcWo4Dye2Oro1Mx
UnYuYR6DYdGMwv2vkeNuYafZRMaJg+VcvrwkUaPyYwtsVsZMmskvaYn2FHhsJMTLs6fZoz1GbhiF
WewN9IBQTPnKiqgLr4PG8XGxtGb91Y2noNTJOUWGIC0iAk1eiQbOX4aMaIxpfs5CvE/wPGRw5VL+
ygFmFx+3B0n1N4/3CxvheEeJX5VOVYaUTFiYDVQCnyOBvw7ZfNptaow9yfYuTvV2DJXaP933MwqZ
3hwlEPbuNTGf0L7iwCf39NmgKg4fuzsre6xp/ropx+Q7/Dtgft8cDI0N4sreB4vkcoVJlPdK4DFp
jYnPARHXzY1DBjumaGxl9HO0c8prr/Nirg4qPQ555MZiy1aMtjQugjoABYLRp2AqMmN8mQlBy36c
5WYls1ooh14ZAyYifpkFgVyfVMhymm1Li3KDwyaNh2CMd7EL4mwwoeeHN9syg94fomRTGgtOL7qc
a+HdZSBgVz0Mnlsa9/PDECrJNxhfKeK/VbUKV+/hjxDR8/GDybmcr7vY0ogfQVG6Y+0ejiSvpYJu
4O7VpY/u+40IZTtj9aL8tjA74AOs3l5AmIgKQ+27c/3cQ6r4o1YY1CnpDIqTaHtvv76f/UMqp5mZ
ll+6BNHB9DW91T0rUg3iJzUS4NPsJhFU3XRVcHzXJ2D1Vv4EbWv16ogE6Tauen27TXZmAey7W40Q
RcHVuZUPRQQ/H1pyd+5brL+1dBw3AXxUmHmO/0jTcf8oSh9kyVaRgm/S3LI3RsuiE8gFgu93vWw5
gTp694e9t4587aZ64q0a1X7KmNqPNsQrSggfm/kp3MNZld1jR/gHtnL3wmmv+SAcf00IwN8iBwh1
arK7afeL5o9PkWm5mS5wgQ5d4fpEz6IeFWN7BO1Ih1Yh897tfhQs4rOo7ybY735+w+O5JvZRB8XC
NMj3/ZbkeKan+FKYQoobDT0eshGGgb3iu/tMiCttdRXutY/eJqp/MMycZhL+0i3w2Tj/d1GZArWn
nB+KFJyu9NJtRD6pMVbsBy2kEnFFdZjOwRdwhogVXLGHvg1y2F1QQ+GJPwsKwao8869loIv/HX2j
zykQAhcMqHqq2Yat+0DkQEGrou0HG8oODxTbzZ6JMkP3Bhf7VT+7s9iHrryQNkeU2Xf31VMZ6/Ns
7CHgz/C2KbThjp/91fjFNsNFB+6khVWibUT1132VDzpZ9j8m5IPWPrcD0cQnhS/La+mBs99OuyG3
JYtpuaE9G/dW27a3XAjohPXhLe29lTsSD0rVasOLycCk7+O2YV6iQr7sxTIOeJaoo65eVT5CbkYp
jWv4gmRkjTM5Aax8ZA/kdSSNJB1+R2kaIGmTR3pcmdM1LmVLVVk+tvAEfHvlQyDXbLlZV9US9qWN
WOyk/A/jtGB4bE9O7t3GO/PpFNn9NigmjObXsyBN/LBOfH/5MIDn3GYYvnVresuXxqFuN/ZaSid4
xdz2FIL9AOWvxBbDObnvEBA4y4fX3ZzuEWqdeDZDoOoaFbvQyl6v2SC4nK7SBTDaDMuwAnbcqP5D
i0e7HSfOnF5jbe3/XE1dyVl9KmWJ2mpP2Pfx6nbf8mHFlCK7km0M4pYFNHwXfTNV5Yhokr3l6Uqn
b1jfuyA8wyTk0k43R26BM8nDWSQFNzQ1YNr8ZiCrY8oQUy9hdcSkgFnX2/xyB0+JXTde886K3GzF
HPGXGrKoG031SYXZiykXJ1/NU3XT5UiVXSPale4T05Hc6Rwka6eyhiSwYGb/8gHMCbxOZTRevAF6
eCEhtPWcFULX7O7liMx4R4rNm5mw6yDUKpphmfxvmEdMNL1qoEJT4+JfGMjgvdzexWqiOiypLuMU
FzvjwbjMwglx+WV5IA9kuRmsiXJ5ZunNuISS5i6UGj6Ng9LIJ3SY1f6nbsdLw90JAfKUVNx6djut
YvBP83FMowH4ORn1QV1sPuO6I+QMwiadlfr/vFXvcQUfaiLt6FEYlxlsRYHykLyO7usGhGpVqZlv
cPa2JeEmcxR4cq9ocSL+VUhIBd7ZLYytsskCH+12V6m1i5Sf5+3KyZ4Wz2b6viMj1ok6gOTW7FVz
U8/j1RrXkjc9HvAA5HbGLyxK6SsGMHezrnSnjptzmNuzMRVdGf7qPEwGW0FRVDajHVrzm0TzU6rm
C5sV+JgdslErKvuIFJ3JWaQYCCBgv1TSSCJP3fgENQylEau3YpJ6d0ZxluCwI5znpK1EW23dA6hn
GFgZbYHuQpEB0WvSlpQHDVcM7qw4FPA9dJsyJNibOW8ioxoPOAY6XdGVVPMJ23kPcuWopIuBnlJp
EYATYhWKTBSO63c6fhGQdCPgv27CE1vo21oXeIVJMNLcNhbHic95170MMwMCUwHNNdTfHvMpYBpP
nfATsr1jLkZT4uviebd4ug9eFwIQR1BMUsymErOkwAZcsV5Ef0XMkuAjIaiyVXPlQNLrMLdQM+ek
rkWrYpg9tlqwmfNcNZU5n2/a9lwueaFg/sV2jJrqkUnaIdO+fLFEjvd1IAJfapoFxw7H3V88ork+
noOHNxEh9jG3IJi7ykJKKI9hRO15VcoHm9FJE5/g3EI6LCMk1mlPh/Hkg6umrxX8pe8VI7dXRF/b
Aeu10Z7K46m1FT6bAVckV+EcS2qQQw7HZwxJSAGBd9Y2v7rf9KV+tGlmLBI4stJyqIMeFjzZ5l11
57wHWVINf+adFStIIggj/h+DP6Dz/lbDoe5B4SzNB8xdrnQXOqEnU6jAWY2P3jr03UI5bz3hBJkq
8J70jFGlSdjCS+WSSybqlShBP4/A7U+B1KMbNE2itunpCmbA9irQofSFdFSDs5vunI8OgJnzAJ5I
p4lQkKu1D9B9GZ62diU+wkCNOrIYWfkd+N84f6KDEPVC3DOeb4vNusSqvWFZvOPerl5u12Kd5rY8
A+GIU1mB39keNRNlwnMVLOFZlK89k5jU1OoQHf/bLMlLpkhXhq+M60qZxNDWgx9W1HLWfDn/PHe8
7y/dc6n9Ck7X7tx8MiFqYH8t0dvtGkHrp3qnPYg9udhACQ0VP6SbVhE6jQ5JzFCvsvjDVucE2Qxs
kDTTQ87yogqKAuiBsdiAaU/G1NHUmqlauZ+7rx+8qSew7ak1igz8JY9AtrfHbTqhj5MAC7L6gIrL
Mb5/jENDlsVNWOFyc7KjV3U8csn+wENhjw0C6/oEJ7IwbpZNsWxWiCRw78iPToB7kQvSYHCvhEVV
ZQfNBuPLqIuS+K3ci+cZhb6ftlOlGGamPlB7hqvLus0ag4bVw2JYZZj2Bqcq68dWBjaTMfZux8rF
bM3infUmYf6abRHh6pu9jlWiDKcKoqpSAXIZqv0QQJTsrecBmxALwJPSfxyCNMYvmRdV50U1LeVg
Z7Oee6rJCBVZ4/db4sWcHi0flN7/y+wnlcF+tuPS+j9SFbIgYRhMANGDQP4wkcpLQnooIGEkdm/l
/xoM5HWEq/mU6Dq/4jaT7CO1gMW4MwmUO0VR8QGIZ+Mk4hq8IUSRzSl3AQQ77aiBdjHOcl5mowZv
LXj3RpOhICWgSCN66FaeGFTkDYUWfB/1FrAkx1YV7Kq+iLTyOdBzqad0RPv+AUkXPkC2Ic+DlysB
K4fvrtuWHABCT1fot2TaR3te3TdjrbqT6i0SZjvTInqB/5dpuWnfmBYza+jK4PvRRerBRtJtc5bL
JlLnGlqbUvkbCN0otACNPwdjRMv1nsJ3je9PP9pNJo9MVSqWDL90V5wA9PL+7ehWzYM85JkPtble
OiQ/ok5WPRHEaiaIARJ4R4aIfZSgu2qMt8ZvM7cAJDTj1AoWnHXUpps9+3gpjPi5Sqv2CbbpvjmG
lqm2EiuxoKk5Si0IuH1h0cy/b7gYaJlvidMEACmvE25tAv+YkZFIPxYwwr3ugkCDxifgD0tZWqu3
uCh21ezp5Xw9rlHKO/aqgxvcAMqSnY9fwmWrn5ZeVHF9UUXt0ehxO1rqvOnNSaudbgudrwz/juC+
oBm73vFoTvxbc6XAekdAilAf2umM+cuMQDcLdSRt/UmjmRDStN1zsgAoQ5BYAr0nN5j+j9NNbJmf
OGkTOjhiBaw8Fyc0ZGe6FUzGanMT20HR+jIYUIK3xInX2N1/ONGyere9sDe90b8G+F6mlvRQa1hT
ObuWoelYg/kjbAKyA9N+ZSiVit9L60jh3FyzWm5kiMIykN/YRzZOAbQZheYuUEHqVdcV4OXoBC3R
H9t0RY1AHYjdszKnplrSO03n6RqS6LvyhK/0UpSNFYpX+/t6B4EgI5dq2PwW6hCaE1QEqm4NFX8s
ehKeWUZ8s3C2SeHs4XxvWyNmpgVQmaj7vqzVzupK6ZhuQCk91gB6X1xjjO/TBnQUzvrsLJgQr1tp
dATriIQeowOtKru7TbHCONCB3lGSuFcgL671MIXH7NUVwzLbZ7SdvyrVecvA67wzX2PpxdoB8QTZ
KWDjov+/YGuTCufyiSvaq3H2JNt4hZPycbDlIW36u2YgOJaf05hZ03MLp8YUkXMHjNvV9XBdvrFB
IhW/UejZbi5pkkQoRSHU2hfTND7cxjwtdGUGsrPzg2+0HONGcpkBwUzvn3KE1SqgU5vZ+k2zAJ7i
963SLiQ1dJk4wH1Haz8Ql3MU/zleSXmP6yJTC1ie8O8y6+35YzDqvhts3yFI/nPK25BqWV4vEuEl
2YwTdlsXbyjmPpP/B8pH3WxbswOxwKRk+ye02904LDupMZDUZT23pJuB1wuIhhxSejU9rzQfDljs
y0DOPacgFWnpltxGUhY9K2n3s8F90p5oO+Jb4NTjhSdNkSNV9o6QFgttpLB+/32HTKGboKYucJJi
5jmLvZa7j1F48kyr9g2EyG7jjqTBYPULF7+bIW0MCAj8GHtGGel2X7gorMc60mOx2spWJzRjNim2
Y4dPktHpePXKQsCP2hR7wuMi8VkCPZleOKmOUDni/iwsa1EeCCn0Q/slUisBuD4eAY78jwB+nioQ
rkjwYyZyz8cbtuu51PbqIDFY6Bo147EGgq6FgLLxlTq0KDyF3XkF0caXWVFs/yYT8/zFEXwya7ql
UGfT5WebZBsGpgPtyGR5VMgqVS8tpfoVsaFtHVk+z9ogZdNH4KBqX67w6JKaZ1Z2uBbm0Ouh4HWv
0++EdmYjfYqR4hYi+TAPhmUkifzt7+Txl+jrRpaiuFe+q63bWhdJsu+EY/C543jG8Xx+OoiGIsgI
rZNaq4W+cruUXtstDgMtyPPdMvS3gYS9RwZcSCtSj/e9TF+HCMKzXP2cxhjvG1Dm7LYp3gDc42b1
v0ltqpZehJV23XvU8STMx/6V+G2l/t8H98T3X40QZUKbX+7oNxJ5bt6+JeS8++ztjR/ENXiXgy6I
J3AO3MxxVRPGzimgeJdoBcdZbnPrroQasXtz0NRc5M7rB/Ka2yHw4O7V6VS2dW5AqO1urkkOtAOL
wpB32YLTtny85DBs6AC2p7f1OAJGmg6Nmn1hufAEMT/jroI4VMrGszhcD5DTLPvOlFfd28JImjuw
pGOqeDMlneuFKHioNEA9xeIVJBnTRkYVB2xEUOdctBMjX2zHxaF5tAs24Hprn/21lfQFrbQiQZI5
WmKy7E4AjG3GCZ42933SRWervTamaFyDcPrBabd2UB/42iF0FJz/hcJsX63KRCwc8tyXb//rYn21
gsmlvCkX3a2Wrvgr4JtEbm9PKrIYyO3DF6CC/vyT7tXKk0ngziwvC0qdHCupJfTKUnIhj7lyELen
18vaO8CQs70OGqelpLBC/3RI6C2xql6mqF0OYyW5ZWBggA+WqDLqERFEMHFEZ7EW0et4JB5D+eK9
zClbpCx3vuJVH3AqIJNwycmJOqipOjpgGFDaGBT8mfqaWC263JmoWZLP8qhKGxftl98+xsp0476t
mjcLbdAmy4OV2m0OYBwJX8Ywj+E1dBQc0SQdNX4Kax66VOnhUUKj8ofeL7hs5NLODKsjOBKQEZXL
JXXRL8lwx0fhNvHVtG4lTYhJekSX28Qj8az6Vs+5DlB4zY58ktLRAOAONoO7jnK146iC4a74dxkd
b6BVRN6h3O/prYrt7iD0+EpWIu7M4I3HgeHbRf8Xia0vfMl4s2bp6urwrpts6/1lqt9lvQZblL8l
uY2/1mCK4Yow4ATe67O4TsdwkBYhcPKqU3rFU8PMfwg5LAYtU3zLGetW6vc7YEBC2Tb6Gil44bVs
YiVqGPvRX0BHr+9z87tE9fTa0jugtsdlkH2LDXADJ0xy/Bp8uoqNzwuIQ4kz0cGr9Ieg3ikhZYDw
2PxbaekshqtjrZxH4PtO6f2Zt8sa8vXy8IERo/ShrQBNeBzYOEr/Wyod3lNz+ieIU+O8aMQyM6gb
esKMSBvXxUgAK9+SuO/lVBo3EEqegHhV8kb26VmrzhKX6R93Q7bo09w0Lr5K4E7cpD4MsW/0KUEW
E9FaTzsYuaVY0r6+JqBKpi2I8yTM46VzduoSmP+ug/CuZqfoF4W/m8erHZ3Z71AiNB7839Du3emy
60xIQIiw7m+I1akiSsvMRjLmFqPscdy+TEP20STVoMekJeShvzTD4kpbe8nU0ZZZB6kxYg0ZNW+W
OrH17BPHRmFOZfPkQjmlZsT9aJwh4nxgtlvSv0qHBPz773GZ5w9yWc6MKpOl1cRzw+8IvcEaZd6u
Ijba8SiZu2ZOy87XUAJ/hUQ0ylhiVgOpw6eUi/S0X66m9xIgNyQvWRKRjUWVit/FWBf4a4wkbckk
MUox/VXsifdoXPnPyuW+LPfG0T+PTkC4fdWluO+35e8ANIWnmyQtsWEugOhrgUlnsOSMhNmxvNZ0
lpVgt5n7InUMNECVh54ItchpHBNfU4ZrqiNRxe2iESupWJLqDT3F+gi5DMmo/3iZeytuFL4tQ3oY
QpFRlTKbUiMq48Fy33WHEnGbHsPHXQ2OPe+Ysd7EwqrXWuBTrTWHNViTvnpIx9C/emZohFeqOHhZ
OpeqpXxmL1rHddNl+zKMWvfER3jTuis7dCaKm6ZdkknvqWK6J6990kMCzmXIgIacz4R66bYAO466
bTtxul56zAVULdZddW2W0gdaFoQVx4hVtxsETJaH4BvZGCmQpjpvJBiRWbdNXFBxFWe0iOcM5TQL
KvSfFiFW2mT6FB+mdDutRy0xTBCNyYMMe9TmJdZpABijIzXvM4QjHs8gwEEL/dClVNL+vK58VewO
A/cihulMoUhuvtIJBfRVn1NxTPQOYC1Dm3S6HJhRM7BFwZ5i5u7Pv8Hbm/n5IQMt9sCfZmmaonAc
2tVDhcUquPixjol+guox45xRjrpfP7S4LWDjCPFoA3pwEAsTVmB/0jmE/kHIYCFsVzV9mO6W5VtD
8bL2D3M2zHHPGW8S9Royfwt+r94w6bAlIkQq3gaY9lUTwaT/fOdJ+Oa4/1mkISQUXbijMwLP26AN
kwrJYKnyIDrhx6+9XjtnhMFXrlTJnI+niNrr8qx0oUXY91KcfXU9f2rfs48hYaihN+rNBRcG+cON
g4FCWAvKo4/O+3N2qUUOXIpojn0BSuK6feu2X70IaZ61UCBX7CLewjygrLBORUigNcFPGHFNymyL
Umw9o8y5POpi5qh7ZK5qvgIUCZUuyehyZiAdugOHfE9TSTOPZrrRT5RgeoI5NDNpprNNVbEEbbX1
vGi10gaX1Wecc7xNhYxsD5LribcZONgq/JgTXPMFC8+q1H0IectZ4Qmh1bOuvN8Qab+aY7gzmYeW
CXITNwGXBrf2sEB0jvU2Zu5N0CDIZJQvicYMLyezHstTFH9HgLyAACMm8VHIOaE0vNw+BfF90kgD
1m2xf5+vd6E9gq1jNTmTsaYmidIY2YiUGPi+nCnqEQoYy5x8/SkdsgRJ9iZ9XHpkU3RvwdGW8ouO
mGWdVpu4ckK4AIIenjKCEWPlQxLFusH7xMTAwZV5Oko+ORZ3gzeon2GlW220Rl4bC/CdsUbRKjPt
EPiJPwBnLX/RELWNPR9siBGNz0txu1stXO0aftqBrEOH3ZL0qyyvdEH80hf94gDOWpD0ibYdku6S
etoxg+6gXKK4z7a9Y6YZcCJFqB5AQ2etO/G23ZOEgqGEeShY7ku9sSMAYcyBL6qBR7H5zB+5cvw4
+zEQqKcFGYTZ3RmXmds1Wi8g0S3rirpq7yJmZCKOxBgLHZwcxXEfdm1nSoNcdNgMfZUx21DMynPi
tGqnmMhqmazaHYM/E9gXZ1y5r0X7cv97ZxWSe3CmyYL54iyy/8CxhC//I92O8ks+0eL32rAtnaod
qtaT2roAkGMxHzi/txVV5nXiGM+C/Uv6146HDeRt93hhC2mg01+rGf+TAH1WxJZoMxBq0PSLwgkA
l+5fgMkmKW3ZJ2WnfJDws3ulmYHwIyqiDSC5AsYKJmsU7+weIDXJK63uSUOjxdnxOUsh9t5rYKkd
ahHJkFK7BnEWHjLh8rNMm01FABVGsMLg+TLXw15qbl6RR0CGWA36tpYLoAMYv9vGdTT1Y2M2NirG
M4brDHqIhWNwTcigOht33OujQnzd4zb6ul0TF7hIuWLabD9+3P/SLK4SA9vLg37JDzEvPQk8Y+B6
Zhll4mw1558WzihG6YYRm14CgvFoW9L8mVcJEayzPrckkhkfqD26qVNuYrINXZJa/t0a6ckMcM1U
oYWgPqOvCYqmDgnkw/TGD2PC1FIiih0O4lfnPL/PiepYjK+JrT/jznlFwTJQQgXgXnbFOQlIGHeS
MkqqDp6W0G4rt4vC2GY8njy6iicLY2BbCTVEfMPQLviIRbjVidOr7htZTfjiOES2H4gu467WwiDL
z/nJwJ+MqscTGNVmelny0CnwePPLwzkutnFrKfCQWyum0YHY1Fy+6briASvMQ2HZ5AdSeDt+Gm18
OVG+l8GIkBmlZcxVAkeOmhuGknFnasZOuC+NAMCClYPm5RPmDwZnihEZrTwSDH1d/s1uliqqvus5
haXfB0TxonKEprxZ6G37iSQq0l1BtGT2StHovzxvUi26VuRYaDAIS8PVpzSEt2wyUqdWS4y7raPb
GsRh9j1x2M4yMQhbZe0MilhtfEGHakz3rPrXQh5XDvUschd171Fg8aXx5BEf7N26NOUZ29+NdDh3
J4H7/q+Vax4/oC+qzPX0SPqq2fRdo4R3sNYCemDlpqxvjlZpBxiej+/wWiA1O7goUd/cBhFKjQHH
FYrnzMhyggSe/hWtC6MtT2/I666okGrAAHPHv+PAM4EcwW7IdYZcFUHavcjynVSjXjXtm7sW2xP1
IVRAeXvco5Z+ocevIEMx8JQ93P/ZO3FW8y+k2o1z7Vc3v8Ln0rKjRDIqlhyxWJs69vBW5bDilKAo
8hWipf5s5AT1PjD+fcSlIFk4pqEeiz/y/ANlmDa84ShlvPnkBnFjD3YA+ieFDdKnyqneJ0Mjbvzm
9vokloWKuWGxz48ja3K5dGm9mzTS8ScKn7yUpdpC+fUSjaKMlBDWL/RozlTux9Ihij1Hbiiwc444
Fa8M64eniczVJAFq9Xk0Kv9fhnc0vLA3Ixrey7BwjCXjHt58mfyebD50l7Q++d/Hnow6/b6LpdvT
7iIdfkpEHlY1euWWy1ZyHw0f1b0hGYNJ0djv6RbXYKql9Up8VHRhV7mXyf3Tbxbx+JniqS2aOMQS
geMLAd9uikD6MWCsji32OD+C2gSJJks1vPvQi2C9zyudOgna6/12+TDx8hrofPf+4UozVDUGFqtV
tjW2b7mYOXASPnE+qh9jTpoIkws/Rc1dLW8s8+ieMl1zwkhxqmpRLtMIWcsZXefBnhkIzolz8J+a
WOT14ywajk8oVZUxUhEKanWTNX/sIAqihSbRoZlobAL1/IzdcTfEJP64kfbzunR++6pKPWO8puOd
TTe5LFR2pXsdxm7o3er8KJO2WSTMBSUThuWI0omyeq9SEX4wRJQseZKnkFGUlhBy0OhrAE0fke44
dsILYuoe02dP79XvA88KTl4KMV20mYinJAWkVIf2hBNJXRIkbNA2TFgyLjGH1WhMwtFzVBhr2mcY
HJKopToS+SQ1KFaJoR4j8lT9XFPM/1a7htSggVPK+GlrbZiaD5tuXMWnkEwGWgaErsQUodFratg3
EkBTgAGCqLPfA99lezeu4nzNP22P5gQMrzJaPYEDU8XVc5wqFiQrlVCs0xFQhK9GjV+8hIDFUpC9
b/ZS3bIOombndkOtJ2JIXhBV7tvJJtr6mcyGXS0twyRum9uRqJc5pZS4eyQXPXV1BWGFkpKqckCg
KV1KD6OGQ6FEbk4eW3y9BrNzFkWdVfLPwBaYzdQXwASMkgApVreMY1JfbPmQA7ZNUE5FGTHj0CJa
BS2N3xARMyimmN2/BH8uMBprDFvGzqNsbS0TTP78eYkF0ZoZM8+uhxlXJKeczDux2NjhOUVxngwg
GKM10/Jm9JnZ2DPQY7KW0vJ9AmsqChZXSMJ7P0LH5mReDpfLh2tgACSFtxJJrleXm8gEmTdc1sCV
IAwu1/xG4BzJDLeACYEhzpsasH836wc6QcIqV2orE3O2DqNme6Hfczd27pt+M4dvfmeat9bCM2Eb
8U0KbK8J16Ucoor2PUY7IV+PIPoPBmMf8vrDgE1Av/ZsleIv4pifvA/ZbUwkf8QIe39MnxxEytbh
aHLffiLD4+09uIfUt77oIxS0gNxpUbaaSPJ0jgN7QtO0BSBNEoq256ntlz7SQl0FS8r7S/eenHXG
W5boMN2VC3ZMexuFmgYdqgc3Fm8N+qDpL+l/GwP6zcPa41X00qAOvZk30w+kwRRKNGkBNtodwsps
ObhmzOJp1Nqkt+fl0P8Zr6/dFxlfRJqD+2IjGaVFPbzT7D33QtEIHDBc0Im7pU9aUWZrcvcnGRTB
hbUXEq+zKWrT/B9N6zbrRk9WJuLBZajLWgVXphnCJCOsjBpy8Yh31K57+4WpMXR+Lpn5Ki5m4m8P
Oh67OGHSeMqSWgKqIKus4V/cbX2q8FgWBZFKvyNxFkKLsNrUDo5xvORbggnOG8pjbCqrLJlAqsvG
WVBpXaxG4PxxDR+Ovs0H5ehFlwqH4NZYF1QIoev3lG7+qj4t+89awaZ886vNXm/Jvw5jJQcEqAiG
v70Gvg1RavTMQqDX45ISMGlwdMKHRnpVnNXKH2ISRkZvrp8Qy6Fw4LqohMlR7y9mpwqERXwvSWHb
7EeEp7mstlw08XfkK3UXjY8bG5y8H+8A1tPIoyt57RXsrhcuwaCfrc+7UA4zKPCE+tm/rktVhyRn
b1WkHmez7N8Il7bbZjTUC3tcvZG5jH+8TIAFSKLg8GHO5lf27RLd+VV55rZrFsZh0CXERc5fAh4o
tXzd5WLU+d7xb4gtRkFU0U6obhddrbtGqInaElzRnHJujgKef7HM+7FGlZyRvCc3lY84cA4kuH+Y
WZgVM21xq3LMdjnheqkhxFD2LnrWWCtLhJrBECw54WBBNvj/shQelEsjkm3SFaaT6pR7xBHNEShL
+lbC6s8/27cgWkz+iTnwjhffWGpgJLLQxX5kZUABKatoaOVnBkOSIcAq3A/AkwWjB3XehuoOOlqW
bMFscz/zxcAP/ZDlC8pc/6JjSipohgJo9R8zTMMsB/TUuVD9Audp2z+DYUXROYvtGwwsg7STFtOs
XnJVkVtIPbzuzAnbiEkguXdDBYvNMIWAomte+D2dmwYodPZSwi1AgMQW7c9GTpr9BB4buV3GQkWq
NZ9yWuAv5l+BNYqct9fChtWG0ezV6J3WJM+EpI3KIHA/rPnoPqhtAUL2yK3LLFnCuBUrvzAyN8Rm
EyPiVltwpXeUfKANyu5NPL5ky/eKsF+x1XUm5kpejP9JoEuywfp0FDJy2EoqvpKE5dLjSZXEYDzJ
bu1l9+apFwZVXZ0gIxqBfeVkeIm4LvHVO2viZbbhr7sOp76HGnMzMYZTPHn0rKoln5+KHSKCyT0B
5P8oyBpPpF1VgBlXc0M95+xQXzgdJyolzUV5Esp1wpR+Q5zff8PUbofBy+HN/SW9mFPN04uX+bTO
OEUeXIGPLIQ1vqMI0J6n8EAqPIA7CElloCp9th4yNO3EV0XWqHtel+SsSI+PE5LodqM+PNu0KSCI
/4Pqab4QV+45GD0b0HcYycshanE61gc7bz0ok55TIENQLYGMS7yTLGpr7UqJNdxqEpKlSC0wQYT7
h/DQe1Fl0PfNDHkX710Tk0PIAyrTjui2Qhhm2Qmnq3Zr8vwS1HvOP96kheBAedoMCgwYQe+dcTT6
5YLEE60uk1fTBgqcBvL2SoLK0mh+u0wYW5MaCQJrWKXscmMLlUJQ92vRp8GGY6hi8u21WavZINBL
ZAgAya+0Z2doIv4HZnn5eqC6Ugj3hWzeJrI+VrO0md/9c+aGK6q+5f8ntQ9JSoO9WCG1hjcOudaD
MsR8igiXUVEf3DC+G8nV3QYOEScXyhynYNaMLpQfUz/+UCnu7L2QlBOKV9JAYh5CyotdCuWGK48J
o9q0VV2VWy3rcQ2nbIvJZvHAxa1LRLwxYvPabMwzJZs7jH2yUs7wnbKP6cUQjVyrxwjkeAbYv8wR
kMjW1NpXmbdPpCrEvosGEMf9CrIO1gywJa0B0HtJvG2vyoPvQTeiKMhkrmxm3q2hpaPLHVhp4T95
akqher1Y/xlXBJfFU8ASG2lc1Ekmis4S/FhgsJrN5HnHL8ktsAJW93Jq96QsxysK3OksVQ3YeoNK
BBSPkV9mzVF8dxnEm2to5UAIP+PEP8MJXghCl4i2xjsqpFoKtJquoBobreW94CY0vRlQ3hEqsXMz
4mk78BJ00sXWyyEbL30NQ0JhoLUdBru+JyF0tA0fyeS+FP6l5exr4MlS+gOvD9+CAqm6qao6TSza
hFOgd/z+FU9n4X5xAH236EnUowPZkoIYIwwZx0sDfiqkQ2SKTLg40wpjt1eyKJIuafnXDEMv1dtq
6KG36cEN+hS9/0XiFnhS6mRZaSgZIXXkJVCJQOzfaMfpLKM9NOso/I0HMaAVbkJwjON+ytD7JM+j
+WoDCm9SJaf4lCuE+rato1N0bGCSKWsorPKYkjLIwiTKyJczL3rsnEBiRHk3owibVasj4DGI+q4Z
mw31DWT9/K4Yia94w7Ipqh4XSDoch4RPfnFVNsTe3mrNRXIKDBM2qqGMHY9xnG1EGLlonTblMbzA
DGBH0738BTGh89qfIs3+i0d3HsfM6ys77lHyZ4/YHtzJ+yt1oTV8awRH0R9oq1Ieezzg8L7pLilV
ctxq7X4kBIYYM8wjiHFotjVYX5QkSZaGN/6hsFzfXVLW+hvr2DTdWhDwVME6SBqChcYWqVDyLES5
dYnaWJtYtvzo0xFiHPlX9YUHwgzM/w7gcjFTXaZ1eLosXbxfiac1/9ASvdTcgLO9VYozwV9U/TlW
+gpu7IYNEhPn7Z21g8otY2EH9iE3NNSJOYP5SXMdzLnW7B8hqDqHzxE+dYkq9CoNjFlGTm3lOj+p
Ak2iLFEellIMSw93evkrHX19cBAi2i4+1cVpuVmZD8Wed5WGaB1nvJfGW/CvUVAlQRvsq1tWlNAm
91LdFVhnUf9jyU5gtG5JuyNSQ07sWgxnOA/o55kKvu0QZlCJ5ADpxbS+UAv+JJLSsAvXtDOrLZ15
8koIUSfGiOILuYohLZyqDXl9cFnANEXdgqDBlo7T2beB409bZ6OiRoz+rlAxQnkR4P0bBf9mGE5U
0aChPCD/ZJ+m1T/MfyEFddutkNODwItJ1bdx/w4FjWiMjke3RnbeVTAuVcYjgwiivcOxAny9Tn1B
5Q04e4lCh7oaZlb6+FrV2VLZQIoXf5ate6jHDNxWIKkct18GvTec+nHxIaBpGeSnqA2sjkIKCfAe
eq+SUKVWNKI3Q5MZlH87IBp2cqnAddg5Wa2KwcSdZr+xqVODQ677XkqjE57YkE7Ol90xvlb8mocg
8VqZ5+r2sxj4SZOwiB4iF6/nootd+gZwmPFTIdHRQtbYClw6lc0Zk2tX67CR6kwkae1sSIZJ6cJb
zYJUqPA3Z14gdY2m7KKqJZo62ll/KSjEWhJhgLAi4c9wBp/9zniPs1CDBLNor7MwZd9/pXZvp2j8
QA5zU66g2Nj0OTEI9rGT6AbwAmLUGQUWcum5bNH5D26EkiIJRpnuSIqFMYBdUCpuVYI6rqIQovgE
3fwkf7BLQNmsUEQILjPZ7gIoSqwdaVo1uV95r8aERpikrtmbT7ptCcgKpXk0ET+3L2wDEeMli/bX
yLJcixRbp14KxvZdZztodu0tS9aqZccoZX0veyg+BRVfU7C9GEHFWhzf3SVMNn8u19EVOXiLso7a
FrbGd+iahdUcIDdvX4Dsq/C1aUr1YupiQIt9kVkHaKnTdwkVBeJIoikDkNpLZ2AG+H+aD505zY9L
metcjG6o0i+TFYKtXu/Vf2h9Ee0JlqVdvDaIDVLzBjpUePExeYohr79Og7Sa2dgxa0RRLRYdw5ir
MxnxWUjblbT8p2HMnXMOW6LGQgCcZAOuAsSJpsJZpR1IhuoVzPRFnRiHFZWh+7ko+Bco9huxFizY
vruKse7tacu/zCDs8ceOnwbvpMlWLvywGCNZJw3ATQ102FDnicP6IgT6fVab5FE9yRjKMF9fs+RA
t5Xdg/91YqvausJveRHhTBkYxCREUZjR+z2+GGUBl5OBhkxhvwwiDYokOUrEuzRiE75b14MWbs+A
0C2Yq2Cb8gVF57dPji0UenBC4cC56XuK0deufUjfyJF7esd5AirZAfo23Bs7yjYfmHrLI1CLRct3
ScGmc0c/ra0teasBc96/yPtPxYSr734mABGWELBkAETWMVTDzb8/eTO2UXMWR5YTtOqTfXGOkvLh
sKslcJwZD9euoC/g/zEMQaNpA8wuyqaZK+c77MrhZGGj5w6pM7+DkhVufCEYD1CK13oR1xPcWdGE
qEm7/vB0YHzUt1aVEvgjmW6knIImEQVzv7zABVlLZdBhDCcGVEdrXNQYSx9lG97BL9UttbGHVNvk
Hesne/IV/fxdszJGGI62JTLWCofjRudbHWlo2GAJooUQo/mwXgbTNnToX2ML9E0CIC1FIbSXEdP6
aQ+ZVuP69+viV48mI2D7sP0h0H4rPfX+/YvKvr05Xgsoa/ibzkfs7RU/8EWQyCfWQIuVNdZ4J4ru
bZdDETma+5W/tYarUY+MG7h9bSSNzDO1vprL0/9kfhWFJKv0n6v2x5pdcETZTIKmDaqWwbGwIjFa
XsY0kcl6p8WIEiBK26MqJHu+cFAKt6MTPxuKjJcDYF+af7X6aIiQDB1fG3fdbSXxoBNl0Int53UD
BtEaNSJr1XnPxKN87/XAFtn2q7EZ5LIuvveG3E2najPhGR7UxI1u8zJtqxakfmAi94/Le8ndElpK
uqwBdRgZToem4mZUYhMhQtH7nb3l9PN3ClqIjYEkABElqcLxUc2JlLOIvb4E/JEJosiyHucSwnKk
tOUgpVj7429FEMAumrGic06ln7MtIeDhxOOvu1osxolLuPUjTljC5liSuwbZDszMcNMepvExi7Nr
bW49JH+sYu6OVoNfrrBiQrnUhRmaSJH1OgcdFJ8vRTk6aXtGlJ7jQepQgSs/Ry5ldEaQgCEYp/hy
a4YOjVOKXzQmZiOaUaRBHEsrAZk228X6FjO3e9baDFzys9rUHmEicXZtsK3UAuMl1Bt0fbhY+fv4
GtmCo4uc17AGrvv0B+D1sW4ChO442VSP0FIRqRFxBhf2aPiWHwU4qPDRVY0JWX0iRY/5d7/H4QSm
c2JjaOFOu0owyEWjQYxEVhrAVWMAL0/bzvTKG4o3nQPgBQKq/WwpCZubVVBYDBYstzTxLSZl0xqr
8mOWOWtl70a+XBa2abi9NWyt3R0bGKL9xbUeVNOWda8JsvifxSmODHT+hfUoQF10Sh37bRGNe90b
pyke4ST+cSqjIk4u05i8hFlGWFeAHJjR0LefGRqLZbG4N3Ybf75XAi83TkHIE2Xa6ZC+WVrxevJV
2wymVyZFzekQd4RnINm+RMiCgkjAJ5+Mj4uKU8PG+LMVwUCQpHyYUoXx6LP35yCZPkc1etuHsj7r
Qe7z+mjp1fmOdQ1iIcUuPkbDL5c+GeSHOZYkTluECp5cogGeP1gND4XyBzOJiVWkBiV7rzCqg3Nr
YMknxUEzU5R3rHLaIwZrhwIy08knNPP0Z1ygHC/fYqfRHRL1dHOpqvHyEEjG34QsBUwVVoU2Te20
Zx78hQxNCZnDR2FCsBzOFqgey2VipwLaYnGVsS5CKT/c2WIIioP8yGyPZuBjTRtmPqCwzkUyAk6M
Yy4YYpHUa9Qrii/vNXge0LY++poeMwriNVwla3sEiL83lDLldPwgRxdx7s2SF7NNasRJvMpOKdb4
AD5AXGLRuiH7NvZZFANHlZAaiWRfe3EVZ/6zl6FcruKhBDiGX/pQpi4rUdOf/ejv9BbriTqrFNOQ
87jXVOX1GQu5Wxn96oEJZ8V0aR28pauRFGuCXRpfEjNdXYi1gI2RIrVHSa0dp+AP1I/lEnjGk+g6
04SD/3y//yjqf1b59X3d0tBfOcZiZbsGh6Mbzc/+b+1wzDqdtFIAAWqVYgHXmLYK3+Y6a9tu6KVu
7g1QRcu6uuO/DIDY/DB0arNlEt25P6vpyQaWYXDbaEdwYqn53WEDZgA6XE1mjh/T0nrvPMG4PyZJ
CB0VzzmOzVyRWolScrmmtRtHMzJeKiadinuA29l2dlbo/Whecm1PMYEySBhAhH4AEovfGN3jto1z
O1wDcTUpBLuENuMgesnY6979Inunv0s3dqzpwI4HjIBIgCPqLvrbgy5y1qGQd1eCRtMrSOJfamX6
i4p/qeIhgTArVoYPvzF9xKzaNqHYCLLXXAY9eOivAcpox9JXDlcfzBrbwHGTdbMzQUuX6n0BXhdR
D756SggCgvyZJFwo93X2/TJd4YOWPpQWA9yIjg3g0kw/2hjvNGlYKCcBhnDWEHIX7AZIbqnt8y7q
ra+lHe18c+RnwB4Sdo0qmRQbqDvl5CwNBIwaOzW3po8C2Y3P1pvQiQJCMX3snW3nF0/nzukJUB19
5D5QQyaaruUAOZyvfJqZV6NhUU6/UHqBfz6ZlmLMNMjEIvcH4C1dKq/u10RXVcsi/4VW0u3NElgz
iEI0SqYAnsm21wpLCZW+Kkej71akZFy+ajb6eNp/xVLHVySOo5t+yxSIOZCv4k4FrELhpnUQaB3H
DPnPRi25LTqy4mII0mjrBbHijDCVtdNbfp2kQ+yKujMGIIZhauOPKwmwS4PU/8CUn/kkYcT7yj39
C1Cgrfqa5+JmQoTI80sTzc5hP8PcxrJgsgZ0QDfpuL26VI+/VmJxsPz1gzNKmSuQgUNww+VV4ADf
M+RR4qScbdi1lJmJj/Cf62WQHukzpB2XFWUEKuDR0P9+or2embENxVc8uya0FjEWeQ7fVBdzflz1
JOPysOcB0XyTKKu2qQp0Xwn5ob54dsrKKHWFSuihfEnvScUcsN+v5FcvjPfohNewaJ8hjWm1y64a
pYEmgUm5hg3JFWoLOBeRFO8es3B8AQXvhVi09rWPm5HMxxpKCPsU9nf3SyfvQwMI9UNDne9tUROE
YrFk1t5qtRRaMfU4fdzq1QCh8jkWGFVrXxxYy4TLGp0qfmud02UjbuyPuNywMecVMR4RJTGtV9yo
DJZcRP6yY8zHz5r3qhb7TlZPPtlMSHnBz9c8bu5w8dsT/ZEWhjxJjVaw1mvtNlvS4rktnH48/pHE
FRee3CF3k/hpI8j1I52Fl0iafCXYiLdYYqunbeDOkscn+6XX9wRp1ZnvXgP5jdtA76+Mp+xYPr6s
eohuA8rY3alos8QRUmPh/w5yeptK2RU1gBSRxa8dp8l8x2yEMVPBmldX8Ny7qdfEqBSYPzEENKs6
xQUPIPUHu2nkZNpiAcrgQoSBqdRPCEHTqU1i1SiV0cL3QmvgN9k/AOSNnocm4Prhxp/o/nsjJe6C
n33aNLusU2H9ksaoHS1sUpmPc/2lAgygSTCvgR1ATwQj2RMTWXMvkUmp2/klCUuHIZxigb+Qb9T7
ubEPzntC8+JjZOjAh17fU+9K3hTZDr/UBP0rc4r9UeYpKES9EVYiqbFgG622vFIPsZPumhzt/F5Y
jO8L7j14VE7x8zOFdHU/XdVYT/oFiIuRfpxRdMrySToEfFVitgqqLyQYrUsS2yxDjPaAZGqDT5+h
0MSwxQxCywKY9pU6ljwqOVFuxcWu/ANNCWFntmRyRPF87lrwxYeXjVzopAwxVKOlXn0yKmWE2mkB
1gjs16vma35nqSrCNAUy4E6dqTSkyDV4A9FGZuDUM5sFdH/Tk2VlfJdWfK29p8L0nIUNlNMuf3Yu
MS8PCPiHnlDClgnh8Bgemr/gSqcKY8A4U6bWpRC04FTKsU0YnlTlJbHfCk4XxKhce0lXmDZyNAIB
c3w64P+pvoWTnF18clyRrpbgjRxGUBT+hM7STmbFAy5e+bCF+w62+ZrcwRT2w/3wEvTbmYoE985N
FwBLQ9CoGCnVtsumN5jMJZK00hVHfmx93Wxmepe9X15nx9XAB/FdJn+IdmkdazUg9ew6vPhvrpN5
IgbWRlpIS4Plub0+zfgGAlknaw0PEPBWyvhhcSB1K8H9wnTDXmKLP0gfo3tCo/za6hT7YB7wavIF
L2b4jbyrgd3llvYV70N8c9iFCWBvkY3bJUofzbPcfUrxngzd6bxXaGalPvz13KyEn9hXK8wvX0AF
gni/J+bq4+8Rk64LUVuQmJVxrSFlMbudvonPttcP+teP4opWYNBmFJyAnEurBGh3XQ5Mz7YkvPxO
LLaepqh9M1vMGofBXj95RGU4MubrIsYXO2rlsGn+jICA17RM7Qx8C5d+s6B3L1cLwIAl082R1l7d
izF42XdwBE+7aH0fOVcFdqY+HOGvfaugbWhNixokWzTN3+aQRTdTftbdR8ezBRhfqH078sWURnDl
RUH+VcThscZR16pDiG3JD/yP7z1UDrz9oV5GCXtRDnRs80qji9nl+v+rVTU4KelfLewdOO198Fqg
k4CQ0noidgB9LyuRZevElr76EQqSMn3c4qziPp/4PQFQiiUC68hD3KumDuV89dArYhRTZzi+vMXy
b/CF7KThgXtaazvUbZ5fbUZKePxtLTTz3VUR+6ZPVGljepbHedsjvDkhaISihJ3641ICpN3cO+VI
5Tv3xTWzuj/x/ul9Wt/Ql6VHjfI/e0kKYBZPcraq+8h3HEbjulpk402QOCjsDpFd8taniy8r1jNw
7bK/P1ADBkvmNdJJRepFDxfPsqe8Cx84CJV7o+vSm/rHsWPi5IxpfIUN/9B4VF9yaTa72dZhx7hc
Jab4TLcBwjP4iEozUZoM0zAeV6FN5vkdMMVdX8J4GyO+yJ9QlH6sbaQNT9Z+mXopLrLnKlKowBCo
AxPGWU7Fcxcu6fwzpXqylZzQ+htxYPfnB69vGD2TOIDr0LEN8Z8S6V3VAElops7sB9vPliYPjnmU
W2jqBBe5r7kwEEjKr8GK1DlXo3zcgM3eryKHXFPPjK53Ok1IfHlJHPzKp6w8rOT8ws8hqLqOmGjs
aPv+6d6U/+Aok+sFLHBzmG76SgUGIpNpmw7T2/opoY2IQdE8wZh3Fioj4ank9hDfkI0poe68JJTf
uRHoaqV26pBe6f1V+0BEn0LRBkGwl0g8+lu2QMH9JEapoNbhEyGXhIjMkx04uVuRZ+Jro5RnFewz
uN7gauRzr9HZg5RTV6zMMuAgXAtvStz3of/yBHmV2LCO5bPICbnkF9e7GxUaVzk3qkGn33BGEpYL
zDcr1rjjUIWBK/clb3nM7H55IJhHNsiinyP1/FzscpLPIq1zHze+28ZR+85Q+0wMsVeeaQaaXX3v
gTktr8+tVt9vr4myJfwp5FE6WE1bQe/g7sPm9cEEjM82K7Ae9DubfRGa9sYEDU8RrTBY4Tw3VMP4
bWabI7xN0brifK5q8f+VbekSENwG6tEt2lDFY1FChbQIEjVg2sGB6FgzyreD/L4Mz4piKog82A3g
Pn4ZpIP6+sO3/EBFFTETyhJcs36dXAXoG3zhtizYAJ7rYQ6DRHGuvTzuFTXqYCzcuKhALi8TyB7Y
WySFg1g8utrcqe3beGXPfFR/0sAjQv1tkSaf2mw8wshEtrxWugo9cWhNL7Fi0MhDBpdWqj739LoE
aRuam6UsoXvE80XYQeUJJU8nestiS2xLRENDqoHjs2LBVh0HpJpKfHMNl6jbi2OGP6QJ9p6KxRmj
ICYowjHLPJT1rjxk9cV74tGyr8iLAKXxxQKKWSLquS4/tLtlDvbq03igKo3E/hVOT7wJd6U73Ymd
Y01ho79TlqwUnhOOrTV56dx0WTVmdSSw7cx5IbhGLJjPD9osKQ+RDyMseQhXkImFu+VmdI99fuO2
RNg5ZIDMV70u1fCaXio49VUU3xelQbNCtAbt8x5YCa+7AUNL+RfopRdq7IBHCBbaflmB1bXAzyFT
5nqROPMUaIlcT0jvqP+xjAjQR0ynH/YTEUNalKfrTX7IRufG+etUMjQwoXVz8lVC1glbavLtMqTi
QiI0pE1pT4aWcN9N1h1TkhFRlEZUbi+EJhfPXiL3Rkioaogk7uo/8roMxldj402iS4z/Dvkv7aY9
9s/xLWqc0MloQfmPRm9ajGfEjHwOYN2JPmsX4Efj24mh8126cuPfuj2CxpyXT+sgLNjowd+HKjVp
pQLyRHjNg6Sx9smPepPmih9fh6pHHR7wNPUzZ273uOmgIIuDBW1Qcvx7DKx7YZ9qfj38gpfn6blW
lB3yHOCkiR8fUUP3ufTUHLoNKll5Ie7IHoZC0QB8Fb20OTuSSIHk9/HhlbZZFnLQgoyCvTXAkzbf
goOIzz/idIYRT2fO8ARJ1N0rK/LUSUtn/+j+qOBifwt/Xn1HRXJhn6hQ29J3uiGUpEZYZA/QWXSm
jfDEi7uWPP/s22HH2GrfxswCfh+CXcYNzhgkfg906L1b9O/RXEWPfJPCkS8cq+EZ/bodggL3VAEg
ZYsLv2VdaceZMovr61ItUg9Ti5BmTEtg+HoinRCWn4G9QVwD12GiSIzMj8aogGPHALAr7mCnmDt2
LxVNKJRqBGb8quG91oIiMZLBDeNWWjgzB7PI5Vpj9m9G78IxEBjATsrII9MuRMJNlxwJXgtRFRQG
G3rH9XzccXP6PCyFG72k4oFPOn8KkB1se5+LkFmDmNz/0JGRMbEcxcNE4Iydxmm/9YTYIdXz5U1E
aZHOIG43TRK1cQJd8QRVp9gR7+ozDBztuqwTWgU/SImZrta2wo/FhYX8PiesLc7I0P7XFXOOWXEL
8c/tfhZERn5aMNPslq+wJ//eoXOTUv3IR8yxE++LgK+QRvllE0a2AqfDrk2zLVS6uymLP2fpD15I
Jaw2XMBKdibsrtod0hb4PEvAh0DyvPi7jFjmOsSJbj06bjHdb77SOwDi4bHInP58OsJC6Ygok/lY
PWJS2JFf3S+bsQ5iXT/tayd0T8jnbKO6Pk/LyMLEhyIXkZ8Fd2JipJhWktbgtdYx9qX3Vk8SMihM
JwQcLOBOHo3L9L0eSPwOzwzqTcTAD0UMcI7+Qc7KqNZd7wxDz2rf3d73u5mqz/VFE5/juNOCV3rl
ZZifh7xqbGHr1O69RvFrAu71PsDfjSLPoHzxczYlZJZV6Fw1du7JHA4L7+juJSvXbZ9wYDiKafXQ
jGZIUbziadHDwPiQ7hK8jh0PDpNvY7JAtYLEWUpAQ4VYwJvVAqIo8jVVa9c3wSTUBryITi+g/cbS
4DcQrTUKESBBG0wePkhMK2iej81TZFIS7wZgh2O/e2CVRvQf98usgHIY+rinWv30vUFKoy1haW1r
N7cykImfB9yZDRSVAehlkekSAdDBcjda0VM2BedFa3HJOOBtw1cIN5AbEstGTjsbYVn4JteXG11Y
MVY08ZvNXedkKfNKeEyE0E/OtZqAxE3R0TG1OBWS8VvLZvDdF/ttxFrXj8NE4U7VzBd0Y9ezwKIM
Yxa8UXLIDr76EXtsdpuNrj14YOySMaXFReB9RB1H1QIv+8VQ5sMnHu3uBilK3suNqtJODwQyWUmX
pTRgkuiKKHMAK49MkdruhuQ8SLk6iNIgOect8QNkCSpcZymArJ56C0ydTOEt6XFJOAcAaY2G9Jil
QBdDq//ZrE4ob9iCvkioPheCg3ViSDVpwjNaiwjro+6jJlBzSecy1YySWwiRl2mivFR5AP9kWTzC
nqQBTbEhKvqBsaq94vJyrpMGr7bDA25uSEpNqb0HFOiXlF1yiRiXlf2yvDwwTddwEUiMGJl4XLho
tuJ9cLHlPvEL3axp+UGaWZvrXv9hc1LqfgBaZxqm13ncpIyXzz9kJrkbJY93ByzIwDjYSjsTuYjE
KTnmKjqjxA3TU0V0FNnNYd2GPRawoaRKMnaaww74anZuYGlqUKWv0wfjJdRRDs99y7HrlvlDyc+6
6ztFL9kTnwCIRKhoppCvrHvT4DreaEBsGgVTy953Gckf8iBYm/WB6BS8lsDDNnFAOaGoba24fzln
ZMHKCFCO4K0XBTUdbsHBxmCi01of8M40udBuPwnOn/8dIxhWYuDz04d6JkY070kl7+ysyiBDzbNn
CONuT2a/QueaFLHgmbH9i/IU1HLc0/yefkuiHUMyBEJ/8UbU2e+IbNAkFv5F7bltyH6dIKMhTyOp
zrp5XM0xoJbqDMIaPHGUVrJte/7DvgrJG+LmK+mNWAWkHekcvxbENlldM+/f/pDBV3loJ9enIh68
UB/OJmxwnmZT3ZMTe2G+TnwOCGuJ0I2wtXnj04YrOZo8Aig49kuOIsyn7fhsI5dm8SSxeqeapVOQ
HknJfWWPPxC4U6S7G+oSATX0GhlZC2qljiAE2yG5vVivcJPt95hIYLG/nQJEDmya/a5yFZ87nWyZ
hjVqxSgtit62VjdpGDLCjYOHNbf8TEhqr34yEHFOsGkTi0GvYJJYf1ySqTJOFMz+tzV6kPi8dBqo
o3RRtQ52yrgN7u7Ortu4BtT5WVvqz92rtJ8wOTOB3li+hR5U88nG+mpKJ9Z3qSkn1KPY49l0ihfk
y8bLQwzrVvZjsGkGSEgUHDPV13BebhG9z6sokPoYu9Z+U4M8+55FiPHUomSZoxb8Eb/QG/PnnrK4
brYIJJ1sMJIfGXS3o5xdG/rIRMajGpWYudG2D/5uT8grV7SUoO26ryfryxPa7DZOhkU6OuzuHXxi
Z9GId9x2OX8E/s2f3ETx/isIUIwzr5HqDu3ex+m0AbE5FBRhwYlQFyOM3v31JlkzvbuqKuiokO6B
8cfd6xb58OaWAeF1zvuJ/0gYennsUvHv7PUbk9tEKZ4nNIWYtVQvUeMbWxgUhyyX65xEnPknFTAJ
FAauyHBZIHhmM74nUOvwnH0gCsxyYPRQ0je9nfXymOceLMv+NqHQfO/kBmVDKuz29Mywmiq0semL
GMpXHXixHtTRmFZ/upxBmzaLjfayx0nlhTN0oBTUe2yy5/yGcrEHRSo1lrI63iDIzudPAgS4aaHD
x/z3LuNBPztxU4TBXeW3gN47mXSWo7PUp/f77aMcx+TW7o4vAVgzhTNYw7qD8vMVQq0bnp89KzHK
ywp+xwF9K8txkUTr81ecGEQE3Tyiz7LhW8kxvFJ7uZ/bDLA1H6WJq1+1Wgg1qdd7WdwArVu3o68w
eMRx/ltpxLIT3O88Tb7xamC+dY5amFqdPdMErrIeGPMMSXqy/s0ztfrXvYyoSjLvuQXdcjQltsgA
L31LyDa1P6v4LC3mWqUh7uO1ez9dJcUmhYjqqCjh3Ve3X6qJOaYQpirqzEpYG2tAQD5dafXXRBef
c/6Z0EsytOz2/1vryIwggCjiKK1erWhsCx96ttRfpxsPUzfI1Dkjv4a3lrYX6GSCXWtPAhOFjxDz
7uxKgxXVDxklr6iKsOdyvP8caa+fkq3KQtx/5bj9WV7K6xbB5lWFNT8qYQHHqgMRTBSh/mNjL8CB
bEIMkj2GB9jPuyzglmUyJwjFf7Zhj12o2ZEdrq7Qb2EBBtKFoPf+10rxFZSAvunReEeUlgUhMzq7
Ioe0P25oSAGAZsUw+46qTBy6P3kTkn6OlcnlGBq0+0oGwRtGR6MG8y2JuRObOBSts6tmjCg6/psp
1BcXHvYl/EFe22A3/VI9kL2nmuqtS14rfRnFO91dY1T0VakOQz8LjhPgIlkAfIh0ZRqOGlpqsTrR
KG1dnXOYayyBkfjUYwSObwF8PTOnaIHZfJUd90Y80Hfbp/w7fABnbQsWcL+5ib2P7iZnbcyBLWtt
d1R0Y6XsGmri4llClzafCPG+gCX9mu1PWkqBtaiK3eoMShuB9cc/M6cPpZTvZm0FiTVQAjuP872M
9pbb11yFYr2uxQt9usB9ZSNw8L8FmENBvCbS/KoSLOHl+EmniL0SerzgNyHycoGkHN3a4kWlJx8Z
9Tdo5pZKYjSjlfkIWlFhXj1TdcMapBJ4hvHDYWUGCaF6RGY7GGgThb32d+nREU0s79RS7RI/On8K
UTbno/vErhUbEvaviV2EkZ6odBY4HKfWd/IEj0/JjDzlL0Qrilnx4k0iszno18JAo+0dgnWRBCsA
TWoCRPiY4erx9XQ24becoLtSJ5UMfEsIujCPHzfO/jqYjhW0HXhrmAR3jaSkgGHUfQbXBym3Yt0W
4n7dN5wvDNG1Up6937a6HkHLTMhtBueoyuIVV7bD/URNUdEuVirL0JPPtvI4a36Ms9fM5sIMkIah
kyIjAbJbJalKApZACTR4eVynehNt6GiXRdMulcJcTk1mpcvFZA/DS3leVkbU+9OcS4NRwpsKMYgI
DWEyIIUioFaNZxl/3s4MvQquQOKc+ynG1GfwYbUWSE1O41L8yRfSHhya3ZC/aUTHXXZAJ9OyAK9u
T5pxkNRABFS/LBN9XRNnQLa/b6M3fMgpXRXZRcIov7OrtDBSOu3rVeG69gl3hjbB0aszsVEBiUku
jvDiCokC5c9Z8LC2wSLI5zi71OlzzeKbwudxs0uD6ndYYYhiQd/tPvTSqMJe0ObNidsOYuWAN/bS
EHrzDf0CQml15miveCLvYJiIy42a3LwdNzRv05wK6W/49J7gLpO2X4FZ5T4lFi65/BhwNqLbacEj
+lU/DDVzUjFbecJhNyzr67UH4Qns7dT2nBHKThmqJjdahX424C/PtopjhhYJOEnIoJosyUU+eVcW
etdNgtR2hPB/dx6tFYKGtVIYHPKAlzYxAAefhrz8UON3Vu5a+spHbGnuzBCA9nngM3AhLeFcMSjE
v5XgYy7JMZ72I0KRJQooEScTdzysRiKqXz130DQ89TCUurw7e5Zg0Sm7T0pwmckkVU174ULPMUcr
CqO91uSYUvffVNk0l+bWKeWM5MEoKF016xGFVXkLcoA0XVQhWCa5ADOJ/G79G6QH51biB06ooak8
Cpn2sPpI49MSPnfNANTOmxdKiwI+IxAGNsXgBi8TaPXvTXfoedq7Of+qso1BVIFgh8oSr+V0dDWc
cDkHGL5NTP6x9wTcbZL1/G57+xlV4/aI43mnfZryBGGczwz4AoX8B1SRmYFT9xjnAFNDFia79Vay
u0I8i+1ilKplHGMfuyrPNfSjIW5RhCO0CijVwIx/ceE+zOfe5oWPRmLLg/+khpkEJ7ifgt8aU7ao
ADOMiTVSReKsaQjjVMdhCdQ4HG/ua+G15G/y9PkZuesSiLQ6alwZnZHBku22xOhs4gHQcqRsVc3+
z0Rn5mDkeAaLM+z5foRBvYCxXbbdQNHoLbtadQNYx92iRMlY98d1vwKpXqHEGCjHzbvfyBObB7/U
2YxTdJKRjr5EIZpOIBs1OTF3NZJdJS0mSz63LIngbyfzJmGpbc18SJhrCfEZ2TZeVvnm1U6oYEke
866M70qirgGCgtNbs9wYh3YYN+vqFBPJQK4SqL2ORM48n57demvTg1tW6yhg8M4sds218hBamBPn
uPndyi9MF1AOO4ykIU5oqjIh6q/MZIAWGHXn1/TO+4HRlkLzLxm7XPVhlJ4xPJLJw4H288BWU1pA
h4AuKv63F+5BBCRVt2LVFDNdTN6IHbArMo8J9QCuH93ZSYYAdQWr99hAl4aBw85WXYbjlNK8jS2c
oNP36s9uBp23F0oYpOFksepQ9GYntioS17hLMi/HpffclxYCL7tqyR0RKlILe9HmO3P5D4ZLF7S7
fP/BLl64Qc36b0LnN94ixdZcQOE3s91Eai+y7weNyIc0aBJICBCt4HIcQ3b1LWgAUxDDtN22XhZD
c0+857CWFi92iF9nvJ2WBW7DHka5JVkMNmYZB3XA022aBUd0S/ZwoxETjno0XzR0jISK0UQtN6Ti
dAcN9KxLQxemuWAJ+A89DYpof5hRo/a/crVszf/VMlKlWGaAxUwxQmVD9uD0yXOAJx57RNEIDrDE
WYVijGhTCT3X+cQwLHfmW/OpcxB92C8lEnKdhBfr4Ve+q2pMgRvfZTNnmaSyOr0Lyk3RDrvKiKnz
BX0L6l5lgo9uJKyYnQziVAf9twVntzV6RJ94eqIytly84X0SweE+hX5t2NTCllTmppCVi6WUZnCC
I2G7Oijm4f+eahQ0TPdV1hos8WxmmbXuprNAblEXCfEAz14bye+jy6AGLlnANJ6ISCJJCzxx5qUO
zPHzgsERg1lFYqC23TdINOihFDJNB7zNGABsGrr0yeyRsMEIp1j5ViJ2VmeS4gj/Zl/x4xFiUov6
2i8b9bA85ERyOwF6ytCaSO8zvh8+exz9vvqsvnN8sZsJtlJDNnIye2Shdsj/oCz5wWnWstVaFBTq
Ta/vRr9kazj8cQot64Sp14euEt2JvS7CW+PuFRfKGKPBuENevK7MByfctSdrKML+htsapYWFF9+V
0vtDmVkYMTFlo+Tj0HceI3fTMpA7CrjCh9xfjQtlIqGKP+sTLaHvtQiwc/IlmotbcPceT+KnifHF
Y07cLRmLPiV70xsn1fSSBaUT6+meO/Yx67rR7vly5QQQrQNEYovrbTSOZqK1Y/ovfahcnou00AcL
NswUVY8XIPRhQLxLDqtxVDVDtm+sXxHtsCjbGPfb37D8/aLfZxc/wPt3bawYlbkLzuaMdVI2dXXF
S9Bs3Mh1/wElVWslVvsqpwQfaZqDp0zq0O1sMAN8WoxhCPHcERJzlH5zyRQgqbgfUtFWGLTtTcLP
5yElUmdfTEi3LGnN51vFtIzOLdt22YPwJWOoeVFHNgWg5qxQ8fXiCAkhr0NBPx3Vyi+H0khzqQbY
zK+DxyZbMRgWxRsUJUs1wWXRhtUvTJD5hVmY79vXotK6mYJJWHdHENtKIK+7pTlq/Duwq0sIGQ4k
Yl4HDp2QWnWt9S84nPmtLe+3ZB028KaWzGbLtCr1sA4kZhzHcythm+LRCuW9UFBTrags+vedOw9q
X7zzD3/KdZFkwmOypdlhf1Zteh+QOJKspiLAVDMJ7V+i8fkcsrtILAehKtDQapresrOixBNi+78y
Sg19++gUZJdx2sKdIRfNy8cOEneDyDW8LjAmne9jeki9OuWb+LNdbqZ5BXLZ+WoDqjn7nZKXoB02
bKFzJFwzd/meyRCBZeII5fR49afudLJEFaEL3xX7+gLrkl6wFTbVb/YbY+C8T1qP6E+dEGWWEZkA
CAP7/AWWDGsS11Pd76nh3SKWBD3ex4VCvs2uo4ewUGz9gyrihT2Tf1vjl4/W8cMcXN71ZkUjpYzF
vmPlpBGj9XeSH4hdWBZbOtNNs6QY0Ip172x01ttQlaZivV7IoQAOVo+ndUOjbvVNEidROkrB5cYU
40vG9hg3nQLk+W3PmI/aw7FXnaJOk2wFg773+qmzpTCM+XFu2Bp85hMAGIkJS6zLXBOrwcwlPgp1
zZAnLIumoDEUofY1JxZ6QpSChGuH8ZpoFDrbF7N8nezYflZIZ4KvOjFpsHiZIbdY/0a3tRdieCR3
3X0mQV0pxy/uKy4UyRmmTNKhWALS5Fp3yv7b3h4S0UjKgbEDlznm7ncWqp4Qme2nw2/nNE8KE2mo
BmQS5QRG/Sr4KOiyMsNVumARMRIOh8sEeSmWA85gS33OFg7YKKRwUHXvxBRdRlNjBejuGV311jSa
N1UX9PrqzJMI3nPrE8J8ipoeeeEFZ+VG2YusFkXOuxKqa4mhXZhtoZnc3wqBglOC/v600H4m3ROP
kWIhQro4Vw45wHkUMPJRiMfCD4p0p6htJF9adPb6VntdZSxW63z85dMqk33JiEFR+jEe/IQAw5lx
WxIWJSDvdq2WSd36FrQKefNBN3zFPigCUtSW1uOa1YGf+W4titvI/XVAy/yrwRFXfknGddd6+Qxr
1rA33qex2rUeeuZZ7GKSYDCzoJ+t25128KtCpb0zCfJAyZO6c8UrtKhGfv1d7gku43zaCRdMvlFD
fXs+xNG3Jp7Xg51IcW6obGV+aEX9Q5GhsHwVFl3DOksmTvgaLd1LV2N+sAx3lRa5nEjpzPy4X8cG
G6ZqV7KqZIkKCoquwl/HoPxG7dMD/vBAWKAnXub3epnKmh+JdyKmRteejz3luNMuXeE0xWoyYjym
PCGyXbPdYYFHnbyjrSPLJJLMk4T85HlPbNqIcnh3g6l8J1xAi2tCSAOBb48faGppOoUFgNb9Sa1k
+tBIUSHD6fahy02sYgfB204HolB1YfgkT4a1SxGJqFscFMvFY5TZEvnbnGc1lcB2uupj+lvRB0Pc
zOurIBj/wDABUTqw2+Yuwt12kYf/BXbvpsOVJibrIoWgrH9mEDx6pwoKXQy88i34wjstDbURz99k
K0s2I/400RxaSgkRZQ3mmR7uBxWDxVlQeh5VaJoIBBhrTg1pjvaFl386oexG4bFV8yt75GPOFA+w
NIecWOhutDXT+q2odAG2VUdEmekt4J1mmKqRk8g7g6dcd4LU5tlz+3kiR5hvX1XVFQXbbbf+JU83
KaF5PfDO3B/eeRBO2V3sB5pDFhqcgzeHmj0n22I4sDgvsksWgsTmNBmLYkuxfKpf29ymV46spzAz
NMapy6hGPm2mGVGjjBwJ/Ppzhu2bVgYDrq+CWBdBJH1EaOEueLJuAIJw5AGmKW0VmloaZ0WbJNsT
Zcygu2K3GSBhryGClXNnRugQCSwmbknwLIoDwVItJEcLVOVhrEiNrxPl4zZlxJICbmOr0EUcY+k6
1vjbYmv8HKTNiza8f0dPICbGSm2/z/qohXQyBQ1LewqAgOX+N1+Q3vTjCwvV6L0doLLcFq7KnW9A
yzB+FHEaMkaKZWXHAZY55cHA3IlSF0vGl+rx9UnLWQLKp8AaVfTvUnwO5Y4V6bwpjW1pgV/r29Z/
n3faqbg7Sk7KsjP5eE1116mc9FwszuyXNyLo07XSISj2yVHW6sM0cacZ3YVZi9mkxeopU2Uom5jk
lc9A9HVdNQeN/lQ9wGCl3SetxEVsj91blK7u2eYwM306YroR8XFYNjAEr2Iuzpr4MwjWi1loN5sA
UtDK78GlOS1tDcvuAzDOzda+Ksf6VGGpk8Mx375HlAU+o6A4JOdrAuPbZD9RmJXTd7mHi3Vp2tr2
FSC+/nGvQuEcndP5icJSwSackm/Z3SUuffI9MnSH1SdrYtJklw2gKJ3mwUHh5SxXhCB0HD/sLYtt
OgQBaN6fh0tzTKoWbfNhMHYlmAczcbo+cxSjid8ln9pZ9T2STlry1tN6TAacNSM7VXRBKdBUcvpl
t0BfiUGwd60ckyUYY1D29GBIV9TrHOMJ4OQm/PWmxJAwFK130oqPQG9BYv0tx09iFQS9ckaJhhJk
TCiiGXkdUAb+MOGoanRb1cCh0WEUsrKmDSqD74B0yaXL0bqja99l4FXHfRJV1W8kovUajLyHeKBH
ZlJDhmLsD8xkJ7/TKd93O9OZVHPnW9cnoq8zYOgjh6ISdXun3seXCZ7K4K4SLzXD+VMMlPFKXEH+
ltuHIuQIwuFG3a57+Jh9RuvG0deIPk6+cZFlD6+BLx44k9g07FY81EfV55NT7RRpNv06BtO3qc32
Jq2iAwEVUt7/IgqAKpY1UEj2/wTrOFNubHEMSsStv/wRmSo8W5ELeEYRd/42sA6zyoSVaOdNaWBi
p/Z0MX8CUGt9qHaUk0eJJUiGedX/3bJgXjw3K9hKDjcoTowUd347KD06Uh4wip4cRqVhuYorkEzZ
pn2rypHO8/rZM2VEBhCAdiZChNKWJ0rGE23cIAm+4m+bdsExKU2QKSMcBsUDt0jSUUlfBX1vXOCM
dPmgU1PbEG6DA+4jyThjaMf+tAm4NRVRbtk5HnYEMynJGS6Zfk8jZiYUG2HRloXp4kLEkJGSlo5e
1Gn7h4n1ACXdI3smqvWNOi2atQx/pa6nOd817N69totvPjN36VmHH1RP7Ji8TJs8FM3WJgfZj9dh
kH+bHE57QnGsTNyswKjfyE4VDBrZvx1T5LPBiLL+4GpjOHWHYrXy15gK3SM9dxKqgMNPL5Dx4QN8
Q2cPgYkt+z3+ajugoMsz4bUot/hCyuUO6gMi1HHg/iFTl9nXc8JygAYzfXScLN7BB5AQ5MRRYDm2
je86N1gojWYUnEJkgv+pULL5b4QEgaKaS+koM3+10C9rHYCi0e/HaA7bMy557yYyppgnkUzxy0Bc
tdvmbA+qXN6yogJSeOJXDt14BgYlsHmOFNnNhhBM4rU9g0zqgt3UcLZz20ceSxrpON8+y8a8pPb4
vCHL/hkQ+8yseerxpWniVB4d0Iqp3mhxK/12QwRh8r7UVJ98/THdYP+o+NMop8qGK3Gp5yUhix/S
YgpyvknJf1Zc/TAyTliadM2/0Hi8narbCU2m0quaJ4NeheHGc6LU9P/Zuu4T+MwbmzTgeg0VKOak
gsWYQIaTpk5GoRzzXF0DYMnoU1tB9/70VnTlPlWJYeqbVhTlCm8woqzlXyju+FDGrI/vPIk/5Q2o
eNJHBJNxXCWruNcdT8DfoIJ5/KYRiLnkafopavmPzm7qUR3PZ1YmBlzn3WT5GCY4xuP4+MzC7hNa
BH66UuGtfeBQmgkWxliqcJQUvZTwoHt+iUgzJd7Hq1CAWUCDArl0aJ24BsAkcmjohsnWfEztVAZt
ZR5qI10+B7TLGP52jx9uruYpORbxfcGFmrQQN5xuwbs3vaDB1C4VYn/SqFTGMiknId8Q8yI2llau
oGmnQXWOJJBwSMaw6H/rctBLlnbbUh+2nkdd3sjEn6v62QyQGLPp7PKDbaBEAYI9cczQ3VQios23
dLMEma+DAAhhNafVAIPUQwFKbvBrXwW5Gn9hcRp39SLnRvmPMf67Y5fx9YCWT9/rF6gLPuHAAU6H
O5e85Ux4zy2eAgLBrRxODGdmjVw9YI47BfcEhTgmFWS1ynMOrLKQcosSe2dGh5ReHX/uRbitZCeY
JsNLELohidB6l1RkxevIsRmIKp/tT5HZ9LkK9i6y3S6RoCMAipXGPvKZwmpbOQ0y29nCaIKQdMbN
r1X2FNsPCbaUYnklvL6ofj2XbNpJnIUlMrEdDoKMr7uCF/kAFxsE3To/TztW/5eQZItEPSM2hA/y
JSjdqgU8D3JYL5NqpE40XYhomJi5dobIbAoa7KshmXs0DiXRWOkNBzqt724pbcB6AMbhZc3pHmqc
nu/FL3DEK49Z1o63KCAKlS7/oM/MYfAmLXmUxU3imBC72GxdO5Vmb9QY1Fr/WK4sMF69QS/rumOO
tjwsT9p5ATxSqmM5Wm1VACq7zhz08tMw8aDVm799GD61llwL1DYq3EE/yyAoRIz9jyFeqXFv0mCh
RB0n59AojyKaKA39CfhiVMLMRiwedWQj8zG9narnOGWu6HGZ+qbWhSwbDiDI9Sp6iTlnzwNNBrjR
/GNWk2ytAq7Vo5TbNPjHFIujPsNjyN8ZDUeG+h1xLv7txh/geJaviTq4F9OaDdco9aGcfiUGxPYf
gxWgEv0nEZCeMtIcJeIxFotzKr4MMEogSLve4bj22rlw5WXVMmQWv31hk++NKj91Ww51Q0qDgZI9
6kOyYwyJNT34h5BuWS/VXt8is9ZQfb8AFXH1Yp43OUYekR5bbLawYr91dvnCGuq6yAMh+5NZlajJ
cQGBYG6TcwuEyySWAHKuIMsrtZNwuptvF5t8VcIzdv54NZq0azd3QLKDumdEqeRfBWtRW8Si3my4
5E3HQiwLvPfx8+kyTPBualqTE93kmitY8BsQcaKdKc6W4sDNbNGlwbvQ5qiyboLUlB6rdguC4inv
elXcUr8leQU2Lf1jSLUM4CzglNpuTEiALUtH9xV/CKK9TLxyXunHPBMFvHxLXVgk5LCbXz0K9mN0
W9ExXjxo6HPnkStkrC/3bk451UBpF3iJgETDQB6LufmDv6TGEJxfLiYUt7t5vTeNrhtVO0pbHm2b
54hF8s59uzYPFUn0BwGQbE/4nYzxTLnOcXzIXtPqy5zymHlnq2SNzpSvm+Dbtnx7vMe/XOm3yDQI
6Vp0BQeTykkD8ofHTPyUD4BB+tPs0V0aFHDsL4kJ4ywn/j5sj37ZwA7dHSnhVEq9b/6hQrJST7ed
UZFyvj27/4PHCSZYYh/+7JuY3doEhTXIETJ6WsL8DRMw0TSdZqZRvZ+0U+vKRE+6UHvsIsCE0W47
7mzs+3A7tQ2Z12HmqF2TN0XHzzxfMSXoENR+e8ilYKpCas7DH5mr4kzp/BHJAilU6Zgy1mBkKYdE
M4OTsI+UIlhDt6LOsObZqLYWHZ73pvCE4sYiE2AhEjHW70tes+7zrKba5e5Kymk6XuC1rWbPxqEs
s6pa2866P1Jtk7A6dZAnyLafRPAYjnlVT5SQvt0wjvspuu4HVLn4Yym8U9fQJoEMo7ZnjuoNbwAa
+Co9coHYQtvB/BpfbocrqYoghZHzjoADvOBIFamoyVeO6nTCvzdGt/GrQGOPqG0nnoaYqbGAtCxq
bn6kHlYuRmSgWLeOcvmC7RwWHsU09cMGVn9IGLxaztaQb3XYSHxSdBAR2A9yAM0nqQBtnqdboqyB
514WOtNOECCAJRwyLGtQjw23LFjXtgZD6u4nM4uLrYeXhejdtXnWmyypVsNn/KsWRGx9Dqhmf4QO
PegiLZMJ2CLoq59/fPwOK95tsW/E4KF2I3wBnfaDcv9t8Yn3fGvnYxZnmTtnFwmFYl10mNb71sQy
k5aOjVxUK/g58fwzreG/2pCFYVnxuXhM0tORieu16Mo3KHr9KEt12+NlliEJP154nP5J0cNnuuPo
xinQNLdbN9VhR+FUlhmH193VoUAt+7A6KG/gUuwJ5PX2m+OlUQ2IgJ3Tde521ErrQtld2kavhKml
RT4D/+cS+Gj9D8GUp6egZlhR6yrki72KH4m2Rl7H1lja2cBu9msuOkd2f8/5CZOjc0CUqw0NBt5G
ayN3kS3p2Rch03mk4WQPPW12K1rv3fc/sQnQeB0Io9Sa4Jt56nEbU829bT1+3lD9VgzTXfbX4ZU7
LJUYYcF2lNS48N7Zz2FMCJiZsjpSGBKEklrceIkALs2ATOOXt/btBdJBFL8aiZo7+ERGtIxw4sgk
ayLTafWGC6ZE/0kdotXKn1do0k0CUEFdDC16P72WwNEzki/NRKPwbfmPZVeYS6LV+YzSRuQ00akL
jBZtU+qXbGReS1lGt/+XcqbY/FvZjFt1Q2yqwTw+WeLRQV89ye5uDbaL+8jQnJWLN0Zc1KfwIrqi
yWrpA3al8kBU7upFJwnHfnqlvMEvLNn2K6V7C4PaFKvFlV8x9XZ7za7tLuudLsMfiLhiV3nAXPA3
mvtPDt/63pmQgENoYS5sOHZ3pVVhpkbqbxPAG3rqqj+UVqgdS+dW711S1RTfyQ9ix5el9rD/Pgl2
h4rz+kUj6nj+Hv42rQloz71XxeEUGbs0GH8+5dsQbMxePyn+5Q2UCTEKf57ZuuJMF3811oSkihLL
EEWBF25tkkNfErfRveRR4HqiBVcRjzoNJBKOTxLWwBpegU7Lpz48DICitTBm6IueH/nXIq3JVq6x
ao00FpGxhJrWNce1VK/vCheXk2MxwAmW/h5+7vfZJAHsOe3+ElmLaQx6sv6QsDbeWFC4ZlsxwLQV
O7TgLcITFy/J2AbpqyuxUJkfQU/kZ1LNET1/pDavfHxxM6STSN7hkOEJ2fTNh7QWNF9JKkAhy6JN
rPFu9uPUtN+45QLDt4m9qbeiMtXDb8Zo/rbnejvUcXMJNuSuk/RjwYvMma08XNWJivTBZVc3nZsv
T2uAn4mBr7LMcMRSS/82YV4susc2il0cndCRllsvsvvcBUk+L1MIbvS2gt/Y7Pz7qSxG1EZlOe9G
X7OcVkDWYuqpzk0EvmFc5o2wDIQzssdp8fPkobkc9DVxToaz5et25B2ZZJiVeW7evlZ8wbTpv4ZF
zcuIep4sZVfNsLQyWYBAY8rBNuEWhswBtAw6z+SKV8ycB5PkQaHHL44XIO+vjJKuWUb3i9QHZ9u9
vgW0dOSKtMierCi8TYhqKIAVq2hMwg+cLAjfIZQxSjJGcHKmiDvB9eFl7/U4rSG8Rel2dfHXQaQs
pifVsabAt6dWdolZxqf7pS3CfSjKfnRN2cQNc4IKVXkxin2aQLxIVsnCFaFMIROhpGmOxTNGu2lK
DkldOZrbjbk9G7/7jHNQCYvuoeuPTmeC5h8e3c2SKDztmI8D+rWzmgc2gm0f1y3iAVUS7UF+KYmh
4AAD8wosAC3tNHxgAHfiWOYCUEhqg/zwSaF9TaSQOgqDIVPFgGHfmVAan0m25gYyECeKTDeZabJI
HQaa/cON3wxtkbs6fnW6522LbM49ONsa6L6hm2qhUBdL6Ftzqec4JgbXlZ95huRhy9RtA2kaaH9J
20yEZCRBojc4+eF7lwgPCPIfCE+N7BvYiznlQVYdvN0ZvgEHoxqH8SEJZtpli5qi69f5PMWP+F2A
3rruNYOUwPAhWILAz4f4WGCgS7IolTnfVzTOO3onbRUftxryGzu+5QG1FlBWW5wggSbmEmdVWra9
+sD0LEyX52FiMwl0SSRmpRenpClUUiLkvuqHIPDphqiVpb4X9C+2DeWZK289DouQrViT8H459vTI
vf5eYJOI45hS9yUN9mrxPfeglY1RLBch0Bj5HtLgxJk+EXZAzUsuYa342SA/lGhpxy7AnW8Dp5tw
ISpbUd4kxmhSgrTWqwx6jiUAhYGUk99jXVhOeG9JhcbiN3qcAjkBLvxs7s4KcY5JLocI8FBf+P9D
hRo1LxJEMuosdJVo/1vgmaSKQ3nn7jM69hOY59CXbUpZZ7NEMj9FopWGfkjmam5l1/CsCBDfSLzn
Kdzu9v11Ra2vItKd0jjb1r5/ZNWT+BaPdPhVCrxr4fMdPVxJxAzt49z5GTsD+KhutEt/+IbZcziC
ZEAEYkc3LBmx5q1e7UWPXbMZtjJ4t/1ToNziVfhzyk0NexkyqMGgjeUoBJgdQ6If06DVx8Sl0MGM
4MMpVb518D1uPSShBTCqKfcjl1yLFfGUvhFubd9paBT673VCCgHgLrYtNb90neP2+gX4r20JwYtO
C1ewWJCwaAQiu3hBXEhEGwrtmgIExMU/SdinQKHV+n2zPKPN17cq74btjitA08UjVdrTBczh/bKa
/TZZX+SujjnTFqozglOCdMpihJ2uJtckUQvqSGMp9f3hfVbwa/Ld0Yw8wJb/mr18aRdnTDgDdwin
Yh3zf6UiuFfG5BEoqWKBC1qOR0DCFxNcePNo6tjAxTHfFWyECy/PjPcWxq6yMIEa5V1wJvnngVvs
DiIEHd2pcfgl7ZHl/COt2BodqIIS1xpXeTl8Lc0DctkHEkX4+kumCt2vlGUkZNl9ry0OV/dgMlpm
Qvgsiz3P20rgPJsV+LoHRUxu9qKGKnkcooJsfQjAn9EO1E9yJ81DpvnPkSJA3UcynXbjIZN1OJh8
H+2oOZ6LAnDmn791JNVaxe7kvckI/q29yDUykxysSCi5cn0kRQ5NrXf9yh/KMrhjMB7CApEhCS6Z
VN4qHZdGx6Qe+2gRBdvTBfDwlZ+1Nm8rxtb8jvWKMFcMk3pvzt/ZRQIkdisSFXyAfIpKdAYr73Bd
Xo6/goul/Orr6DeDTrTdBetUifHmx8Eu1kwMzjZsviQbXvZBuCuALY/0ttMXgYKkiP1YwmBWHEKK
m3QSqmfyB4TObBSdFaMaHpE4Yss5faZqZ5Ze0efKvk54vKFZ8QpDph7oQkZGcNUyzW+pzsuFJvp7
sb6CBOG3Pp5uFw/EP3kHIafVqnxYHAIRz6E6Q+YUsIWUw5EBLPFNbDN0banwfihWnoLl0YOV+So9
sdDgADbU9AJP7heZLVBMeQjCDhkgkqiXexvVtY2jup9KQx5Kh80Bfu15GkzrrdyG4c2eswyu3jN8
AG3h+qLOq459jrj6vLkERpqzxsM7E03WoMQX3/NurX6/94WCYDKMEZa3ZYzugf/7LPmi341VuSAX
tRMBp4oI2v3qWBxJ+IZ1cDgSiDAg3dAxnyEV9FA6LfetwCGjR+SMAMUbrqp8b+xtw2i+s6zCwXeZ
Be4H0WCIwi+Y0oZVMw7I6y8tZM2xpKaZCecLauUfMTmz6zgFGvKa4vvMOuwMqpu3+olZ1iidilYW
YvdWWCClOGcx615So/Ia1jOy8QlmxcsJPhwQ6fjJdyGPNYZr2HDxGyax7cw6WLmHZ6mcB3d2Yi74
bvAJjVaFiXZLMxkLtieIdv23hIkH3urjrWbdx3OuphUgDH7rV9W9YRo3DESoynuB20mhUd6KTbN/
10rxHYQb6hBNwM7d3cI9HGkYJKT8OBXhOLRVcnA99qrgVJuGtgFk/UXWnRSs0zOuiACs7pqMm7UK
7uhtuVDr3V4XPbylPgTg9YaN/u2yBgY/KqBaP0qZfFa8Ac3XxZeHpzLvYMKpDfvgt9zCqMdyLGXL
HN1qzf5xAXh3ygzMM4AdHT/b/xOJP4rYBebLroTGZNbjQcYZTMska9ZkXjKrmTGpS/+ehDVhnPcc
40KwrV8eBetU4jp7ATaAUAHXYkrl/7cpOmfSnWET2dlN3RLdgmj1t7sQDyoaI3CKvQ0XppUmRCw+
JX14/x17/tghdGMqPb8GjaRdtlYul8OJqX77eUPDU5bSbQdSO6+/IWtwvk/boiiyT9cDHPc5cW/X
RF+v83a8PqdDf78rcZmj3/Bg4aIHh5sRvYWNIEaXzKhksGeVGsNm6Vdhnn5V2LBPqyUx105GiVM4
ZLhBdYsEE9XhumP3bpiGEk2C1fZolTrmF1md0VdlwtsRu7ZvIu/8T/RajZZ054jeD5/Kwu1pqsS3
GhItBy1FpX7FIacfm5/acd/fjRy5SJKy9fMMKdPhUHCC54s1fnp0GnhufwiklNIk9ECc76Dbe4/W
oZUAnMF2MFben36EpDvtKJLKwsFboXXb+a6Ru8rKaulYG5fxhiouDH5776G2wkvUCMK8bjbDPCrl
D7hcyhLbG2KSQQtDClPeR9RzEJATkrqcceEXoauK02w69K6WhCX080mjRGD2atO9ZgaTsEyhgQ8C
2q6Yb6Ww22tPqAwPT5ecRSVsPTA4gKQp6LKRv2r4a10IK8QInh9Yps8K7qTmNG5WV1yWmH67nDUL
gVdPRmuYpegEA4Ky/jgfv/y4P3XKYN4NrgNiRa9T7cXjg5AxxCXmMwlwZr5ov9Eb7scDVT17jUKY
Iw81gl4fU7BFeueEjRFrPPYxhM29+3Xx/U2QI2EmPZ6RU+lrTwrcSRTOlukWcvbuIJJBtwyF6NvA
YfctT6kSEOJ2OnEGGZ+Ch3bG1xBKcYkvj4w60NTMnqviXcQ0gW6KilagEXiDGMDfrkAB0jxAht6y
Q7dJBPlVu0Bbkxxzb0G5QbdmEzv/zsUX/l357L3hRJVwibNpIOGInUcmOEUP6kiba0IZIpdZMwVt
PTXRiBktJNI6ZBa3PCI/U2FPawKrIj2K9kwFO9fNhEMTgNd1NWdEqqq9msG4Hnk0HEDKGx0cTUB2
4cXxgJf2oHk/oKNZL2zjgcQSxRuyLmxCfabyrFCOzjbUMknxmVZxv4QhqwCwSYEWrz3ncEf6eNAb
cvVHZhs7RTnrWzC+b8TpIVC+wCpaL+SSUaIj2P5YNTTe1sZxShGV3vgChOjSLgmBg4WLgOmQJfcV
CQMJFwvIA1ituViIML8KGH/ixk1zUE1gpoz0Z73JC3XAZ06hbCUQoFdTlVfj/jL7W09xssFMEUst
RZEP6H060LRJW3B68tIWLanKisWnZus8Wi/ONng+Qxe0B2vk4JGkDpBE7RRr/WRrR151/pjUVV88
b03L3nzR1MwzKgjHLgDZbedFDs9TWUWKRDh+XyF4xa7UrT3MgKHtp5DGDIc78KM6lZT59dxHO5Rb
JRNhrKDO0xI4SdWQVdSvFWyHkZ3gVDSEDsEDrRTRGkB1hB6eh2cI1txnGJHlKdA59Q2Tn5kXCAZp
zykTV9Vx1jjx1hxkrSGoiucrz53Xgeqj3QI73GA/HhOV89lAWVBf8gXSMgGsx/bS98gmOVcKe7+S
gafU8l7M+yPIAxY6lJ0LpJq73WyrRm6DRyaVuLTcBL3gVAr+YWTbTYukT0/gViSIk3fn1lPCI7vk
My/Rl1ZGUWDli0FvBiEfjGakQhxJotsD+TPCGnR3UawwGqNYgsiixEsCECQbam/GzwAut4RUthKd
Ox+hsRy/X4mchkegoUzKwc0VLkUJ8n77JycGIjpTg+5nnD27m1Y02trFOHtL9W5oDfiezph18EOo
eUO9HsgczIeNrN+rPilU1/RKVYiJhHjHgUoVlbgkX68RATeOTBawVlFiYzZS8xg8fQztTyAAH3+d
nJrplQrTi8qOKmOhiCiuw7Gad7ULro40H5NItl6ZlfwUCTVc5GU1QY9qmzKMDRKMFCXEqlDGaG/L
RQpxTvtwyAk5FzFQUnrdPlILkEN9lXEDnYRZroEgluKwaaAITxYdNPNtW819ReO+ePSvbzNqrrV9
uogc4eWGxx6S1PwwnnVQGes7mBbYOk0yO/Bd1F5WSpkoZ1BlmmS0hatsLsY8Aw2JL+V95ia5ONcJ
Wl+BU1zQWQk/PeMtnpAzWWqq0JIlyTULDqyZuryf76mUbAGivk5pHdbt/iu+N6cj1oGH9hoZ6Rzm
CQZinizWngo3UGnWVXWhAHtGC0hhxdHiAMhvFPHw8cNlQE4KbNL7D2utNWww9H6/JuKQdCaGHJ/M
gIP8R7tAP7gNC1B3HZfF6WPwWNjxFzlU4MTtz0pMLrHjpuMmxOJVzev7IKXeZhXzaWjgsCwwRMPT
IGPy0KZ168BVspm3PkYDMpFsc9F4KhhMz9v+NxGVn7ns8OrlBCZTl0dGiqkCiq2Hifkm9ZnkP2is
ggNDIu/WXIplSIhwvsR2iiCUJc1luz6qpx2pAAvzTthm9PDf2/h+s/nYOSFcLQ9hzUuQp86L9kwz
DGOZ9pwi1qYrBnknpcE1dHlykfrKf1Cyo8GMN9ESbNr+LvKUbNdoXKeETqanbWapWbIAP+C2wkIy
pMqJC8uDdQ3ihRn4GFUziLLOSukzWUasv+6JuPTjwLWTWGNj+F5AkEDRujc2Qnq07IZiO8pf0wX+
D7slbGB8bGacI2GP0uy+RNmSj5x02MI3czfwuNSBGGWZy+/JTdKE9rELSpK5wLPQ8vyGnSHXV2k1
nmqaoM4qsqKqQiJwqnTxpbGxkbbFORN/RUIAHUMwXqcNl+PBufC1sxXA5Q3t+MRpTEBmw6dde9oD
CPgJBmVYgVRRvNneYsagqYNOeqXlvQK6N/0gR+h37BoF7NoN6Aw+Z8xjQNp1waeFJKPPwr7Ml4HB
0uanrmKwtEJGj/0pfpkvfSVz1WYSynXXLVoKf3Y22k/g3OtSHrqnyeBRtVaQlJ6WKdMgzAHMonAP
SeFgQeyl0QyamRn9dVZc7Xo2Rnt67Zn8+B2aHO7auIt+jl0A8CoAPRBfH3EGxZPPw6dxyiUZLHj7
9FU2GPbaHSTTRmk/9vAvLvccd4T1Zrxqtp+2rrfZw9vHwjJI15U3Z68+zIGRTLnEo5+A8LshtsL3
TCHCSsIzxvMuhDpQh8evLO7B102q7Ic/K2VFyjXKn/Pfdzmdr3Cxzi9cSwA7HulD+rPTTrkD744y
LDdSL9KzGWyucuZIlabLEIFnXH6SMLAYMuR9bzXgJ3CYH+6WXpKnCojSwkemYc9Y5g4S5k+YQpc7
wdkgrv/GSsBdVA0wXiIqwGEUoQCsOQEqXN69LdZBz44273cX2BJwOhHqOl7v310mA3l9P3mJmvmP
Cslcsdd8QKk1gSqJKF1sTjTb1GV/HbkBz8fLtQ/e6O+wS85gt0HdAOYV5VZfcNbbz2UdWduJUl4U
EfqPwaJAV1q5eCCclvcOMKQWgp+CYWJpEJ3WNNCFEJTloFK3Yw27FSegUW0v4BuVdF/3tkxz0TaA
ulBtJhD13Ys8f5JIOrbE13Lxj6sIPfbgd3Hqyx3FRfoEk2nXWRtUMimIM4YbVejGCUpc2lQPa+cA
eK2pndqKkRWerjJlaiXbdXlEdAvzibiDVewmljwnlNV+XCR+wsnIlCcxE4vmUO4/AkEQspD4W0in
pDMu2fSlrNZUaVRDkHPM2TP1khnIdllJtCVDyHmPNf0iGCjB/kHwTsjHV4ft5Wwl3xO8CuPJw/Wu
gbfUhiavVN7a/JhMPFcgLBYHuY+gPX3IqN9HM82cP9Pken1uZ7EPQFRuueIa+WcSeXBzuYg7I/W1
vGV7WjF9KCPZGHgjLQDY0efSfBYW8q2rFQcDfstx68m9w/QJPdaQ069Zza8NLB06lSdMGHCgKpru
/Lmp0LvXP8pQcXtciZmx6s7pzlnQUhzrsBdmv20Ic++a1oGv+hVr148ZQ7fl4eIyqaQ20EaLCT6t
HnoNWYmG2nyI6mNelnWY0RNuI9cW6J9hAiXLd3qskKzU8fDlABDVIM9TgxmNzu5nn1aIt435BJG+
+cHNKsziTd+TNti1vbUwfYqLmsWSBt7xXgtISxCfjtadXi/Nt+4L5YJ1EhWtJvFEM4fFXQ1AcMxj
CtuktFyOiNni1QUzI0gfgLlD/OI5o8Quap7aFAidOcj1cWXvBxNEe5r8ixscbF35IiHQFfW2ibCy
+c+8sjgz+VimyCXth51FIUpLgTgk4zMwgw569ap5c4I52851jP0+r7SxUDb0vgwhi7zv14vvjc0P
ZwcYygOfQOXUnOVQbTAdnOt9lvkcPw27Gwk/dbJsGbJb7lFfdXWQohAVFicd148eR/swTbe9l+bk
5C1ho4EjfM5TBfDJI5KiZmBhx46s0C9HNY5kj5fRLUQVd1iAVol9PKc3C/zyfxpnFeTgJmzROszs
4Cw8xJ5vUXxPyFSxQn8YJChzY7kORAVWenAK8pV0qD7Pv1HR9/q52IOKsbCbsd3bQ6RjskczmmI8
2zt6J0u654wSLEr/hNaUfyaNraD94NhtkM4VFtRL6JEUM+KSqGmppFWFhtfcJ9BNBtFNm2F1YWMy
HsLiVqofT/hhxKQIv3SfCCtih0PxBFjNcXUBW+wFxzzO9Lj7WcYtSh4pPP+pCoZAoJOwAafnsHNY
Qw03FmRCmnDxv/Q/quafcOOVDPWjdfGwFz23zd6vh2EqYnknA/TRepVBjx+GVtmrIpIN9cbWTH6l
aZCxpa4awtOL9ZofdLmPAceZPErT96uyJWC0As2FMxUCsZDFxo1mJtPR13w9nDBrqq9Bst6lGU8C
eu3xEbwMOqu55chI7OMH+EPhme66cGFyO9z/ldXI579XYw9qOajP6rnHdU6IQUTH5otCfGRH3RV3
8XVWHTJLw8s2jt1mev1FIxRHvcM47+4a3ZaQe3xoFHn403wZtG3DBmrOGSrDcAZdoP+VigLG18bl
Pn9NA91rKPsTMAaSnHezO6oit2RcI9BPpx1PyWVuIYM/994yoirjsdx/AWmlhf1UQ0yvx5fdu9Nw
UXzuFST2zUDDJpXS5ujws5jXT4VNflcnAg8V5zHfR9YZT2KatWoVhUl3EPV59F+P7raokUUAKU5Q
hFweq3pwroFN8bNm96tTKgi2Br+0BQJSUZUGg4fYiUinG911SHx7RzNcNHWeDhcsW2cloPmCXOi/
O8VkAdldy03HQbYJ8VDFIWUpJfwJguCaRPV6lQwayeF/GYBp7955aOSZr4oOORL0p4eJfbGV4L0e
sy0FUSbEcTOGTbpwSQvctTjrHeZKtWOsxu3BqeneLbLXk4y+mB880fK390k+p7mHI2qxaUoeKvkB
vn6Y7yW4ajmUzy7P05acg/HoBYLQ2uo0OIGnX6Fh9adHYtj5g2x2+kW+bS4IAPNaLDMCsXyXasyi
kJIs1GXZP6xtfDUi3eak7ysDnXehkRPNbtx7axwZoHyZvT57ds10Q284dgOKCZmZEzXT6/lsxvlK
o0GGDmqhZq8SLDLL6m+3qwfRmkYiDGPodRaXpVmePsflnSo0jwegH8ToRZZpYFG+baAiNqhZJCho
VrDAJKQhPptp8PY+Ho7VjY6HcMR6LAjVv/PViCANpqngPMZHdX7VohYUexDtkNXwZ07PXEqnOR88
X60DGGG6tXJWYdtTC3vU2nMdt0NzRrY6rHBqE4/UOwX/9+DPU/tBm9anaPDdUzScj4uPpUc8OtQD
Y6JI3y3t8WOpR6eB0tOp5+g9skOG1kc9qUiIvPyt8W5RhXgUVsLVR526EG2NyFOBxK7d6xWKLlGV
/AfjYD7YV979WLv2GK8DBkkUqB2QyCu0R1GOD/TpekvwyzclCVahqLH7s0tjTi3A+9J6RD5aqFxm
bT7rP0Eyp4R+V0rI4Xq/o3DiINZc9wpolbU7HM25RfRgNYp63eFX2h/mcZAViCsuC3M500kRuZcH
bMCKStdAdMKyzOKgWrFgouCU8BJwzBi7+BDWzrvKZkiCQm9r4M7sAU4oXU6XCgt4kVcFpcOrxSiY
4fk90h12TwGQR6sblwRYtmGVCo9d1j9dZ8l3I6tFtKfo1mDbyE7fD3CK77ZZxj1mS552N1BUaV2m
KMDegabKYH7vqgMNu9byhOCmCKAby4VRJ7Og4fmj48Mkaj0u6LP2X/BJ9Vfk9y5D2ydqZiVLCDs8
HP5cifv++R+GjKfhf2l5v+Ys1WnHcg7AYBulhJT/WrO1dnndC8PO59JDUbCk3WXSb0ogJXABSxwD
7OjvvBLpUKq0CVJrK/gdvxbNWksqFyHu7b3yg6LfaQl1epDthaJs/NfF2cbMg2hOej5yWoUC5lCg
uXO+ZSgttKLFpHg2I4Ggo/7mZdF+Kx0baZAB6m2lK6BM5WRIfFj1y5vdUKYhIO6bjFA0uXthBTR/
1qjqwixW01DBcuRUbBG4JwiVz3jxW3AO6X7AaNoZHamkGyDW32LguRufN36PnKkU/FGTOfq14ib3
pyb5trEnICGmMAgZeAIlJvW1oqcoBUDF+f5j7njepOO8eavHh9ijigI7GOqiuI1LShw/5R/DwPsn
J8UG2kBaZ4JHxmDFMJnNV4ndbfOhISvxz4mm/WQ95rfhxAhmVZ++n8YW3UfTZ9xY5D8NXAbUvB0L
dZ0SWnU6WmBJ+38/ompKxDmeXM4lnXaYtiNbBfUxE232yCwYVmWBZnPY0u+xI94rXvTJlbBWZ+LE
ig02yHaFL0zxkKc50IOTY3A8Tvqnbu5fdHauA3FG0Yh7hp8vSATalwragWp6+37hRQGikAPs5LW/
1ijMpqnr6CQBiFqeJQbtdVXqNPSNfhkdGCia6+aa8n4rICvABSZb1Ryr+XD5/v8hSAx4jqKs/qSM
c2qAPqU4CKIdlU3Befmc+yxw437mKefozV1xC8cZVzHWMdfvrAd/UJPmSDZe6usxht7w1L6LU06A
JEqeq1CdozG3F+VIyDLki1eIm4EKZxlLXHQ0RST6MkeoksDTxwVi07/6DTSK5/M7xhTdWEdJHtWn
gGlJ9zt8jBsKP6G3f1UVp7yVF3qFzQI3+q9r65aMLObso0/wYtSXS83tw0jp6qMCmASB3sZo2UmM
bXPDV1kLwKPqHVK+whzTN9sPu30D//TWlBjqdXMEEjIF3iLCcV68PzbDKyWKbble35e2JvUEnpdJ
ySghqAQ1kn1AEgFQEugL7tUxDo4Rvg/CpTHlOcBgUjGYpS7OhpFbPRuw3Ymm1X5waIDXPg8xFVV+
Q6mi1jG5bZ/ZvvQ1WRBvawgBZSAKCrhTmk9e95Uwr61jkXHlVcecuopKSwsap25v2VpKwUINZHTc
cTgWrMwj/AA00MVSJcmNa2Jj7oIrapYt7X7QDgXirEfrIKy2a8/3JtiFxFmYiMDlH5X1OxM8dDEt
7lLdy8u0vo2P4R8V52hNOl28L7aSENiNAk8Cky750BZh9YYTxRqzT2uvjxBdtK2EYYIZapjbSz8k
+nRLp+Jva7FHXgzqmaL/5399DvACEVUdIWthwTSVGk5Rsv4lwrq8zakyC0ouokfyqTXscARLJqFJ
Zmqd+9ULlnTPvL+2UQt8rSabjG/F4PBfI6/7kXdXnF00n28umL/gEJMJNQb9XPpvgZl6XuZkInza
QqBVfP0g+ev+kfSTYbsHBKkmn+KlzXlxbLjY1y0f6rYhviRaPzWP0KBQlJNEcef3GusOO1fA5Mv7
MJHKx1VbU0lBD3ntMYVzoQc4skw8tkYCPZ4NbMdWsmxePUTuteUSU05ayX2AUQ3F6sbHS9ABcSZb
3LkPWUUeU88VqlE6R+pVZAiVyHu/zVI0kednpvbn0qHzDIXvKh4IBQhB+DOebAAcExDWgPMrwok8
6CPDbg4pviMcdQv6GJHsTZfqfC5wDqFJouPx69yqqSBo22VrVbq3W4C/FlUHali6qc4DJaH0qK6q
JmSU7sm7ad+yV+jTXxW8nNLO8ESKq/vXFGYpmqEJ+0Ryr8ZyFueordEp155Cil7D8vHxRX5U1j+r
B38TA5Zgye8L0EJBCCR8CRUoaRT+MKjiTdlXlQ+L8CfWVPa/+gEVi4bXxNoo4ZcTJ8PXORdBrFn2
wNdXqo/hT20txcLVtJOQv6qR4m1RX9g+wemT6mg4Kw5PZi07oozfH5MVPYV6P3UzW5GdmBRxZxYY
SB4qwJEFLrK4gCgvCSLRP1mouZ9HchXtMyZ7tFeoGWlt8jE6FDSynEuwfO2yAyyNuh7enlrjWjwW
/TKxXvKe1CWr2pB9qbjdV2V446numZ5Fb2DHM5FnotitlYWDTTCfax1njyDA/yLW2R9mGvv7k4mf
SX9k04cjRUOLQMBhRvOXVDCdyZ+auCknzWYX6i64JpCwpVujhKUhoMZDjc9xbfRmd61jq53yDkG+
R+70xGqW5sVOG/f89gLiJVe0tlt1/Jf75Kh5uAmr4uRJYI8LQ8l6rx4WS+g79RlyAH5cEuDBsLnU
SJu1m97UlVvL+ML91xuc/fTLU2lqZSl+IV40yz7bnLLBtZ5Haz7CfpcxaLzO8Uh7He5GjLI0GaZS
Y9GM3ZaV7/spOEdImwSnl1PIW+66oOlsXRMRggq8qndRIxn0FI/ILimp4vvNdgmLCKK4gRHySH6P
uXvTkWjPdFTBrfW3vRZxLGfviC8C9rX5qG4bsbE+OLGAou7TqaK63Chm6mcM6dZBGpbUfCwMPmEu
fJsMzdbPq6lL1bixj8nfEuwZigIwkTV7BPdksQ7fsxHlfp8UiHsfXYkDl2q8YVkyHwGCibA3kQtc
3qSLcKpfPI3FzzeyGYrxGJQOYZxw0Ep5AjZW1uov4KX9EAdgG6HeY9e/yHcnPAUuWlr71xsCMptS
T6dTpa55l9juKXqYR4hrsfdN/nZVpBtAuIZkbxmFkzXXwONIG5mt6/t2iWPyBisoLvHJBaoAUqkE
m2ZSG5+YU4FQlhSJ084RHsY30oNW2ZExp9nAJAwUmITB2grTCTuJD/+fUUXXGBjciCwC5gYvguup
WIbRv7KWWofZDWRv9xDivQGA2yhg3BHB3rdq8sdIk1ODwKu/yJ+l3xljWUD/hK4Y7dZe/83NNwU9
dOUxSzEN8uzzUAZT5s+VGSkPOYRA3YT71oZCGiQyCUMEqT/n8w/+hdSERPVzvHYzzAG93AvrsTmQ
M9N7hlPqV3Px1BFF2rE1/E7ZMVBbzkIbrAfmjtUXG/d79yHO9qpJ+WpiUxQvaaOGfplGl9XoJvQh
8LGJ20ENP+KpDf0tRrFAACDDH+F5totOhP8Qy2fse4gUZjG+ADHfCczRWjd2c7inRX84yO0e6z3g
0zAGVhLO1Znlsm2Pn1rdXU+MP7+JSCSpFdmK3yRsUD2Dq60+1IkSplIIZa2/yryw6LAGG1WZHW1Z
bdlthgyso/Xee3UgNrUN4uPPo5BFho1P6aJWha4GTf/DBFD1Av3wtORBuLWmfwOPg8rjUkyP8eEQ
xJkfw2e5Lsde/gM484prF5OmVNHbNBRD9xf24OwereVFRqyrbGf8eN6Fu1mNbbCYVtJAjLt9RjJs
hz10M6YPDmQvDu2oJPTO3m7h/rfqPzlbpRnUtQ0RN8cq+cGa9X8O7a5ih10P6OKgGEgtPdpdIZoC
6XXUt12Uw2FQWLWMhDot/H28cWlqJt/zuYlrSotmdi+KBinCxbKwDZXguaFsCxfEpf+wu+EaK058
ZjQxv3OG5osrX52QLThAq5jzeKpwP4yn9mockR8g+eSEbBFLk4aDBBqh6c21n11i5p4hAXPjIZiG
WF0aBLSiOwlDk+kmDLX1gBn+nGoaNR5Deao107h5K8qzfjk4tea8s99Qih8B3ob2lbhFCpowncDm
Cg3u9q6BzO84u1gWFULRj9PlCSZSex+TWR99exMukpyX2HECDzcQp74gHwPGukJvyWIEUTDIvLdk
uudTRV0fCh/7PMwqUlMomMiMnL3Z1OJP+v/YesltNdJmvbptBoexok4Lr7ChhOEMqdsdEl1o4ba/
3OyYmxGm0iFph4APLLTMnRCzsyo4u3NJPb8lXccMeK3goGClejDjabDmM6CNCyD0w4/gCQKaJojr
7rYHGM1f7Cra/TtMkOqFyXUWfbGuNcXTvtz+DXX1iwm+BkXOA9XcPEBA2VWIi62c03PO91w42a/Z
59xS3Mh3O/eKMa1z+lWkD+wwOMs1GcwCjV9zQ2MQS1wjRTywVUToNKCmr1O8HA1sSKeRN2sGV3pU
pds4fTZNZu3QPNZaylSnx/8j0Tm1VHMug4EDuXPlZR0dTd99RVC0p+EEm1TjOUl+BvFvco4SkQGB
Q/jlKNyaEsR5nM6jOH2OF9mMGljuAW/fIA1C25xDdXWwcmi/5jKHi7OPhIuIQY/6A1Z+YX6Pzzsw
PBg1gWUZGa/K89f84PcveQMRS844mUofcKsvv1t7H6bI/eSa3DtQdhIOUlpAUfIp51vBI9xIdE2d
qRDaBNDOfFr1qdre463bK3PukymdyYW4gzruxl5vRhU/ue9YwNeFQEsJgEwAy7sGpivfzNh3fl/9
jFr/Iaf+zSiWQwz+5+c9oHB+zaKpqbYKi7xBkmwL3lT0BWwVLCUIEm2mjLJ/Dbez5u+bcWw0U8i4
QAQbqknNmS58yDYEB2n6mlbk5o6JBw6cWrQJrsq4Nu+fMh19gKYVdCE7Ikls55B63hMR0A295Pgg
ZxT84zmabq54SN/NgALkmO9T4u0/3/2IWQ5HeuYSFAvnGd04DnGPIDqoQYgDxBfYzmZLTj+/ZVgx
vvAo/V19T0mdYVUuSrCxHYPWKDLIsonPK6suDxcQykPVlomPf7xGXrZ8ihvxW1jJh5A8tNltODLt
p7m/5zQCSOkK82I6z7l6vukBLJpu+JcblH2WebvxQjL5rq71r1BuAEn9mHosggYE9fvuTmRbQpO7
yQKIK7PhIVvAxjAoEcf8mDBj2iC34ZA6NRnomhGWEHdsnOYcaoaG7U4rpxrqxQZ5IU4y/WyFfDFs
kAo96IIiKFlplhcTjN/6stRIwSMcoL1NQKk8wq2x0g+2Wo0MLZZUS0DOlY4IXqCEjNoovoCtNt5b
zfhAihl+zgu8SRF+7SbG7T9aHVkxonmsiVNgI8+PERDJCKjU3R+HRdVgnazoReawerCjGs9fy/pJ
jSCIGMEDeg78wZdr0Apo7x9AHc3+u4bfe+OThqzfktGJIPiqyQvxPlpkKYQPaaaJL7OyHxvnySVn
ROv+7ydwpGR2+TtNy6EAL7zVX+kMLoUSGvqX+VI4kuMX8yr+Ql1wuL6k4X+ipzpmKmCJWgKCooVI
wMr/erVA4T7K2l+uGMlQuxPQ43RmFvCvfFcEUuhqOAtDau0leRrnLJ8BTEtAKC+nZuzt2pT4Lq1K
wBipQWNzTucvZX2AEtxGdUomrjJWGlZ0i6BoucGyLublN6977Opx1gWJ7lzxzvitOCe8joIc1DQv
TRxGXoWc+J+teZeMP92syxRWXMIHOOLgPuZglEUrxriD2gf48np7kMDI0SKLrqAQxNB35PVyHJ0I
10Le5rHZjT7d/8KvxkANMh+3c1K9Ldw+Qo2bYOBfxehU0LvwHUmx2MscSBDy+3fHsL4bjojcWEgq
7CpvaoUay4cjnOZ9MzXtdmE48Bn0iKfbSYIf8VPPeGuish8drNaWRLUbvOH33hUGdHcCbzGR6f3N
NIyiVP/jHDBc1qc3gr6cY4js+YcdHxuNyBKREvjgBVfbNpa266z7vlWsCARBaUAKyDXrgNMCEm3K
KDlJ+Cj26XArwDx5FJKznmoT18YkFW1V1PAwcVuOEdJeA+W58ZNnRDO02/ojyC6q6G2fBWvWmmQN
eji1A5fNUth2BD2HZERWDPLRoZNLV64xohaT/F1KN8NS/XkxBw7zJSO3bxNLijsjrngsZbzDvrZW
kNO9lyTRLLcWQF6R3NH/x7AtdgY7nkCVXqb130agIDJokmY3s1BSqSTZP48kylX3q3udklEJ9+JG
e9xZAB2fXnoicbiTTvub3n67dlxwKuGz49hwdBaQ3Z1ldEiPmUCIGsXRAtGNh4Ma+c7pqpwzD7kP
jJ7NkaIGhyBBxlY/QX7W+MjnvLyFVkUmZTFJcJWsB3xNeRnNJ11noG5ATaulwHnlGd7PX3tDyKee
FcbPrS2E20LesoBpf2LKMlbHovlgqCjHzhlLZOv6dzYsOH4YugmtiL2uhCO+ojGvQNVluiUempOD
E1CBZy+2y13GUA+Rga0GBrjyj+ECfSzUE7C6IDA+4yObyv3J15X1cvVbTEnKzePxPWM0icO5uUhE
Z2uHQJS3Tg5aaX4qaUgF0pBXunCtSJXdEQYe0toVddYkxToTDhWp8pfgEDfqzNFoXJvbwkF/z7rk
WnS7VAr+gjo/3iov/IfSbuQhxQAjHR73kJNIsgb/DPcfnvfrLDbZvNW7EcEpxNOvO08rdiKHcfEk
5SkNKbK4qxMvAGz4e7yfxalMWpZ10aOOeVCB+ZLKmQXWfh2beeCsI08Pft0JbA/L+fhOG0LGG5er
VIkrDSA3cEcMNtMdBiBr/6q/x0K/4YZTd7YHcFGXjOt3azoUiB+cdBZroua+qNwTMKIRxDG3qXVl
ABVRhtgsJVdfmsbLqEo2HP2JNhA3OzM7oA4Im0sT6ufd3YLUkk6gGj3rPY3nlTbbeaFl0uE65w7I
lX0n7w+HDl+Yuc922RF3BcSX7XRD0WRawIk5lXUQyWpV284csfoMwDMW0qMKirrEdxw2y8X8NyWw
M3Pj3cQzIqwfqQDDgKHzTXA+zxPjxhvG5a0JQDLwDW3hIctMfl0JV7iRss0iVFDSv8JiF4eK+nu6
XSc6B6JE4UAj9xWYgNC+aSsryIyK0pvorEUoWgb7WMFEPeN56AJ/Rf2OfmHgXA93GyKisIWcihCd
KwRGUF+5Ta3I0CZS7DUGBPCFRs0Z7KPzXOo9SA12jteY4eHD44WHTJgEuntvyeMaOYEsVl3sU6u7
PKUikTl87NiZszHjFU4lK+cFyKlizgdCxpFZ+lKfLOwmUs68nZvRAbwuucHidajVUYKBDJuZGpge
keoXoRHelb6NB5PB7a+sNaBrdSIn8HJsK83WiywWLpheNdjoV/ylat9z1d/9+UZ19LiQKFopeVZI
iajJO2k0owEXUyo3BwS2ZIEk8uhau1kKK/EH0lhlh+NZ7qM4AGxJA+DUn/sO21e7y19QE3wWDnn9
wKpQSPuloxliXURJjUDbUN8CRf9rtjHwi0BBs4eA4VEtiDhrft4BcQVQie03+xLN3qtPmGUiV84i
jla7yhFg5HaiDD7m0mgyxzjjQvTcWFJO4rrG3a2SkNeqCgFtbfTBUtVhRwDSCl33C8yp2J4QkTlm
rcpUqlS+Hm3MTcee35OtqRsODSl5Jgx/rQ0wGbEEkhKMrAyiyC6vK3qYPSBGEewa0CmXjAc8THJo
IPrWifU9XXay/Vz2wqShN3ddqXASKM66VdVdEce0ULW3oLGzIrQkvxBrOo1nJwDHACQtNXRd6pnL
hjlf3LrAfRmOClSTqHLLeVA6YCYhXviPxPRtjYZsB+M+CmOuqQIj+hAsU0iCRUmqdlJL8+vxYAiB
cTu8ySyW1fZ725Un/RNS00iSPmk/YBrV/etGoXtiWDNnmC0A+ksN1+2K1MKRh/bm1qZeCoyCSC0L
BmJPIAumJhAHXv653WTupHkGolqAawhrYr/gKELIYEi70PYNUUGfjwP/MjhPqjOSIoA4H4XZ6QOe
8LKvRzzuvgdjHdnQnaYC1wBOmy3vBJF/2pLNOFBDA0gQ4fAKk8nxut3IqYd0OJqj+9Byn4iip9VG
nIS1fNNOjaBuzCvSB500EI/KOrC6nY1POogIj+G9+qh5RrzKdObbGuqUouipRhLiG5sLeXYrWBzk
keiplnry/xltOtqH6Wv1RVDVocw9RXQ4IXkaagNtOBVdYZxQhZHTGOu1zWyt3qzCEzLf/olyxKLv
HV9xbLYK+uc/iFfQ9Xft/edO5TkHOjzKDQrcNJPCQ9OzA3BXXYeSrq3PXqFQm792BfhCbeWYGYv1
l7J/3GB03O4vVesC2Ojla2kF7tkx8vY2s1oUVLwcCvlap9EPWmtwF4WCv2HfecQeHLXZhOCZLESh
Cp8hnuIh9rAphddQ0XibC8DYnRmpzFwCWAb7afaMcYxTNwnDFuypaiwmquxVTSGT8RMSpt+dA9kI
5NLU/r6Jg+Fam/pCd3rRLtJ3UOgE4wRjllnnHTQB5RZnz9IkA+mlVhl0UUgghkmRo6alQRLw0zpu
K2qCf/pLj2gD9hAhpiI9tN0/FF7o8+OTeqW1g9RoEnYLT2UyUJ47TauU48YJO4CXPp/fuHATr1+Q
YBxH+zTWNAtI1Qr4uIz4f4ZghA58wYz9/ZzLJjQ5xaSHjDtIoGZMxRJol+QqL4T+tlRDJEceKmF0
VV+I3buV8JVU/1sVqEad2GQbR4MSVMIrUPd+yANTmaEzGLWPPea0z3B3M8jk0SWG9p9BC3XjhPIk
3cG7F7wl/rkvqcDCroTXHYr8i3+jTayLETgYXhbu/tNry9VvALoZCjCx5zVBAVeIp1lQ6GvR48AD
oNFeZrgf9gQIUY+hDnk/ZXrCENrjPW44XGznELQ4DKwua85UZFs9bm9yDSqwC5kHX5QItlv8cAt6
WIiqR4TNVHpdSea1stZOE4ZlyUzOWLZUJ/YB7otgY5zdJmusvYrr5/CZz0sRHTEwOriKZ5i2p1fJ
bIcvUFbMuYghXJ2BmcVhl86tyBOIsqJwqZ5zXiAz20Zw/u5DuFlpB/RNHqQgQHuths0oAJIU2PBV
s+50nAM3Zp1fttieAHh3SzaGwxE4H78AQ84J957mIyyf01Nqx4XXVRZO0S/UFKNbmrQOKp9gCXuo
YAxSuR0g8FWSguojJFlHAykcLOg9Ecav9EGYHXutz+K5JFvliCACnHaFxenAtU8mdgIi9WDLS9NJ
QtPRClPO/Ro3kBPe2nCi5HU/E1cRFnfGPXIXrs2gb3nMSYhPSJMmVsooF5ci8K+MxZIoyIekdG8/
Hbtfhf2rT4BydcUlG9uWCXvCoCMETg1OrWncT+96WnEiU4ipRqfaniB6JzwyYi00ENWmftMPvqsN
xPi7zEt005sMpNwoUR0LVNIWbPpSAGLjd2OH3MoexWdh92/ZmxT53h7YFXjA2dWwVfvXcZhpymUg
lKbQT1ByGiecVp8J+zAkAvZB7+cmDjJYyXUxVZmjWuQOf2ITvs57iGaKy/y1hI0A4smai2ci9W3q
5GJtB5u2QqCVhPrvE+5k/WguK47tTM5mfqM49TgAjoZZ+PFyNIPHdIxkv55lfonpFJVZoqBIgmL1
XN/OiGCoALNJiJ3oHQRzYqf5/BJwZNTyqVJtZPm/ZzyCWnDptGcvrvpBrETKmZGSbMurHMTr8Uxd
rsOPv6hojNDROGJh02+i0TBXAA9R3jyriLwSrpKouw9dK4a9QWq3/7x3YEsuGQhqBujogVA6sxGa
QpebF8DkY6R/C+IsPKPauK2rWdvfiT7FpeE11/m3qI0XQpg5AIOrSoPcDMMDZy36bjDgUUTsRDLz
xcXkB1AWuzOvYuBAi2MNs1oGrx7L38jZGgCGe3WQB9c1EZTCqCwOwdm7+ufVmO67qN9z4DH+KxO1
RNDrQrFBUBQ0fWmgztPZDeGW/WTSfb1daFlAxpyYRPNa4vvoN1ibI/9OQAD8gGLra2dde9UAoyou
brjg71WAyJZCm4zlLFtrKiJ4/z+G8rbfvzqY8pXu07tQDVjCAGT+FmDJGu6SYuPhLTVak5G6ZQre
WkmFHq4+7rKiXkP93c8iyWZGYujDdjegROFJS13RAhaTB4r+wpBBfMzDp7DLBxQTMD6n2PHo2XJF
00yJfFiJ9iLqngOfyNy2XIA1cipDC77E96z0PEihCDXyCY/r6ww2AURP6NcqS6Qu4wiw8WlFMv5V
JX46MskZwlirNL9o6s9b2B8vP6I1/WfdGhQHf+8MiCOg5VEmSHVzfTeSdTFhbNBKHFePYfZ4MVAa
Jv9GljyhGkl07bkzSfqbWX5b8twvcMIbLpYiThEP31ymjB9zI29pdl/4ryy1G/6eCQKm5ifDAo/0
hFq6STToNSKdYNilAmVIl6gUrotWl5TiDJU+z0pbmL4pkCR4elHZb2O122ognNykcMmSHo8nizQA
eSZqhHuyB0wTvMcxaOU6hOFj9YJkFnZ/JTl1M6OJHDFekIHMl31122jGhE+DrkYmXoHLobs+ODJ3
+lS+GYK9zUf0yTr1AB3ms4v1I80mWjxw3Bur3uO4whx+WPaP7sPBB0PETKsShALiNEgkeNhJcQsr
yfsA+jajNbPeHXIBUl38IEVO+cEWFhwKGZ7Z2xg5r9avxfRnYKweGvt3YOry3acsi8lGAKAwvajX
wG6YpnDGmElNCcAkCv1nVcPdZToFR+JLTYrixT1sxTJcG+cwM4bQQHnr5X/3Tqs8ZFj7zI8V+qwa
IjHzfBaPNdOfPSoiwNc+8jZVneuhXzjk1k6wKFoyK4hBt2V1uI6W97hnnDNakBti9O9qW0oRp+qB
YfHT16htf3W+cwoYZjvFveGkzdFRJgMnvR9eSIxQVCP1FJ8HeM8xbNQyzmtbdi5q7lt2f97PPx37
RQPrhnZuL9rVOxuZhDqaK84NGjE3qj35ZaeTN7lkNELI9I5QEv/7VSAufk6FroYamX934NVe94V+
x1PSb4jENm1rexFTwhK10iKMBcX0FVdHXMWFS2b/Yrv3hA+mEnDsl6MvDt0vmcJFPlEOeg6OBqts
Cb16rMQVM3bh1srgXfntTn9v4X+WvCHy2endb/tUU450Ws9OBZjUCj8QJlAY6XWe3B/svhyewuqj
zuwfaDYC0qm/TZzIzv6F9IVs+ONKY9YwoqZyDdnNqRK1nnwNs3U2Dinyqis5MF8QJiqrAwUbv19f
vKLY8L4vK/+dppT3A/OzFUXkZje1ctpDga8MELvpzjVPbITkL5Vo9Ds8l7/Ey7hIsqhfii12/o4V
wD8inJP4m5ElqxgN01QZqO/9jhUWezYGJleGVrpfV5neSzTt+SDCm6KzI7eLYKprDzmCenoyX0yj
VhzvPtF5ke2nIhBF67xQz7Wj32WUq80YqibqGZ3tb5y/Vdd7iwBQKNk3/rHpaHXkspfjQUlLyIGf
1Ttz9TjyGI7nDgMKadWXWniQAomyJfkY0F7aCia58FVDm+OWEOzlto2Us8TRE+sBMXvzrPGa0Ar5
leyF9JQ69aToapTc9UmfEJG1dlRM1+jJ/WvRqj+RRVMHrCP0knw4IyQ6AanmIVygrUAISgUskho1
gUhN1oAky6dfSpoFQrTpAsWiIEft4IRRQAMX3wkvcNwN63X5h0YtfbNz4UvgmRhlrMYeeOHI/XM/
0usMljd0rLqEcX7oy64VGY8R4a84K0I+XjseJqUr4iSoesJ1gTVCob7PapVQjFow6guhbYjSgskJ
Cs9XZaTa0lFSdsUcKXZQdg8xP4yOmGpmjG/dCVJX9/U65RhS/UYTLEsZH9AWo8NXWncwnb5feVuf
cRxD4yN2tlp6Yrbv5H+ad4EfLIRoO4SG56Y68LUzduwRHMafVlcYggW2xJKZBUwSSTTuGQ9cAdyq
cpPWdSIbTwnuSrdEhOro7NAocCp1zt9fNVv5bU/XEjbw+ZFfVebrvZGMmrygW/ZdpJ1Qkl3uoxT/
5+LZrK2NYcBTUMOzX4S3jhTIJKNDyDT1/cCUDDlry2n6OYcl1AAkQB8301YFQk3tz+zoYx4Z+gZ/
kbeI2p2+Z3pf3XEkGlMPZGaz2/gCmuJAvcUx5C5p5+BqPVf1bSvt9/Nayv82i5n2MfCdZQVWc54V
hXOWfGoY57U9UDBfNbX3qWjZT8JunX2oKcpeUVyzhEM5lDZUEfXDfYbWRr1W69ijc+6qUahZAIPL
okM0kqz7aUv3RpZObEhAPpG4imqhTg5hOcp5W8T6anZzrhEDyqiZmOxG9Th/JRS3Tn3c+lCX5SYv
3jGHlLRbeSuVqaz3ZrOEM7R2BNP07i74xyjRyQWgO+0a+kd9UzKkJufXFKh/iQx4eR8Ur/VC18h8
Az8gShZlSqcx+jlwYi1pT9GHt7OMtNWfxgF5Y46x9AtlW0rXtDJXNpZ+jFBPDG5A7eTTrxdog7Hd
0TXA9zZQFdRkX2qOfuvWYqsj45U5LSnCFxRWqyVxlqfz31PzG5ZQwJe0R1C2zXymQQaHsYjeVW4j
tkgaEwFeHpA5dTwWlmsFnQetNth5FDb6bL+N4SmEyUVrKXrLHTHy8Zh2kqmUAGq4oTFVpggiEIhB
h6Byw3+lOkf8pgrVnbV/ZCuO/BGWM1ERX0v74wCSnD49+zdhQaPAXxAcG9+iq2zsFLgSsFgZjeNS
fuBtiYdTCztfRuNgg0Gh24lXoktJURdkhfILm4gdPiwzC2t65RxR/tgvbLvXMrB9SpRCZP362yt6
u+CAgnJI7nYpxgNQCre/3AZVNCUtLr74UtOGSWBfF2XhRZVKYvkMTEZbDfkUfsdR7TmTDbsFTmli
Pf+8SUMMkqpCCp5KtgNc8MNknf5N+1KrO1RIWomgGZiWIwqj8iJQu170XnijFnmhb3o2JG+RN2wQ
OKNLO2EW/DuHkTMaBijWs1fBvy/TFWBU0VLahNhcf0Yf2BFdQn0tunlG1qoGiocHiT5fu8ADm9+N
00Yu5+SKxLzbUMyuPBpbEiOk94Qmu99A5t9YBu9vmZwmpJ/uDKXpNWnU1lUrtsWcJjOvW408VagO
G7sOEQJi9xtw3x9uyoqmsF4srvx9B50+68Ubng7lQ+xltuyUXOT0m36KpnZsq8Yg/uZvbHnajlqB
waF469yLIxkXVVBVTlATa03av9SEecue56vfUewZwpb69lqnq5ner8mQavLJYaM3vEzSMu5l3jHB
W4s0o5lxD40zJUdIkVsD/lwEP9iNigeJ9oj2wUfyeSl+REyOqqsEi1I9mFpMtYJCYdjU2c2IjYbC
4dIqS3meCjZjxcbJrUYQsFlzoySt9sTkKL5Hev5/kfihZtvuBD4glUxoXJeaFB1OL7+GlJKrDsI0
lfGvaPxaBh5qP6elEyUKS+hPtn251gB7K03T8+iV5ozBTF9MuqAdRuxVvW8PzMhxqGmnEqhMn8a9
37unlgAB7FvnswbnOiUbITqG/kB1cLSxAq9Zi6cv+itqN4VYpVkwvON2zcAHxQjQf5FhFJN+IeNB
kN91t+DB4IDG1d9nxjnZsXfUbC0ku37S0OMWlkY3B4Oo/San2+ongIWuGa5MTDGzCoAZtGRSyVd2
1AfYAvaDA8cbfsNyoaGAoWnZ2I6XWBzhRQ1OEJUkrXa8NApfeHbPY9reb/Bu9T/CzVYUFHXsa0gK
kSY0htmlRBHv60KyYv5ZC/2/R5hJhYJrRmL6pgxxZuXwAxndlm9+gkD+/ZnyZSt5KPo/bvSMYt8t
nw/7GO3ZimJZkdyl01wU8Ek5Ma8o3c0jsZ1QJ1H6BIuFyave1xneCELTIZdN0n+5zWKd1SkbwXzA
MACwUm84o7Agk1UIk+SUkw2gQrIb5iPPtU0Am6Mwea/AjFrs7NL2WNKm5T/7I+tc/2+ErtagWWAK
2WfP98TGVEHfg7qhNLI36p/la2ee+NDAWitdhKzG/BjfW7M8GtnFEEAG7q30MPqpcrLdGEKNwNoi
bCSqoAo3TgaXEJtGIY0zgwlDS5v56a5L0764s1p+9NbRyr2gTg8XoD9ECvq0cOJF1IbDcpMNHx7v
OlcqNArlq6XqakjUwPj27apkw/dJgaVjQHwj+rLCNcOz/rd16hF5OODZNQ1f2Awvj8WH37Pa4vGE
tOAdlqaFOw5vTCgvIdJ74qT19YB5UpqtX9EeX75ljL+AgmfjLPCZKStF7pd44Pm1Kot+9zVtyzSi
WQzJlDF7u2HW2xoWw6bbCH1RTgbaLjS05swyjONkjcNA/L1J1EBQKLSrb+EMw9C9OMQOmcUw9RMh
+yPYXu9UNi667IxebJOF+hyvbilhuFp3kJx5QzOoR4AYFYADng155V+s+Q3q8bZBqAqaIlUbXBTP
U6FEIDQWB+topE1scFh3HlDdj2FOgOOaYIcW1/MSxVRgV0hfICY8n15NVTVmVbcR+5QhDFEdXATw
M8gKbdWcOhFxhpRQdZpfghI1AEgSKLmtscM4z4dBfKeHAdl8EvwXDOPqF4kwKDssmEoSxWHSN39E
g3lgMhUq4CFkVNyhgxxlH4rNraI12kpYCfCmV2TDnT0aptlus/qrd93CYnseHAh4E+zz4yYLeiK3
v/55gGz9L1vFWkFyyw/RnKpf8OEpAVx2PQxuhPerod1CG8YyrbORayGH1GP5Zm13zi2BDiTdnJUx
Pvs9H0LYmmHbjTlVl3M4SHu9tmJoOQWz2CMrXxVDDEe2g4ZLQ3aRM9MzCSTPhcBCs2YachMvIabf
uk8u7bwbwrS0gfMeTlm1gTHfqbMuu5q8catJEMAb+ltODG1WgZwCWChFB/axU4JxT3IbEhrUGnOn
DXIRPwJ6OWmgSVey8+cMr/cgQE/atkCywS8MeeQk3PMC24f/vKE45dWV0qTQ3Rqr9JkuOtQIKyd2
ZP+YfZ2OSWigTHIr5gik3r5MwQr34IwHWMm6HbY20QLrQbu5mZq0p+zdRzuslBUQX/u3F8J1eJ/N
Ppo+9noGaGPFKQLqcJu7w65GEbl/Zre67wYJpjhzxC2cJuKYz3Hcry7B+xzb37BsD3eneBGWHo7t
zoDYN54V3DbXl1mnnv24KyRWIYCulM+lW1H3Uea1k8DkqscRza5LxH3coVpr1+N/L/Ew4GIwp8E/
JSbE86NIilosPAPYIttXZBmU0Lh4IJ7evk3h16tApIrwyG0r4sgTcEu4kiZ6IcqoLsR3LkvU3kQJ
Y2X/cIrSEHl/0ZtFjWoFa7dFTiUNuU0QxKxHYURUkLJGfaF9RTV1cHrpy4kBh84t3yix1csYzrzY
mC9syNFljISipwIGE1Ye2rzyVUil8z77jZB8m5QYmOu17IIGj/vu9Rf1LW57P8dIa9btZ9GD4wGT
gxyzGbrqCNbZ5Ac+kd3OlwqZ4mVcj4VL6KSoukc/w5aHTCZZlC6BvjaTHgEqHJw2yeh2Vx55yikV
r0SAlB4uiUykt9gx7xRrsfJn5KJE14FkEtX6yfGRAqN4voz3ii0qlwsa/FkeQ+Oi5fgFD/pHFZ7O
Dk5nEUZ/HjArHg8eA5QkyspsDPZ6oRHz/qJUJGY6OcEW1TPpMyOkpkJ2yAQ4c1qLm1Yrbtr+S/4v
C+fWEuXShf6swdUT27yR68tyziaJ1+2iT0NIwGiAO/+Dy3CfjOxijNG2vrOU9dLHGJSbJRqV8Y2i
/6EATXHjCi/QLzHVFGZD8k4Bht9HSeT1yHHkJZDqn0kpixELT5Pe5zoi8D7hUhyHlRGih+lrSOLh
DD+gAs6Sf7cYT5a93V1sgeEbsb06mSD8VDgRBQdoJLnbHelF6R2Op5O7giPRUOUYZOpsUpa19X58
NZIBDFcgkejDBQMhRv09LNS8rtkhcHZ8iG86jg92cJlfNYXyJpX8qNxnInnk7Yzo0r9qvIRk06uU
M6kcmgd1lyT99+5XbA/4lv3ykMya2+8Q92NB3s82JUf8RbbSxjNJZaeu0ORvYUPAEy4nXZiKuwb9
E/38Z1OqTML0UIEyIp1Mved0v1DHBNmXceYBtJMu4umyrX+Iw51PbxI+9Os+zvZF1GWve1GgLzXf
7qbVa0NoGlQIwRby4l+WmA7qFhDtHm7d8xtvmuBzmGY55CYtKGBH0J9+tPWNFdn2y9z7bCMTCXFF
u9XWTjbDWMzJr7Fu86O8SxSD5b1gncNPqsHPLaJsFuAbYbiGZk80Z+ZCJC5At3aCbd5jLbv3TVj4
+KkS/n+UGBhqIt5u/bwJ/IyLzhxRcotWBAL4DKzuq+FKYy/+mfWneEmlysxMuWceXt66KCLL8Xeq
mG/iuE7fVOfHoSeCBUFZ6KhQ2oYWn6Yd84onbl1NNsNB9nNcuuAu+0Rag7mmB6djGNg5JYcbLk64
gCiVy+a7Wk2GI2eBkht1SkQ5ayKpmJt646k+8WZKt+IZa35WcLnZopDYwBMH7+3M6QKOOyJxMpb9
+MpTEOKVEgpWQIWyUus0wxhb1KgOo334yilv5J117JkTTSClNTbY30P/wmpR3zA84/4/sZB0vSoV
0b5kTOms/aCM/Injy7COd08u8Yum3EVVq3cQdi5dT41ebnzdK1wqW91yGchswW9laecz2DwjMBsr
ZRussugLU7ggXv3MBpwZ9zfeHmcLsFSsQv/AGx36KMzyiBrko6JUorZL/8i0NAVkvH6E8UaEnUOk
S2syv/lYlIcHl6+G3LjGHxo/BQCPfZtzN020RezXYWjTcCzuLdAb9zEHk4w6DcZAYN4Kyr1D8cXT
g5UcRnpERZcdRWI1aLFNllRjoByneOSfkctTgpQ6ACN8JA1+eZJCiuqGOu6Ra8vb5uuJkrdiei1j
XzUuFvk/y9/7t/hJyuJSnkR948ByuJG4IBQeApwTtb5XnzN0qiXfdQY6Fj5ZvhBl5VJl1hOT8DA9
QYcYrvryTli0y4JsOm5m4xlz9bSGyH0r4wc7A/SQ41XCXLLlLmxO1kCsA4jf8pylxsb3SFiQ/3HW
aESFKAGdvlV5QFULtIPCxyXps2PNPZsYANIpJIPbISH+ZQRT9zB/wk0Kxg9zsj9qcqumx1Xqcf+z
sg0KyQs4ZIs8WHsOZ9QAWP1ta2BndaGJwSvXASJUAS5DbKtwF9P6tnRDjJuy/rvWflDcZ6mTyRQC
EFdSngpnONb9P7wGfYVk3dT1uXLrClu+wwCjSljuUrDfmnRXL5ktv/Dk7BOq8+AirTiYTlIL1i7b
dpCAwMd3sHF0VuZHNbwGDXyjHW9607yn35MXGi5dtfIleYBsa6p6YYVmsG6mSu6sUAuzw+1Tlyaa
Tey2Rk7HHmLuwowaqhN7UuLLoMnZiwJlahGdNL5Aft65aT+q161mJzVuM+CzUz70ClVl06WTZ0uW
ogSH64fNfec0QO8FTU7tCcy3KaUh1Q6J76XFZEooimiTTR0n9dpoNKggbWMXBiIO2SU/KNGJJAjt
Sd9tDN/YZu2bKboba44L4H1bNM7Ds/qmU336j0XAiEnxxcByQIn3Y9DYOxWh7QBawnatwBVaYcta
QehVPyCn91wE8JDZ94OHJX4TqjykbpmJBf0wSnCW+Z3YmO//k0xkOTCoMD2D7/P/sTyxGx3VoTnx
kLjzau0TGL3TlLXYCdB4OdPzBhrVNve7ilJBRPtH7oKKBMZKCdzmaLX8hCuDqg8QL29f0fK5pkmk
Yb21jNieAWHq5M80AbbD2YMpXGMjPaJXY1lIzL+5hyTqpr6BfphhikRa9VnSb2KA5G0EbnYduIHW
aggjDECSD8uNEdyjj6f8s7+jFOp+YOVqoyuIQ3k0UpAsut0iQlF/tueYj1VJRZ6rLyx/6vPPbiXr
5sDlfG3x3hoXg9SUqcSkzxOSRqNHmTsv+SU3FDiO6dboELejl2ndAUdN8N6/Z7goiQNa42nLDMTW
vkmqgYLbuoiMsTywye2tbWygCqaki1PgMphuTzL0rtQQliYYDlzyRFfbua72PTjruRbnoJq74B7u
kOiz6nJDA+acnWOKKYyHcpncbU+GQFhJVAPb6AbB9+Un6wb8EPdybMJ4Bc6UpgtUjVKgWh6C8K/f
mp//NPT8WB3TkU+83VHgkZ0bnSNrflpK/ziLNTL5Nx1NGPRwSiJpezuf2MIMfDS5wcJkB91gqA/2
zuV4UhX0/bbupEJglev0lnXPEeMmt0k/gG0mhjJnRXZe34uGRq1ys8rKLiRkYXh7G3EFD8ggzSYL
3afwFw5qVOO/s8QUpY/4hs7xNyhuPYk/fuO8LnoIOF4oaKwm7I7dIBTdJUrA6eiAbLxoKBKxbERw
tskDYjtmA/lciBp7njqWheXOXj7A2jw/bh2BiOvCCnGxVjbL3xCBHWkJf2myoJFcxu/5CGtOg52a
fBxTVkMlvRB6/CIkB05yrGxnw7Lz8CcaxkUrsFuNOM1t/2jAx6+elH2kNuW5KgSZHNpwta3uoIKE
Anjl+OAxUeXDNG5rxBZzBb8yYLdaQ63XpaSnvAatUdha8zpafnCLmvTZdEVIEsCKggIoULy9nHkW
H7pyiliIiaJ0mpJuiTvV5exzk76lBNivXfim33A0Qw7tEglzVNox6HGn5JX4pc6aDevlSCaPnrUi
cMFGEQd5d2Uah4CZCdIxw5ZWJWcEf7/okm8vFyCmUIertmW6XqQJ4o0FRg3jJmDGxcdUwfLobiT1
cvWNl7tI8N7xotI/jomnMx7zYinTfai9VB9wVvfKgrsvvu9z8qSqcra3716WCo8JkO0XJHCTxCjJ
6TgJyzBu2uPpyaEDG++enrwCzZjAtu/M45S0O5CwwlKgnGbDdrduuMiDWQRVG+8dQ6bhtgnVAWoT
QCmzQcpSjQVRn8Fc0FEdMGxLJM4OAQvRByZ1Dn0tKsZAXjIQnNLOluq8g1fATEd25VCbNI0PijsD
QXdFTgMa/88LQ/m4F1+G5PQiYNlH2P9JECNUtFN6Qa4iWsHZfVwZeD5dKV4JOJw/h0HJJVnyi/GJ
JigMpgtRHr+eGv/3ebjO/MY7s7agrvZoKBSnHmsBcfyKA6HDaMd1uLFelryj0WTtjgmYM3vhd0va
NcMwnc7RXhkDXZ6h2Rqsd8etl70lVBucV2VKN3cd3508H2b8i/gFqJAEGy7P2fYOmR/pp37hQ4Zh
5tXvwICYDOKIEjeDEHKmolScLZY1vNp3U2zDRZcaY/jajfTl5DHoBFlTgFIMZZhG+76HjcduCSnD
k+71Or6vlwLQgNDRCCc2d+3DZ8doTlNPG6OwX+tYQJQpzpFsPo6j680Gt+EninodSXjxOmTd91XO
HicCs81ox/V0gKreBceC76kazvg5khb9BGWT2Es17i+UovGHMB9iJT4mX+63C4gWwI6yPK8mPkfC
ZzJRExmr1X75CwPccqANBqDiUHV48CSBjbTN3xTYwSTGOb2bkR0WaRY8rkgt9PtsJVEvn4empKZI
X74h5Iyr0c2aiQERiDkdekt6L+r8XOifQfHGHI8qu4F3B7b7c9hNOsbVygYZDloiHGkjbPZwuRXc
l7cvnMblfNFdhv45KbhBEj1IxXcoPQQRgczsWSU0xXlhCLvWUgI4ZTVhBo0hs0hmAeVmA6jsHLnI
89zvtl+Km4m7wxzXSp1gi6HSfvuDr+on0V3PfFi1n4dXita+4D/QDQAXU5EhEOq6/XKX7KQe3sSJ
QmQjNwtbcy7dTyE25pvEv91B2ZaQzSEnoGzSTZSiXLMKhmnrIFHKpfpId2TkVXvcc76Zh0d6c3GG
1VQNSMa3jwFcjP+6580QAcmV0Y3cWe7UV1+aMjO3jNZKssLm25DnAyKLk8tuk5i3nwJKyD7h/zs5
/++wlrGyfIlRewQ2AXNQwDAf8QnmA9oIPPBOGdSeMb0Im+Z5a5nwU2RaaNfBpRZuFl2k0xT56SKr
KRuj8BqedG0wO8bd7l2J0dfDXsGrH0QMsBW0TNECZPVyjWXIhwLc43ftqColdBDhQtrIjRGgg1Eq
5hXblcuI+g1JBR+LRU2E9vOBZBDn0s09460mUZqcYMKy60I3FpEzzHXPEG6gZSl1TjYF3looFbzg
sVXO0Jt0k+9HQPcqiBoBLrW6xnHRp7rBr74UNrR1edGgW9A3srC7ltHydP3Cld8GgawqXf85LVbz
MCOxi+/JoxtFHUdRM7SC1eYr57jMhCYjmwxsOlf3/2VF7nGtZYqR5LdqPiggHxo0j0U8OKeNOGqG
TA93tDsouf5D2/Qjw9NXjgZ0P6Hj4A72p78uZ+BZ3zu2S1kcVN/LczU3tZqhx5CPMyEnoo8J//io
Q7fEVpr8SE6YU1VPoG/F6LJSYAbGMJUTBXNN+r53XsGgJ6AP1/twYUWzuyxRBvBVgoiHYIh3J4Hk
qY0dgm/KY47dE7RV71jcxdzAo2iSxpUgpN6/QWelF2YVP2TI1YUNGd99jeCNObyj6rWvqtGafzzY
nb3/NCRuTBmve+MqITp3BbMTdQJYECPi8WLv7iAj6DmusmgoxoRhW3+5W5MK6ujpxGHFDFFTb/dv
IeokxK1VY0TD6aaWfrlXBA4H/eXndxHeADzAneLS/Xu3Kx0hWfKP09mOHeQb5dnSUs0lAGKnzr6Y
w6wotigaMjhj+J1INctADgfGuaP9wI9Z26NjtbaPCyZZ9inQUovhacw+qny5q72Un4wVHlvjRWsU
pdD6Z/37vtS24YZOLYt8+dYWvAWewAzU1jl+u/hXCsDgdYyWRaKT/ccPCdFrG9dGwDFuAr8zsVgS
16U4fG7gDh7px+ETHaIYwYLFQRauQWpNLHqEKcVYGKrCI0i34sz2nPUCVUGkZu0B8ocZ13ur6/H2
HiHA+vCUmKop+PEjt3ub0Ply0ymUPXPOTOOAI7RocCOwWsBy/Ul3WrFoTBMprqCqqsc7oScY/6DW
mJpFLSbeaiXuEDUZBGa1N2dubD/mhkAtd2Wn3UrVIgHR7h4vOOQf47hHvisx9I9IECA4b0pj62sq
mJQn51p3o2TsLtPKaCR9mfYc3cZqC5BGFc3Fd1746/hlaLTEUHcw7IcMc6hQl9hkWKXNOhq2iq4U
yJA7kPNAu8I1rp7nqApMiK4xLIUMn1NXe8Bw4X6JOudVBPgjKhaxcIRbLqCi6hUcyKd5D+jSrwAW
ThvscZEtaFRHh4gmmeXfyDCiOk5aQ47R0A0+CSkoCHUIWtkrQulrTb93jnlidMzVFF8apv4HMoZ6
a6EF8J3ECWCUwFtrh/pLljnq6MjzY0PVibs2vpqMVMdiAGWBz+azxr/etGoRdm2SEgWTA5Tr/2BW
rWVYawfP9dKFZQfX24ygqZVlfqp30mrkRVOm0wy4viDP/7WIa8JPKQSmjFiJCYRU86NDCc3zspmH
PjtrKzlVSEBWzcVfooOpqe+0B1uCZzleoAgjn/mUilO4+T29x9H1t7UYCMJWKaozM1LmcYtirP6+
+3cXqQOlkPoMojbXxKz1+JKZsyYKg1w+UO+GVrnGmSDf8uxmb/Kxb1f+4WwnLl70gwPd4UQuYaPx
K1m97BxKq6RGxtQgq15o/XlwAZD6gtSBGAFcGPi8pEpqjttKqC8+n5zSm8dUuhrps/kYM5VjUIS3
cXrzcyawYc6iBLxDLY/VtH9cT48MZCeN9v1HJXBXSrJv304O6kbmDxGS0HMcdKWhITvj7z1JGjrH
KM58K6/yMSIr5k/MOqi2QS6MnDNPt9f2bnjw2ZEbfSF8jnrocCsHZTMeduCQmcXVkGjXJX1nPqkq
Yc69I6Tlhi3ZDbXJMOUZJLH55HVbf+O8Cj6bhx5GB56rQV6l7ioAKoFevtIGlc/5GGKod9NZKmoz
c0nUajJoDIYh0jwQXFHK1kyjq/v9vV0ZIZkB/XEXoS7NAa6U9B776wdkxfnALXsTImOqwZkwqOlA
ZkiUokt2cGtkl6LXlbawL9Y+Un3uLpyz4jOkp1/wGa2RPfBBJzhfIPnk7/GbD+RQQ3g5Ihx3Xz2T
OupqYFWEDb4mI/YVFC8X8b/NH8qySo3e2r8haLwWvShHZfL9MAkPZaY0QpzPg9zpmn4hoP7LUlVr
CzQHwTzxV4a56L00OSTBVY3RaaSIXckHGjSOxjqfV6ozn3hfL54iorkNIZ2HSCf+6dClA9edBSLa
sB0EbcljfOM5NCTYeCbPUgrYWJp5tAMhk7IBY+shl+RgGP/yq5N5ujCuWsC1gFn7bILdRklHtYDU
xgSZJKZgApRJUfn/4EiZOS7xq5w5WEa5BbrHOMU/UrEgKSJnv/VaGcqwiXSYtId+NekQ6lQOisCk
zvVjuieOG6s6KLF7pW0hU/EEMv1wyDHBNB3tN1QbQffZmLc543KsRL+NxwVdofhetHg2n5duP+cM
5WAXqZJSgt0iZIr0/5WJijlImeSZ+wCux8jWEMv99P1eCt5aGvAF9eb1Lg9YOR21ZI4taROA3W5v
x2Zy/NCn5Ib9kmMXiXjOv7AYJn3aTJjmhQC+gE33H6byoE1VzFzRYaM7RTyDKV+lhyvazPq8WdMH
c88KUDH0wrGxWAv3rojFd3cfmBhM/Srvp605U3mNSmUNcDNXjyXgeo6xIhir8vnEUT3v0Mi9gn5y
i1X7oMTqUcRw8LikDOjtbA69Zg7y89hrx+6rf5QPq9qGHkslWnuPyg/YTsqL9WTRok8wVsU4ybUR
E3nOuQaZdcBKNcd4g4UE0oI1EF/dlZ3gcM+jDnAYLcTUr6Kthheg/0lC15vH4ZAqZy7y9il5qBWa
hLpZdWhPHwFnUuxZ7tWTDZrXXqF8oQUHn7ZdjvIATErCNt8WDvfelwzwxM0Kb1o2rpPVzPvvgPT9
PcHUD6oxsHweJRxY2DMCONMQu0jBW5REnJso/0HOB9gtmsJMz0/KC7SubK+YKEnPpuh6a2/zNFO2
AFmGsvBCMPSrNico2RQeYQT4Hq4kgH+mNNI+AD2vc+MNu/fiMBZhUp8oAel3nSfk0Vdw8SD48yaH
yIKFrYJIVqoOJNalkmrW1U4xn0DEu4jzUxoLMwsRdWtgZZEZenmn+72/tLGMW+1kjRgzGITnD+9l
9JLYfHAnnGNFB3MDXxR++fuxvu9Ihf7TdnMR70RJC4sqOV6J7fNf+MvCo5XpabkQb+phep+Lb73l
Mp+gM1AJi7Iqc1C254K4BOOyqc92Jnk1IrJvibNvYApfKrTBtyYsoXax81gMsxWyL6L8E4ZRRBXg
ePt8u/IghgMaJzzOQV24cBv2doU3uAusgYygrDz4uvSht5lLxuvkP/tu+lZomi11CUgimA0Bk9Mw
/CvPqB0B2lEmql3Nd47H2ORJSkcj+1wVoESl8PNa9FdXhTVEnxU5hkZrqXnGgIO06pCLkdm6pPkX
w7csRpkFYgpsZTQ5Wo11PgeAfb3Vnnf6e+Ws3IGP5tzUNgaOwKRXROug7bBQCk1z8HMY5PObnxZw
7X/i8Pxq9uDQ28jQvqRgcPDB+2NV46LJvvD98yePC+GZTcKtS9jIjTrjWqmAUApFQEU+VGoElSjZ
3Qy06fTCqtwzAJwYOB8ru+itzQwaK0x9cKGI1wPRlRI3ePHNlACGNZQqKXvNNZPRUTAO5G4dUfNs
GcbDOCQLzirn5arl7FC0uBkMQUdA/LSSlNuFNlIxzUO/XHmzx6w5Plu5FTjPVLwS5kqCZhEPcf8/
+Wsw+e+WisnklgaqgVt7mYESda6oFqKxVd+/oaLlBErEvhQBMrXcud1pfpJRcmsFEb9j2Tv0BCM6
OPD2OiA0k4KGp6P9IuZMJ16hyVW2bD8sfuHkmzaVvxpQHAzIv2Zm+japR8nyP2DhU43eFhcNxGYd
RgH+7MHhfdlAgczk3AwFi/evYcLa6ACnSXQVqQkUwNtiSm/BdH3+ryHlpkNypX7Oh1wRqcBc9CL3
9o+m81CPDmjFYcmQZHED8ijcrITBA/ztOEhS8kZhMISqkg9FiKwLCkekGHkW8UXAozLRwv6/blYD
T1Dd0gj/80706DUHzz2K1UlvUwx/VYyN6Em5lHXLi5ALJwnoxznB4kTuy+g+544IVcrT7u4w55KB
gWEKnGoLOhklbjJVgWmfDlD250qU+eqnRYpMXHgWudUIF8ybqVxyP+r5Ja2w626U5Z9D8CC9SjGG
WokUEQuGrUVmbM0g4/T2DpF/sdwva4Nt8mkKqrBH/c5tnt5t1IMikTtv8MKvlfst3PmiyKnRWgt0
jEzZwzB5V3V0VVfcFPV1oBeQIVr5/YHH4A85ocEet5xTfTzXI+XM4dxbAjikoQ9E1tKztH+jF8Li
BE2GdLH21DrMCON7sq8q8SHPt9XslhfSZWY0qKtvtfxmIPShhf0IH8DVYBmpl7mIqNdsL8kj18UT
uMqEDHzw9Fnv5PpeXeksuiSc1R8qzTOuntpt1LpEblGrgWbJXv5CkyDgN93rTxnRL7FxEDhIRjdt
mkXBQODwjGDrrXOuEjyTW04s0PVRZKG73FaH0h0iMnI2178T0SMiY0S5Ce5C3pZUtLww741K1Bt6
/4SnNzLB78yRH7VpeRXUApmBbltxGqx9wAlIiatG/EKj95Y2NhKwVDoknKP7bdGRB9bTNcdP3E4Y
wEsji7hqUw/PJB2SZFn8Sjd3gp73lykgEIDrECnq7M6oag2BAXfx91ySNcQbE/Vlr0M37FD3erT1
xxoFKHV7/wniWb7tjkuBmXe75vt09SniYqwULtuF2Zm3TqLAUjrhBonQ85AOgyhJAv+6zGBF8v4t
hKFK7K4V9cDoUZPB3ChBnwruLmxsJYGVAEhUH7FD9ftCnNtd0gBhyMGga51uiKxgLCiDTNiuXqPj
/UQn+0ql3IQV7vIAXlM5C3T6YglaDS7Kldq01T0m73Njz7qak6gqAL7e0Ue/KIuXx7vz/7kEKR9Q
pxgR3q9fbdGgLrxKqNF6TOOiE5nMoKV4u0tdaXZY2vpqYTVsFVXatblZEuAIT7PcMmsgIM9xOorY
5LXuYu3hJ0da9zifdJwLkY+gMtgEdWf/v1VEio4wAPxjC5u+0Wd3ISveGMHc41LAtOIr8C1/S31I
zmufBLTGJTkHZjDP49bRbzNc/f2bsZMjr6o6Y1Hxexz0Y9/iSL+j5L4q05G1DyNaXV9ie8nfpgTV
3/ScoSfwVpmkktYr2hFeXC19ugB2pAhHTvktl//AWrztlSd9eq3qM/Ao5VFm2T42jzhomlNc1ZRp
UtU1bHS5ze5ZNMVqW5wNkRAUbff7N2uCeykl9Xq4qr+BVD/vcWig8S/KpwWtlpOjkUhHSWfqUwoO
k24v77MMYEbig+ppSb4PNyyLoPFz9NvQmso9WEfXnVkuQfe4NOyLrSVFG5u81tceEUyWMCl/rGeH
Zr2EBMd8/IBF2JkWenrSpz8zXmD4zVOssIL2sD6MxjpaiiJTMk9Of/8LO9uo2WuAOT/qqQSQYl+A
+pgC88JwOslTK444O+7qMx39Uw+mazaZzUPDArHP7yExR+eppF9sJ+/8IDwpruK/2TCffVdbpYSj
9FkkE8mjH5Nxd05fsDBhd7j6q2S3gNrhGRV7Sa2P7elvSq6LelVN9Of7NOIgC57g8MCoBvyx8XHx
CPdpHKC+6+DBrhKqiO0uapdFVQ0elQ+IbuQ7Nkw1990IKdIvNBIfuz75wSYfOEC4FhgZjTK5R7Zn
5uf6CtiCSIFl/6HDV7FU5hQ3wnNtO3dQR1fXc0U2ga9vgRClIdsuvSnZVGXtZMY/cjPCKkUsTLAo
Oz522Y15LVAwR4bRde1iQt1CiQHcVNVOXiRoe/wdZqa+rc0QSnS8Ahemzs1WyTJJ0EqSynUhxL4i
By9PskHy5T7Z0SemEGOaqqPqBubDZCi1NpeEUep5BAdH5fJgdIQd4nxcmIDWzmNvsVXNkQHJ/iB4
gp/3NBb5WW3TU37nRzMKuFpfQqf+kxDMKPHrTfX1DQtLZ37L5nH2qOk/G5JyK/0wpDB1m+WIKall
i5bz64a4jJuTjbZ+vvNkw0JfLwIjXnRPWGJSYpZY+Eb/mCksAVakb2qUGPrgnerUqZJi9WpeZVs1
rsjnWnk5/kiLThA4y5EOVChXPgB/hRBxCcOZAalDyV3xX9bUfLxjOQF/Uvk0H95BgsFDGg6dNUlP
OGB5vuZRsBB2F/oBYwa2xIBYihpEQoUabIoIHFmAp2sA9FqOP+EBw1PAl0hVqzEcKBje3K6RgyaE
A6+VnAMV130+hARD8a2I+9n2AY/SbjorT2U5z5i9FfHxfH7TxodPo7A0ZGlfSgjmxnwH4J4ryQ1n
Y+JfaZQNFbjtZF2s2jfxfSx1mzPSAHNh8NsmVcY9l3hdMAfYgb0IOAirrZjrt6d7hHUI+ayLX5Bk
HEMbCQjET1zwWmTsb4rSkuht42Tb0Y1fzLSDcPRihEIu6DB4regWTixCDFWI7sUKn0GAyU2H4xRO
YbSKSkb+4J73Yd/QdTKLW9qQ/SzbBQt5N7xtFxFTurhMaKFRkNKxOs+Abt/rpYIpjQSFLaJfhjdz
eFNPl9rPfS1EGdHF3y1FXuEfqvH6RofaLewh5po1wL3BLa9TbHrFUPbhyGa5yD2/dI6joOWxza9S
AjSzL0ihLXVNNIMHzDdXO0jyXb+ZXJvJ4r1s1wDDfbviha5vY8GNX7efHzpf0IQMtYACzXkBtrv3
rLpDr01rges9yqO/1sR0sVvPNv5V11UrCH5oHyLiQF9zR62Kf0PEnZIwMEnDKB5uBbhdCDQWsnWd
vlRVqL3n1bF/gSheLM4z0fHObfE4L7YPB0Wo+AjCd+cfTVA8RdE22+kjqIxuJW/fy0xRTocTO0At
j4m5naqAKHnVYQilHW3cL+HvOq/SLCHZXZSS0T8ptt/J5XjLU+6Rih4iB3czPbyVfC06TRx04dzK
7gHCpD3w02HHOj+3TbdaElPyTwYF7w7AJvZYsEt1ykxyEn56fx1/u+eM17e4enVSVlJbNmwru78u
M4hGDYs2zfIbH3s4XBgBL0euuuy6RnTE4unf2vQKNCXk6YWfVufOpT0jwLY1jaoHdUzW76cLVTls
ZELSvC848Z78HvoP52Hsry4Z49DMC8uTbjpoxBV+z2gZVegn/ip9P9/lr+PFgAWfNVWYSpD14+DZ
CRqvtqY8KY2pxJVqajMs88/gYjp+4v4ugx7jWsnvUnAIwQZQfGvEBX2QBLaqSGlGujsngtqByhIV
Pce/EYZypmsbScelNrEQbduQs/lX4Ii7TCgWLzrOV6jAQevgQ9kkMhBaUhZv4SWqp86AhSQPbuX6
ncmoLlXI883QdYRoeC58ODOk7/n0UwR6C41OklIChWU9TfwnXbAuvcleXLDswdxdJdcv4+hrRgze
zgjDRFeaqevTQyq8DeQzflmdrHmI3uzx03S6mfQERlZL3jym0cv3m2kocli1HRry8YPmnbPag3EX
Co3cA6wkN/tLehqYBFEu0WVdc1PJ71ARyUyAkm1DLhf18GgBMdnXW4t9OpTgK6LD4qxfOK0efTaC
0RcUkKqJp/VasFOxW1oiMF5Kz7jIO59/nRSkEYAwL8QD6jFW2jgIr6dHKGhZxmSk078WBqgFOh8W
XXXehDDMqpXcpn5ZqQQQoP+JEGIHTpuadO11f/BGor7MWhD8pFE2ARgIkONVxldH+OfFyzj/HbIK
UPNxvUZJ8Flgs4zfFud+Aw1stkSZkV2Cvc3ouW6ANfYREzeQzLu40XQOW4kjQ8sj7SJ/m6QWaJsy
ntfCKUYmmDbR2OFZxSyimaW69V6GF2L+EvAqb0+pcI1wOrGVBhxsxiG5QXh3KCt60+Af4bhRybIH
iKeP2VBppXm6yMl0zQbhDeKt+5RU7pKoRPacPA2hVdrIeLX6dXgu+YjpuFpanRD0KDqcD2Yyzvb+
wC4MPJkKW1UqFdoMGOGYslN3tRDySHuTg3IYX5HGsLex+FhB7rEjPgFn/UbewaGDgmNv04E6R8cy
mFMTgwT4DIA++ahDF5p1CfFJQ0DXhTQy+nQKBaiYD0AlPh1G3nU5Xc/1XpdawRKROVfEKyYxRtIb
+YFqr/n78FKMsparDljGg+i9CqxqVHGqFquahknH9CoPnYgRZLg+EfRORJ1h1OOzOJlLBj0ZWAsW
e+j51qAhOx9/mJFet0wOK+L8AgnbpwWHX4PncPbO8FFOSIlQ8VxSXk1hYacqQ3677f2V9BWFzVB9
tHbB+WuKlRGRq6GFvmWV2FDijlNeTVO2/ymFRh624Xp8WY0/Zbc2Jd9DpcoyZyGDfPe0cbrNj2zA
bfAZ82a9K6keV/4DCdRIWDH6EpDUH9Fq5RYWrTD4BDh4E1lmGxWR6FVsEjdn3hAio/JcVUmBCPlW
mDCDxgi0qd7LhdR7UQk0rASXBYblPCzs4eB68JGKTjtkLaZ5Ay+iAZaoFO8fefgXZvik4kihD4Ii
Tla8CEX1Qz1yoHisDix61FFYpVqC75FWXDscO9Jh7DgYPHPj7MUnCyc0dOdi+KghelH/NKFs3W6s
t2YK/5VsEVDsQTSR4aT+yaz446Y145Q+2T7X0zrbgfEe1tGD+2hFclhzxHOxczANDRpbUdW4jXho
MRBAvLHi1WM44szHm0AIbo5j6suqdpsBpwqALL3T7YnhA9PmqNJ/wCCoSSxTtXncvvZNq32RZCjs
ywaGV68pFCK/k0p+f/tbT4mPYsOxXypUnLZO+UYNxpnYa4s/6llaJqyVhkrOBHwYdgdxJBahaYqn
JeLzrCOT1Xahb2Gp0mHEA1ZftmBkdeLTqu+YMhRPNvwJKgSovB2QE7sPTHBBcnGfV+2wCeMy+x/U
Wiz7QlSzg2scN0yJYO+cVfxR3r/HBK7KkuwGJYejH+xk61lliHBTJd0iJ1cSjl9X1FLwte183YGB
hPRY5R2jTOqEWk7/l+7Pz5RT3T59BbBmahD62YTEX0Xxsb4ejJhvDZ5uMZNr6IbCxD96iLZXzSmW
XT5+H27iCykdaVzenLKErxlIdq7z7ARbIdm70hHM2usfRVXTQIRhhlveAEVxd95I9Xk5IoCHSgeh
3dZYOBZzzB+O729lYcFMwNQEZPyPvRRr6iRp/miBPJvPJrkVLW0Ygp08Q05Zbd2b/wP5ZhiD6QMQ
1Mm4xnFtRscf14ZMaS0oo6rEfI+3VlpbZMBpb/jZjGPM1tmr1iJVHFbJMsVJr9aPU9HGsPpOxXL4
v32ibBUjdw9pnzcyPN5/BqJ87ST3N/7b0OVjn1ppmODuFJz1eVUpPTlmqc9FmaL5rbNfwzSZKdRW
1N3ZT3xwk2BKjpnW1w4Sc4zoHWHse4rmY6cUwMWkJ5Ah2Q+3QjWaYz7WXjSEBDnWjoackWp5g6Tn
VvLXBaF5LFDUr+fGfrJ7L+NaFvyDhWQQpYStzVb6qaro5OeM+o6L6XmBGzcHLsbJcUKaFUi4Q6y7
d4FY47as78/jF535WANa+lt5Xp6n+GoVmM2IV2y4nZvMsLKwQ2/ejUU9PrWy4iHOnJuXGLsihvH6
fNE93EFwGzOP7/25Id4rEhjM23vuwXl6ZoEb9XHhVM46gm+trlsUzHqkhw+ayVZEzeQM7t5CYA8p
ObllqtbffY/wjEPouRbCfvgp4EpPvzMkffpX0IXasjbCjCDY0w3Fdo96t5LvDEjzG2LWJz7GObyn
w7/KlWHBrT/DDJ/2xGEqfM3n5+r59wKhWN31A0yznLToagF725wyXzwM5fJavp5n1+ZNTaDhuNjU
To7/u5ay3wgd7ygoyunR1qOyYm12/Jw5ypYKVF0JxSNjTKjYhmnyZD/Yt15Yci7gW8h+GeQRew8C
EIOGODimUgRObb1l/ru855rVoPIPXJyB82ABOPDxEwPCFrJuhw7Dor1plk8NsDY32Gv7mnZ7W4m8
vZp9kqUAKB3hist7Gx7FQLK+cImVuRUfBTOcXWK9mAVi1yHgMQvhxpe6FGxRNv5Sajp0kmMKIUSS
n8Q5jhOPKuZPcMEwrlaOt0biEAi8l8+6ZRsSW9jeYfPDDF0c6uuNVlAsOfPSg30rx48u0X0THOgm
UVVsHz5w2MNzq5R5sneEJa4FXTYHOOKonYQLYipft1UnBz+ot0oZyhAgJdlmYmot1vM56Iq0wR5W
SDM0LpjjgjzLr9xjUKOT+7w9X/6GRyMmCTAnY3zNM6fX9g6YyIBOU65N11PcnjwwGybXOXsYAzJM
HuwLHf+SLZhI47aRsBN8QV2X4Qt1lHUvjktep3JXSXArnJ6K9mOqdKX3d5tBEjZ+cJhUYTxjC+t6
h9bnMKgKQ8pmCcxiyH7apn0oFUo/pnIa8FKBSHkVfK6X9qSAJhpOFSsAMbeyKdH6htRCp+xMtJSB
bCs3MXDjwgfOKYbvw9lSmddXwf1KzZhITFcSy1/knoNJNCI3sS9LlWpKhr3IkJByC3ziLBHyfDG4
FZOmYLNMjJwvLozQIdgnXeGI19GqeZmdAFvJhMyFR4b107vB/BPnHnc175GprFVaS/eJFPtgCwGa
bZ9yfYthRv0c6c0eOUmk4Ga73I5yZ/x3qC0ecRugm8J1ygmWwzLESaQjdxgKrWZUOlNxCYDL9UB+
uMP0E2wdqjrTbN/VI26kbtbM0XdzcBt/pixcnBqAVJzLmc0aHp4/94NYR5JxZFoEu8+A1GeRUsgI
TeL1ujoMsbGyiDWYubK1UAVrw9r/JL+B9gU0ZSrfuDiCtg0qKnSDaNGb8jQWOtW8sgMmgcQKmW11
ACwtyKssSJj3pBdrsliDIvt/S6H/cBwr612Flnun78iBabZFmhOZlVS2hLF6MGEwMgRlLuICY0Xp
KJrnYWvKKshdDMNzfX0gy54lVK2X5cUo58p/6BsRZfw2EuNuw8SmSHV84I8p1rPAbbwqYXM02ia8
/izTG8HxPRZsjTDzTo0gEOJ1Pt09S2PBqW7F7QHwNnz/Fxzylm8TV8n6MrKHvnpGN/cgA8cICywD
GBp5KTHgX8P76SyuQMq368Sd44Z1Hk9E/MUBevrzU0k8DBAciK9A9AzT6H0Asqv60zcSc4wpF3nh
IVVx2flns6J7tcPjClePpueoTJR8wbJk8/GxfwDgGUIcXsGwK5nPnfQydMX3YfSVA8h/Fvn9aVcb
AlfxXHq/yJOHJhqyjSgWACkIEkMkid20Z9oPR+q74XW04kpB5KJ9ZPcPGhMKv2WO+6TaRCF5owxg
eFwd0+OzV5Vpr7QkEAh1MytRJRXi3Ef0+XR7o/YzoM8WGi4TrZfeSVlBVERcmY4vRAm+0D2Dul2Z
otJRabcKHhFi3+qStOWLUIZgm4ovGlP1TG9t+pP45CEZ9I1HXAta/t8SUIrpmtyHuDqGrmZwNM7Q
rbweQFwusl81xUSfAxCWCl5bsdJ4USBHTsnDrFuISPYOJqCVs1wuaGpJ2yoIOmBnECzLMjVhWh4W
0VfeLeETqPEsgKSw913fcv/BTvFjrhwTJqzippxyCNvZTRpNuJKALE2ntjILj8Ktn8GF7olgrzty
H9D0Ba30DYv0eGLlI04+GGwQhy9ObLv4UZYzhMXvvIKurAV4PmmfLnO/BcvS8SibsldVe07RaK0K
bklz7qSwib5Lb6NhKOTqz6lz7+zN7n6ywTgianUz9Ao0aw6/gfLwdRB1+D/6k3TK+7YH4Byl+88q
dr1w7Rcu2LIhEo6gRg5TKePDJuZcUHL7TaX1U0gIs+bGtVf0FEeCsXJHiMgkGZSi7MJUUhOfsZeK
dlsCUWShM+jPRC/qyxl/HkrOK9Xy3xu9K5HMO5AoxuOlzpjPWuf0pIczxkzv5bNy9Tu3oI0MzeAN
R0WR7YhistMGA7ftQPaj3v0QqFhpZaQpWlzsAjBN5NOj7RVikPTyqjGvc9frtCHVYtwC5umICkKo
QgGAcHI/97KeeIqM5d4Jyd3CpQvUU350M8uRq6afnDDhNVq+UPjUsR135gKTDmrgpFw04usxGmrE
P/ZCk7ZLJg2tUodGHseqTs3/tGNrD6iHcH8Jp82V7pKFrSlaaIVMtmK6DsWl+MJDvKkt7E2Znq8Q
gB1VdyI9R0PLsL0U1IvfdXhtRuDTZmpK+B2P7yT5/G1p65SiUVl5uwFQj+tUSDTsT9MAr09yT0Eb
1K2eCl8CuqBk4iHv0pLbk5TdJscjo/tlejJB/Y81n/5zKKy6eW5Bs/Y0UuScjR5+8KXkKCac59uu
Wxi7hltXFFtU1nIZfkTfFtdQ+IT4Y7b5AEjs8O5u60bEdhp05liz6Pf+kmZ7sBbBgu2YxrjV9ESy
C6lTeJjPDEM6CMqAuWfYmiz6skIxKDHRHuDRaVeHbwQVf/54Vf8iyBkTO8+QqeH58maypihpUuzn
q7P3HtfE5GjE+pbZpSvh48KJY7TtGFHyp3VrckY+uE8pJXl36CPl1X4PR8hUoHKiXxxKH87Lb5Ov
GIqIMeRx+9jdP8UMS5qTJ/dmqgkSfujH14rKWGaLQVoEdC5dAm0ReFpGqQ/y/Iw0e0NARJvImtOF
4ZrEy50HRTz4q8aqIARHMN6eQdC/4i2gAe1V09XViO0on7KYNld0pfQu60N8MgoHm0mtA4NYlJAL
VI78LEWHpRVnjKJfz0Je9XaLcKiWwikXZsxli+tR2Lf3yhIQbvhSgTOKypLnau6YaSCYNEWM4rU+
ktQ+IiYbhwfNXqytxbkj6xXdZ0jgn5PFdMruvQ4WuACqqRfnKzTDh837vBfr0UU+naKLg4CB6D6w
kbfO4ddMbMPAxHY5yuRfqa+zf/yFtWm2SetbvMq5wpfhPG/noliY0ZzYvbpRXgBAa0Ti9qmppLEV
RZ1LMTX3r+LGhoAQOxsJdLvL/WbH8i9k3hHuaxNHlr4kffXcBdNkabCJLDv6aF0317cJXqJQKiGI
Gp2ubVJav+rY08XbvRZTvcJLJ7h/OlIfT4jtmZ4a7834lYNzrPak1MON6qFmJqD1gQbyu1YEOUG5
jTdU19HQTwtLguv9WRYcG3IZmAvP0XNqOPXla02CNCscgeYMlV/vV6Akb5+jiW2MkrJt/BuoXVyR
54ng0OnuHfOfYZZuWuIioVvqeLmwi86+mGtYhnYqpovxbPa5gUWwHdP89Uri6o/8Fyvzh04s1jCh
MxKT8xYESWX65rfThuvqcpF4P2K/Yv6eJiheTEQXllSyqgLLZtIlXK0PT4VUsH9C3fF1K9JgvAWy
xMYpjB/RAz3NItRd4xOt8otfhnD3ubZzyOuhcLbw1QphMMSGlJIfavnmuKWzANOLH9ost7L9UWLc
SAX5iBhL/YZ9FVMxhfdFIofSa6PZkm/U/F/GIAtLDvM/wgcrTQ2BOs1JvKNFzAt56IgNJO/Ycj7W
5T4dAf0wmNF4Nfi15qSEUTudLQDdE6a1QDGHhjbgkIJClcamG2UsfPVvq4LZnKOOsiU43KQyWn++
7kMHijLiGhWyAyyaASh2ZNa++k2lxS8amVx/K9rTLkFwniESGTennxwiwpOYASqTkST7Yefnbz8q
Cw2DW2APWpVvOdtkqwe260IWAZ7Xt3xHQuiblxbfVo15HQgVDzDxA1/NCBOe336gH21B9lIIGS3J
wAQc0cxBDo6UZNSlIwsWNL1K34Vy6dJxo1ec77vPm/CJywNOY9nIe5dvzlXOQgptfatNFukuERo+
pB8Wqpo8KjxdnzT0D/p6RKvxC/cGP+Tx6dSxxdLIS5I+5epFLtNnHY9Zh57AvnGi+1u93gZF3mH3
uaknwW8JqcdEQAOf5yqPBzLw9nKI0oBfhplHakJ8jXfBU991b8CSw7lRLicRYWf5M5Tkfk9KqYDE
KUprWRqDPD5O5cXb1uCfj6P9AcO/qhLMQguNIBLYfFU6x4caSeBHQyy7BDN1ZCrO6wrz/XL5PBo7
LIMPAoFUAZqMuPgJWzTW5kxtgs76SfIpMwfmdHNY0MuhkEBxNimoeeomZSTPIVJwWuN5aKqZPQ4+
IjDWhIfFWM4VI6LAhhbR1nJiNeNJfFyqh2iWy1tleWy+xe7P5ilvc2YdFlVQChyG7DrT/jUjBD8y
ZBziNB4p4tYOOk5PFmlPL20F6h77m1tQqIDl6OYfYGXmy19zVWQ4XXqiPYRuJ56M6FKBkKQ2hnjB
q/jk8/B52/z+2KrtdmQjBoo2+HtizZm2ufEvQGd4OlTr1+yWckx0CRlv6vkv5GapIBzNgx0ypw5Z
oP0Xfa1eHqM40qA//QaEE1d9h7VCJ4/1VsgGeQnjzsadlJS67EgYVEuTC6YFz4vX7Snvhks0vpPQ
cF1p9vizLUX6tDVaAQGK3xFH7HaDuaowFpX0ip/71tG2Ui5imMbrJob/EuZhvSBbUsHe5R/lxWKD
UPe9yeXrupVibi+WJyJvusG7UAu5dyxsZnfa0ODm75jxn8fGZGwoebxjAroWRSqyJ6F/nEWzTDe2
j4dXOIs+EW3FAXupf3OyJetz/bqaesok1BVrZsRvmtO9/8IJn2mc18sIm3P/XMzjGo7XA8CojavG
vDLIrjkphVemSRMyHqIee09ACaV4yycjNLxb0KNYkI1RdmetRQ7IDGQHNsu/s11uvW1ZiHZIrBtd
rK3Y1cwWg1pw8Bo3B+yh9gYVnrYk0Sp6QBMW8a/hbLnsl4sJY/ekTMmpH20aZYZP4e2UBcrQDVJ3
rlwanPigkjTG/YoTuXYkYiCmA9D/6R7nGzgVe0jSIQAWtvtgOx5UTnC8pdPHbzFahNeUzxNB2TWV
TpmbG/hxtcIrZhQ1bFi9pllKvix5qjdF4OxfuWAhO268qipdgNfDaTyXtx7npmo5Uf1nCs6hSvPO
QzcWBjGcj0nkMLg8VrvTBuk3H7grCVbkmfEZwG1WgJzsSTRq395Z6JPib4kF3n8VH5Q5ysclBFuZ
TBWPgNRQ4QdXCBrIBf69jGhd3SsQDrgglldahPoDBMsQtpf7m8MHOOHc8pPzVyLYdv47UZXk7SJj
inmDigyLWQy1Qm1qbapAq5IPMhkwPREBGCa+8VKZvDT7cR42rRz5RiOfifB4Nqc8Y0O2ZB9EA3BA
VSMee4HD0QhLSSb/ONQCWsTu2AuxCw/nEsft5Ha+3jPQ4Dmkr9MHga7qZ3R8nAJdHvLI4FO5gWgR
2++GQvxawjJK0axO3MS0DUCaWizjEBV8F08AR3b3Icslp/weZLc92mb3jbMdmVpVJi6w/Hv0YwQ0
F58X3V9Une670g79zV0JoJjRNeYyZcjJq11mvUoVxcSw8xLQwZ0IBtUAeZs0JcedMAcXHOJNzJfm
Par3pPIbybLop9JRDyGUCj1IUvdLc03fQOFpLNeoOcLYEVdbHxHc3Sf6+riIR20kLJTdmuJedEmh
+TtCeNNYM/Cpoa5k9apD0LbmS12kw09ayyfpEFyEMldZ7ODYQToVJxv4Oq+8Ffenc1txBEYBE2If
CcbDcRsp/elGaWcq8MzSWY115JjVgzw3zpQuTK8FwaTbzcGLjfclb5aQ1WQNejuYmiTBpqISPVwH
XlmBoaw2o64z1ubjLKP+Tf9dwJPhUSBr7VE5mEoaL9M9kkXNjXB2BVdOZAazGJ7yuX6MRicyQwF8
sSnJlcMGDYNyblHlk0P4zYKQy3guJ9ufX+tpkznB9g+SdmhXVLIc9hjj0SFyfurAELevLXEOlpRJ
+Ve2QLkDvEA0wSZ5wIU45ZJ5mxoKGmrW/9De3ylie21HJANxcshPeE8yw7RD/8io8GAPyvQnW3QR
n9SekdkTA6lzAufTkUQcdnZdSqUGQkvIqGkw8QmWgM+B2RkhdRE8iKb4YR+rjbUWUSzrsIBDt34E
AGDRDQxY8cnBVXVdEZwuxGnQedWWN0DOPP8wP9GR4Do9+sdn74HUNrBQeNrLydt3hZ4ua2gV1HVS
y6aXbUXuaWz5en9a9qzYVlJ5Paw6nSqjVc4P9DJ3t7iE4VAQkS7YhRuM8RP31VfyRfJxa7KbK9Mb
Hq2zkLfCPvNYExvnLLn3Cm/yI3Az43+5m8nH6BFDQu0rCO9NqqTXS64jlyLqTjMlK19jDnQt91wY
QX93NWBMw/YfDS6DeM/IksaInCMezj9+iLi/gjZkdXSYbdzn5hQ7sCIriO9mWyPlXf4ZwZ3U/jYo
dxBBkV/JcIrZ6QxJblAP1b44gSQyKRUPzozFzS9tynJs0PtjAWfDq1rSS6USYEg+OXe+dVih9aCk
pcgmBi32vE/Q1ODDvAl667S1hMl+v/Nl42jZZIMWqNE+8XjEQTX89qvnJschBAIGF63u1HsfqPDV
yUd9kn/F+j0VtnOp1fE6Fn3Ij+fLA7aJhTfGuasAjkaXDVB5D7pdcgu4Iw2SCq8J7gOeMLRA3Pj5
cPNZwry0xi3uhf3ssxNPGmoGNzkBYC9SvVnRzs5pNkfjNrNi/lGRFM8y+RcueqBQenJnUfI/8bU/
1UaEy+O0l0lABRhv9HtepWAoy49EqlSlfOjxS7l/yL1tPrfa1AThVykEIyeet/der1hf0NGS48Ij
yZEEth232BrwUa+2XJnSgQcTzIF5iUQj0l7yUUwagF1KgJnzVVWWissggZuhzxC86kvVuMRnQZ/1
Ej38vSriHAXY7qQGCgfRt9TI0rTGuE99AixhvVDo0nmNiNJ7L4LXiOigWGDWbEdQAHBDGcMcslhI
H2OCiaJc7mV8EBfwy5/ova5Db+5yojNMPRuX6JONicQlIyn91BZ5M+/kz8omnBlKUCDOVp5XUPdQ
HRIQ7p4om4oeMzHh1WYR9/5hl6E7LRN8/hnF8o+jZoGUYmFtQ/hSVolDCEBIP58DdqdiMVZA3S/6
ipOA5MDAG/3CKZ/dmtSdoWodVUOmH3rwEWoG1IWXTbQYn/ylf/hn27iCW40fdk76IrLawZWPyegz
HuIuglX4LFMPJK8nIK9UsmN2i9CszfsXOOhNSwa3iVJvNPpWPQ9cZS1xDUnhhVyutS9t1EmED6sa
VWtYFSDWLCV61aFlNDDxoDtF+PkzKqjqHmBAhOqHtUZPxjFdTRtD/RMNXDBfGUiwekqGk6PN+dP1
iK4Xs/cj1duHEtpbnG+Ery3r/a3h8MyVXrIhmdnX4IMuPQGS1q+T+2LY3JBWGXyEvV9Ov+KW206o
C4Dqbiopb7w784HFqeCrMnTwvSgU75QC2j2SwSCdjxLDI5Mn9rS9ddjgd9YTaTSPByvweSy4lL0d
iUyjRIjvpNyee1jnhlsroJOCiDpmlTNkz0d76kkXqHDQfbOBqqWHJLweQ+FXejocSwCFfthYWJHj
1J9c4Jl0djGOVghiM+co/XVhbu118PoKud1xUMKCfkAnsXoAEsgY1nx5FVywW9gr13xkhLCGj2LX
AQW9V4doFly9RuYM67YsOBMwGZHWEvYfQ6V875oQmgADtvCaCyWgomWT3TebovJTBLkZUxGZgZt+
DnwF7vyjeDH/90Lcyp3Eg8/tl+rm4gr7Gk9i3LKltomwSPtm7bbD3OXXWXPu9gcPWNNdazzGg7Id
1aUjiBE1jLCv6AurH526K40s0MpPwr8wOkwsL9JHNMr2E2eMhltpPnDALHJNO7Sa0L45BUryBeEM
J0W0HYCVsMDUIBGoQsthl6fG0NYpcb0IXRW+Fadh4jeAPNJ34ZbFbOY0eA3f+l1d7G7A3/+hu8iJ
g6JCI+LSKwiO+XJUFxdnhr1PT/D5X9BYz5hYXcA4COp+cRs/a+myxQ5Hk1ASDFD+k2YSZT/DOD9e
9yb29vEDuB2vkY9BqNbOEh4UQmhlcz/PwuJ94Gml2sbHGluTOW31QR0EvI2MilRHmYSBPv9uV9RS
+BUVJWt7/QiJ3R8y/8d7SKH5VPIrbXjUAOl1u5HOmiTaRKvbfKnT8PGizmeadO1OAeUXUyycI+3b
to24rc9H0CekoyCO9PlB1BZ7+b0UA7Pe+9QHL6G+dxkWKtGRUU3MWphFxUlfCLj8nGoZGK34bCQv
doX9wIQ4bo4e/EfjonIiUyNoLKWIM73nVQxp4eSMPiseQPvbO8h7c61EvMchQzz08RVwtJDrnhjv
RBEqwf3sEf8nMXaBQLQX0dOkFLkQSNXQiDyzOU1bfYBUPvOeGiH7cH1j9Wxgj9IaF4/Z25fW/gDm
2/qJB5t8Vc56kPW/WrQgFX/juccBu+6OJQlFnunSGbdqxzUowaGbdfBtiOdk1Wd/V0xCW+2wKnke
/3IBgDMY1vQm1RXfDv3KyJ6AYNiUDz2hCt2FnF6O5ABhaAqynmbqDNcqLWsqCYbLA4hdDAlOHAqs
0h5RG4NuUMPnWv4L5aTvE0xYUBpI8sV0Ju22FyQWdwBsL2l3n2PFL03o2g2wWGqULVXZOLpRxtjv
6/vUO/kdEvmaLkSk/27wRKxjkA8uDIIdf1Acg06+tiIUtdHb2+AU+eKXTYefgZEXjhtyq13JHyp4
pBk5aD4LWoNdCK95gqTat/lOQXKbji6vE5jCeAG7qc506KgEs0Z/OcNDxEHUTseIfcDSp8S4/FAQ
kASfPkEcp8sKxCKoRuv6znZSQiGVAinpBfE3j/I4b8ZXCo/M3S+1B6twlYI5pom63FtT9honv5Mw
fakZuAV68UgUFZq4/0glnZukeNOfxjP4dyIDEbkJHib4yGesODMJDCSvG+HOZk34R5EUXD0Lh4y6
vxZg4ij+XxgjWC1RpxTtGtTlX5wFBPtB/lR+QE0MM41OhKJyhVKgnLDtgcRiYPoBbod/DB6AuhXF
sUiTlO68TZi8gJNr5KLA3ehO8dxjNqsQvLCn5n+MqB/QDML2NZrG0SzBxMQsqxyHide/PAgR6TUt
UUczgzJtsSd371SkJFLg+PRiskdKN0pdTBwMe8TuOqO+DSjZyBNVmE6wFFTRMka/e286/i1jtcot
yut1ZT84G/Qmy48Jw31WmyiA2oYgYRAt1TPsceavcUGfLVgCL08cBRXBPokrlAvJYuLvQdqR8mcB
6hBEiO5qV3OLQnDYZYjd90VCRKd3GoI9GYGCqwEyXjBi/JScq8GlRu7NQTnfExtgmy8nwnYLYHGF
UMRmF759o0yVdDg02kVt/MeygLbtpR4p/rzn9pDJ9mRqtN2GXSJRdSnEpwKxdyZwRUqo6Utt2x34
EhGyEfY4qqfOmO73wpH4m5Yd2gW6MV8hIPq3KcCb0ykfPP6myeYnWsqDo54B/7z9+3rpsPrIcNYN
yXvGR2tfnuT6FS/NpJ3sC0nocO+vApP1l3ILuNtA7NXfXQaxPCTfZbFFmNbxPMHsyf+nQzC30fvx
6LrSg5mDXYbhQ0W/wNdmeVmpUOrX6NUUvFt0MI5gLWuLUlPzek5depy9Mme4yDKJp+tFodGCxTU7
5ugeX8hfORQFwnJwrdzdRjj1mreRlNERJOYTJoG7ZE2crrjnoH513EFkPzJYS2KKify+n0CzdwC9
anNgiREgjWVhrRG/oBg21D8TtyC9m9lwDWNh/1swmE1U/qMrrTRvh0jfb9tTLQyMvVH1G5ewR8Tf
bZd9+BiTcrNmCpnG5SeMT2r83hsvEHstMRoaihhzm0h2pWvhVtm5hqBdPJxA2rJeWghH3vo4K3gy
FH2p0ABsf7sUvCpoB2RlG1WrjHcdjRB0dLryiONKuq604W9OUOuJGpTN9hcV/jG7LdYpH3AMoWq2
u4EJivQcN5PuMeugIH3qHMv3tf8eibyhveAAjLFEPVLs/v5srauwiwNqkncmHAkU3G1KorhfHfJf
e4XPmJNG3m6oeUX7wjC95VYgk1++yEwbKn63ezUgzBR/ORFOCT4SuleAwQIvNi6PKmT6bgxJ8Xjg
sia9avY0akw+pTBNEjuR5M5sh9tr9jW1/dmdsPDKZdsKs/tfc9YW2lRDgd/ZE5FaeMuQ25gEYEUz
7ObGHKKUSZypl8Jd+4dVEG3MHTyI6KAJ3c9TLksD3fQPjdJDaKDbYWVPc3nq+NhZv0v2rjb5iXsj
815iplBrl5cAJPrHasmrOHwC/5wCwOW6jGZ31mTW+6gVsM3z+vZm+Uyq/PymafiP2HHMubtQJsci
8+xevw5RM/DsoeYU1JDFrSjk5ScWg+Lu5JH3CQoUtuaiScyKDdjO5o4U44uxt2dWxC0cilvzFCY/
tiXSsYGICAjQxCdv+kYsn86vWd7WNp8dz082wIqToMvQLtD1HQU6T+QreDUUO9WNzS69/gQzYhP/
Dpy1Y9agTmHueXxQENK4FGcc9Ehe/A0beFp9KTNT0xkFuauLoEcXhjGBJnMVbcaFLb4wewUQdoKy
WkkBU8VK+FJNjQdfCjuxhafpLGTT9dJKYHTERXuqLJitEmWIP/rZ33RMnktpVugJJe7cSaHcHhJ+
nYWslBv7M4bdApwMUeXCOd3Uq4wU1lzhAUz26WQfgmmZGmkuoWDSFgkHxEPXCTk9hYB63pr1Dbzy
POdn8gxBclM2qIYJVGftGZpejNY4HUEsx7566RC+9k1KzQXU94Ogqio0DmCZRFuNc+hBjkq1eWYB
eluWkhDbUZU4zZf9m3I5HVvCEeW4SlOeurECatuIvbMbUCaSihGdfuq3obYtnUBaoFJAJJYWtDYU
p2g8n5U6a3psrePb1+bgSmjDIZvocpA2DLEsSQSp0zmWuhia9OOKVEpBxiwId5PATjPFC/53HeZy
yZisgcGEQyELdO8cEnOPLPhsF8LT+QQ6olb2n/GfMny4Z5Q+e4oL1kUdu39Wdbznz8GsfXxgn6Oo
fkZf77yDEVAFOjm7SBvfhNycz9jEMw11WJMdWLjekNt8AofjdGyqVgJtQU7uLFzxmD09U9kL+2FQ
6s63QVZ657chr3jS117Rn0B0LE62ulqZSju7GIWhHZLlW/ze04BzKPVzh46CCsAid7flKA2sQ79o
d8Dkt0tFgUqJTincF3PzHeMmLFqB9QzZmWERVkaY2X1MOwyy0iZ7G2aCUcquIbR4Mr0XFH3FbgK1
klkzHKa+Uh3+zhsXMDdqjiR3edcjExKaIhyPp70Y6bf48rPzH+7wop7+d/RgwfRyWwxfFOB/l0in
BXYlIKy+DDa48NFucw7rnLiaM42IrTqrOM7fNp4DBENNqGN/xoOrnTPdvwiVFHwG7dw+Z7U+cT4a
7fWDINAffNv/UI1Z6UISEGoika/ZWz46SW8nNNeO+22jo3XtHDepjkrGeQ0u5SKMIF35QYaAWkX8
z3lj+9C8+IyEhU2TRFPAT1GulGn95dPnNCGaVuXybATifs+4gRBXcTCQ0rLVE+j8Ks8/505ca1c6
aC6I+DxLXhm/SR7oTy1aR89JxnZDVBnsCaJq3VhKs/nG8p++9qpoySnTzlWX09Pqm2HrXouvC1m4
Xp8j9LK1liDCCa7KckrEX9Zn6psHvenYB8rzya4caQg2KtsHg9gplDnVDLGdSziEV7zT3zKOJeMM
xp/vrLPBhxq7+h6Teo15YYkMj0ncN/RhttWbhZncFaWnnA8X1RR2hBzl4CIEABJCn0g2ZVchyQkv
eqIWTcRC8uyxzvR6wnRz0HFJx8CX3bNginscXbIa1ag071djrlcnnMRT2sOuyhmvdDzKHEfSDTFe
o+aThmlfXPsxMqh3JVhT4er3hOppworaWT5nVJfOfomN5wAEe/iUndRsEYkC1OiGAOPXfGu5PKmb
829D2obuhN+vrNnr3oPQHGw6GLjxKIbZlX6R7OxkZeUtIn8Pp+PQICUByxnfbEdYjY0I8PMEip2I
JtedD+h7BwGwxEH64HMPqaBlV8PDqRKADyVp2POBPhutQp2gmTfBfdSYlerTI98ORfgRYmQPAgbb
49c78iqJqisW85/K+obVFW3CyG4P+sT/hjyW1+m6mO9MOdQmEX8iharZGDzgE5odr9deAH4VwMAl
l6O2MXBVy+PvPnjeWwP5TnfwJgdSn9zwl4EQPNarMtG4COChxEO7W5NOpvscBeySxDFwvOOk7r3u
c5uYe6WOmD37SnkA3uH69RoVhd8FvZ/UlZaqlM3MqgWISKaoxSpxzIl442Jcf/pIlK2Xb/GZcBlv
MWWftv0QSr4tW60tpVvuVnkm4dTnqL5JMiI3D5lP3sEZMPW21zWOogfQByc+hHnS22eW6StrjLIb
o01nVrnYNQzOb90YVtSLsjQEyW3kCwmAgYeHGw8DaZIBim4SXVKNO3krGw+qO2bqB8uE5zIxn7mp
N7LdTURSqhuxUskEiIidrhwhA9+HvE8HPez3E1lNL+INSIu39LozVzdXW6Fpjlg2BHM7ddUAwsbl
+Gg1yyhzQ1Oxk6upDBVAAtdUvjJktHWnsuXZYXIZm6zmmp/ZKDYmlegOruZVoVCUwz7kdscaIdjl
M9OSCJhcFUhCru8rtnd0WV44AV8zKGfKhPNLVsNKzItbyZZXH6dg95ELIdgjMfC8TW0RSo7EAySj
xBzLDRjQ174AAY2qYGso2masM7P4rzj5C9KSSjaYc42ij6S3yaX7bqP86LAr6G/WkuFfiuGGu5t0
+YdpgQEidkduPWM2QaKAuZrEJW3n29nMk5H90BNVKXbsvNiUVC5KY2gUbC2RqQqxvYJ/Ika02O03
eWx9FCsv/Y8zcdJGODjh/It7f+a9nXBqH6OYCxsZcndmpsttY4loJUWyX+92FR2+XCUKNO4I/0Rw
cTcXthlYvEd3diZBVxgoDbp5a3yRFdBmg8FQqSpbwPRyhJv2el9eEVGWR5nYkbeG4tOVb12NLy2A
2gjjtjj+XNQvMSiW2LArUh8AYZmkPw3IkC+9yYPjqjCRJ2cPN6DLKMUURQXts1V8NA3PhYGYPpju
vk0jJdGtUps4Tj/gVTG5e9tYNL6sca6d/eodGIFsyIpJ+B3D+pbwUppZPcwL33z1i4YM+RNX4sXO
Tq3GKSPCWKHu9ZJnn4cBMyRWRgVofCD+UZexL9E1d7GI43+ECuLya4tw0SmV7zk+STy1+BhbyRiQ
MuJxPYJkASyYO/9fKQdbQbiqVI/aLfCFPvveY8thl4qILRmHVmN6QWz46icrztiqdPXyIWMvRZKJ
F8oJBg5zrC2glpGrBedsQoWTLR9eQb0B/+6iszzi8ECn8oYFGBQP9XUO31fJhudfcDAd6P6ZnMBW
lGTiBsxTI+hGzby6EyiK6dS2WAUF9zSd/310v2ITAaSehELi7MtyKEUxC50zuZ0434yRA7Chg2A9
lnC4wq9gbKcLIkUPMWL0mCSBE9ll4+n6ayLZTG60qpHgPyKQhRaeYkdAqiO0sOsRjAoaCBq61ARh
njRn+wnFJ03FopjmnVFt9TiatGbW01a+Hq43ewNW1rCzilbXS3DSIgOdyrz+XQyX26epYOwkIlaN
HhwFCV4rw0+AjdQajbtW1V3Ev8s1jFKnGKLaJi2+AarxtYv3p2G20h2Cy31reWpy+k7zgglhtoWw
CPUohNFi+jpb2zvOzShNXAax1MWheRWr9k+bFBweg3oZQGUpdKQZj+i+WzgUwPTjfjSd5aFqUAMJ
K0jF8z/1QrXGgLwuZD5CI4LOSs7ru9Y2Anm+KRV0ODCUR1X2nQV86cpDc7tKpNYld8Hq2CAY/pu+
eou83id2mso+i/cz1072uI0azORIsdk4EYizLM/Hn1py+ADjxZKTM8BKOQMia55DyptifTRq1sfc
VggEvoMR4ClMAD7mMSP41RrKV4KL7hu+QtfKaRrVw+1y/qH+iK7maRRsel9CEWa3KnuO0t+3jHVi
3NvdyKM7lEithpsQpgzoRtFHeJcrJSI/N535MKx43cPSsVh1588raX2zCzhwnWUtvOA0ebhcBSJn
x2gCqYYTQtxP9YYZAWCdWAQmbV+DembCllNM4WFVn1bXf/HDUBfOEf09U+RX2bnP7lBcMnXK6AXd
8Y3w/kuoCHT4ht4kiOX+EwUifC742oZlJSbQlbkh/00CrHH8GDcZNynisCUyXfW1UIGDG21XPOa7
g0jlAMQq9EzRZ+FMKPvv3aaZhZh2mqyB+3yzaRNxloAWBPsZa3gdGFReaJMKkZMR71crFx+dPy03
u+2+JklqrENKScL1NxYp6IH8BCo/9S44rYHAHt4mup0uSTZETxbIFtMR6Qwo0V+H1CkoNKplzqfJ
AuRYAjeNd+PcTjhd2Ba08Z795jGxMHKiPDwyN1Fcdvrt3Uj/8dWdETCiw14iTb9N8uBl6N+a+0Xw
Rm0BhyBiMM2L9PDIJorerLJtn8QTXJlsbApDogkYNM7EIWQ2FvhAy81iRVOEqr9+Wvs43cyzKf0i
qFVdxXPGZBvXbdNv/vSHRYfVIhQVxMLa7xhFd9X8A9as1b3Hy9y1zl9dOyOt854JYUc8UI2xpLL5
o2Nk9ZJtwnFRhKRcCl9F9dj+fRqsA2nhaavg1V1bjcGocW+J5Puyj+I7xNz0mA8o0Qz726p5SLGI
bTZKYLSQ/oIen061YU0nciBWB8iUoWWtoIrKiGRcxzEpJVvMUGENohg4NAlLPz6ckRrOSxo/9CeI
bEmsKX3l9TSUh50hVYPmm051YeyCBujHNhUkisr+etygt1DCMbAIvxK3EG6YASTYiZ3P2yFO0eXc
UyESVuXljPjNp31oj6Zt6pEtrgZabwq1JTXl29ZwltV4sl6TXbyTNJonsxppu45z3WhU6Flt0c3r
5+v7byW22FXhpSYuEd0S2qfHdI1usL8LUvk1K2+lQiwGpTMtRGGVVLmbNHKMZ3fK4WKINNOSftWA
gI87PU/OnviK2RXss7j+iya+LDZmF1NTy1qinK90mANLEJRHRcBXV2xNb98Ex+8tkTNgdlBWDSOt
jn4wrB+cfl9sYPJ1TtNkpi7Gfv1MFxmTCst89bNoLdOiNHtrSySxauiiB3BveQFMBMVO4T1seKLJ
p+X6tnuGkGViZJIvFRGd4U4Y7W0FgMOptCANMYS4emmXJgKmq7O9zywnJqTYCiWWrDrRwxCWsTgR
iZf/Wr00oH0u58cx/rr9cNBiQD9G9f882YppK957pNG/hl4rdnJ0G9VKjf0zpSCWwPZkdaY7gi1Q
ZSHXjN2h8kEW8ihArAbKUuJtez+MAQxj9FpvGbiFVdqhhjOS25jdFt8xV+Gnwr8Xo/Z61U0gsh+I
+KEIlmrU8jWGCDIBEgE+yodW+pRbn0SShN9f1KQvDotf6GM2KNpJqP+Jb5P9uDdqTzj2ZmxUzZNc
14XyUhg74+f9BHYS0VAjXiHdA7emq3RnNa0xi+Mwqkt9ZGQRLseYJyIKp1HtsgrFF4mIPQq1zwyb
xZE5IxqrXkB1eBcoGQXsE+vJaeFLFMvAIBAXjbOTjYENQwCXEAVs9Qe0O8jDYWyiF7I7yx8j21vG
IzuWc3noHScrB/EQt9/XcjTNnHu8qoAqNo37nJNBXaBJUKRwYONIRL5D10o5ZI3Sab5FaoeSkhMi
GiFD6mtolSyVCjGOkfhFDo33a7M3pyfl4Cr63L7j2ZcIqR+882PLGWcvxIcOhs48Yc9nUqUw3o88
qWS7yv38kpXAWyDvwsn+W8Ji83aJg0M/zm5R2SJNcb6ffKdT3WDEDR9V+0wEZ82jEKUnc/mK+Pv+
6on9cM3QyQ/o6yPUa1Y6irZD+RAGGCdKuPIcWnM5PF0HHpG1yYzKJeXGj30GOJJMUJKfbvEvM2SU
MM+11BzERIavCjtUsF1nf9KCZwkpRIQ7Jx3xcTOomSyeZpHCG/DY9/7IQABAX6HNs4lMH335dYYB
gvVpA/k9nggIclw94ZfQUCFJ7QLyvwRx8VKd4gCRdLt4EM2qL8HyzNmhsQnCXBULA86HQypRfh1t
8gc/YF8erXwv46+RFz833EA/9k3prWnB0tVHhykJuRmTwyPShAOFZowyc+9y/S2ufyG9fZkjElaJ
5MP1zM4QRa58fFobsdKnWmtBPg9z1BtFzSRMLee/Vk4uArDwfYeld/4XiEofdeFxKDdx9u5xnaRr
wgCGA1E8f3XSx7AeM4Tt7CIoxvULUhlzukZwOJC5R4lFQLwN+vjmIfX1v/t88+rOIRKLjSnHmRE8
nxKOJzq9HPiv4Z60kgiOy3I86T4CK0TPjK6NjrgiwCMf8vkgjy24Gymsm+md5ikxQWTKjr0iEkRH
L4hzEA1tOTIheyLsa0XKCJoMztW4k4cNqaJHyud+aZLaaOVvzZdx7pvdB5Ub5Hu/5snBZGemwna7
YNvhIYyOUt71owThicZbRE+oZwxoBcdPpqd559Jdsk8L4iJHJkZm6bMTaiR4u2DDrIhhtEg0zKUr
MEPQST3iatvP6yXCpcuzUCj/Ps2qpGGzZ88iJIiAYlv5zHIfyRyj5UwRdpGF8GGJJCd3ype1t+SD
4fKBX8kDL6sGVDRtA8POt9x9AGL62RWFErcRH5lAcMnjEQCXcX6O8pPUFYziETuwpwgPihRKXPXd
WCt6Z0ZrB4XNvKItufIJkLKl8bJCRWliINyNF3Wctto7pIps3uey1rkCYmQ8r541nswpmhTsaIVk
VqXZCIEzPZExLLl/RHMxSsicPrmSYhhaOT9cisqZ7NuKGz8XohxpOX6JqTInEIKA8KIjcxSRkx3g
aXiSJhJl8lfAOKi6ywUjPUhjcCH053Fj9kRvSLGZWGMJy6MCq3AC2iRL2WywTzGuoNBBl3Pxu41V
CSoQy5D2Zmvd3OBiZnPk7ZE+llCjENyrJCc09bc8E9+OkWOBglaPNq2kP4WTnG9fOAnlU9IM97l+
/M+x1MvaatqCK+lmLc1lU+/4lZwzlctsuk219FB+1SSVo+RY9BA6kmDLYROtKZz2KHozgZCVIOst
57IfHhU+X4DZS/Pz/gsma734iwVzWDnc5P/xe3RXM2M4aoIwIdH+uW5i9o3UXgfv43knG0foiEg1
xdWd5IkNb04p4acXO15jjMIPjQTzr/XQwLmt9Te04lawjDpf8CNOqwA9094o1ogLG2kTQIDAPkex
YlRpEWcRx34eyBl9ELXflUCfsSHrJuog37oQ2VtJ5Pnuf1o9pUyrilHOGcGVrQ2PpFSHvyuCbpXd
HiVUaDvLSbOP4OHMCAGV9Kz9oSKtZKKPfBs3ETpxSiRYsB+R8aeS9IdjdyPXjGHqPDbqni0ui33V
dyAdoIA5Eo9xahiJfsQ1V2Ns+PGOJq3lxp+4m3izPcREuy5agqd6TP5Mya41HYbdv9xzgKm/4lEs
CO+wmK0cooG+dLRJEYD0nY5C3HzX12dia2DyMHRl9UU9NMvnFxRU588AHyheRIaMVUlB13iwCuKO
dtLmnO7n/ntjp5tv09MvFDt0pE9XhXtJmogRGC2Qtg62FmlD+Xtm8PELlMl7c2kMCfU7ZmyMMrlb
KvDVRgjWQqYf05uEVZ6Oz6abXUsATL3ijXh93XIvor74SFpWqa8DJ4j5IoWaUU6r+wJpv/iMJ75Z
YSCFHo37SVeHgwvXFhuQrtRZHo6O+Pteyfve9CP1qICPQf9Tm2C0FD02EXwauP92wlDMnzw9/oJZ
l49Ag7IzaI4Q01pPkCMGVWx9rjqIzJd9y9zctuHdgpy+51IqAjz2pdlSE1bVWj5qv+PfVAyOuP5D
1qSsJUyCgI6LJv7YQJX7u4re3rqzclN4Dw5COuhceGpMyjjBLFsCS+zkTprR5vk3rdbDennvOju4
HEHu73c6bNiJ9ynh9gh3W+aCbfAhdifwo+3JdWT4Z3xnRK2UXnaWFrbjmrCoN9/dz+24joDobYa9
NmLnL7XK+Rpp159iepBKbW3GqdrJ6oPasLHj3ngivChVJGG9jrwQdKd4oaxxiccqxIriOtGX6dO8
B7T0mfkr3yP6GCd7fi9wIoX6boDXESvr34ZjzIPuHbLNmNIPqENZ9ymrVgPOTni1hIMCt4a71uf7
nTMUgrUcEX+4xzoU/oPINIPfip2IRmLQiLqIEsDd7Od7UOfLpWGhg56tNWc1pQAe8sn6oqIm6vqx
i5ujwkpAgy3jwkYNRSMp4qoptS8KC9ZUop77vdvHeiNUB9YjrY3u96NbSaPjpk+7a/rShZ+Br4Cy
HwjID/aNzIIQECl3lcYPhbSf7mX6OW+qPcBC6nE3CU3rg6T7NJkDtPl77EKki44Z2tqq907gIBAX
42A6LsDCKz7rmi/jo5vmlM25mrsFufhOXn4VVqUuM3nIXVQ0/+sf7U7sXYlpPReeCbFnPTMwDsbD
9LNWXUEQ+NLg++e2blfbLNdRUBehgvkudkKyg8KDGp+DyMxGIu7n0jxiKVOf0u+oEcfgoMynHyb+
QtWEGjjVSH0euFggesGyk4hw4pnCs65mWSvLwXAfhzDTZIAc+Xzjfd0/J5vzWkWPci1Y3iEs7Khp
MZ1f+POza0VSwsBRnkIRWuy+O2GV0WORkTw95c5aUgPSNvDUAXofYdEWBDwzTxJHJT4acQ09uVm1
/9nDiFUiZAFxbZbkDF7pJsQP532AOowVbQwEgUp1OyKFnCH4sqCxSBGZQoVqysQJ4/YC2zC3Whbl
vV0RdZbhDtfHobK7NlRpC7/ruNeRpHuQjNLDcPMFs3uXH2z7UmJKT5KOkM3TeeqTFs8tx2fvqv6l
NhZxhx0fnsK3Y9MmM+x8w1sX6CTlHeJYaC8TX4bHNsEDnt2Wf3MzM0kRUPqp0lkFLVedJmxW9c5a
j93tOUi8aoQ8rG+HVISXITKtCvKN6/SvPokZnX5BKE5SZ/GBrlE/TGOM1cRHr9YomxwX0Djf6dLD
RP4u6CASC/POSQcKHF24sdtamlcbCicx41LJsqpXDLYISxMPgzIF69xu3LEk6C1uBsq8wPTKC567
oMfSSr9H7vQAcPf/5zpm5IgORasMHWiouXo48495wDVSjMcRYjIpWB1OB1zXodJaD5G/cpaWvN1b
5aTillGJ5Udaab1B/rSGG0EQu5iihfkqbv/UMLAlYVvnIhRGcN3oiIC+LuoBkHCvLos/S+o8Udlt
SEH6XFYZBTSANVOvo4mamVHcG0xjrgN8m6OmkA33Px1+4BrALDHcN6T1LJCNX1O+8wVad+hyTR69
LXIT6kxNgQfF6WUUPbJW2zkbnWjzy9GQ9lvJw3wCdV67P44IYCNfc7Pnf078nYur8Szo02P75dX1
GY/9ZHOlFOgd3/DKIn5Ro/V4rV32tWzPRIufwVmIi7s3uzGgnbwoPBg912NRqlggskfxbBkXyEgS
HejixqWi78rHb9IyuVkWrb7/bjK01UvOB5wUHUhZAGDtAS1yPzXQZY/6i8L7eoQ0Yn6LejQxo85U
FqqOF6F9VaVmJfwGSqcgXz2plUQ9QtR6MOMOlUpzsnqfpQkABsUE0zfu+UmJ7KTUm+XzXzSxzsan
8jApcwYB5FfYSA7vMaGlN7f+XtSaLaPTK9olgBqWas7gR0l8uHxzXEjVKLoJoNb9yAQJh1jGtjmy
MKY+LHOp9/Mdg+XL2drMw3olevKJoiLes8FbeJtD20lGzY6MhH6xMHZjXTGFGEe0QhYLZRvxMdeF
qq/YnY5qvl7ysNK2jlg+etV6pR1GU8NRj2Jpss+ekrlsx4wWyrIX3Wn1Vtm9nBic5EtpA3wf+1sm
NvC2H5whI7RbMIH1+GhxmOOAoMuMHfPW0n84TOJSf3JiibdxvxZ+rJSedwgaX02WXcG+7L/Sdg70
FYYtUDd97co14aXVfT0xVtyiBW7k/MNsfhbNrwWq+7y8uW4F5BxwxPhnEuHY818F6fyy49fcFbgc
MgRQHqvxKrjwTLsYD59Feb4Nt6ny89zVfNbqx0bj/aR9ImqIZA98C41+PwgMplZzyhF99OV82jz3
DYwSTMXfulLy9PUFfNl2c4IZNIqcKM/ECa3HvakGg9d8R+5jnFT3a9rMJRmxG8r8qCfMPsW24wGe
t6nGJ3zEcwNOFCO6RShZXWRzdUZFWsPoVA24KCLirtcvNQYnDaT75d/obu/oI1FdPCJIki5u9SWA
V7amUc2qcl3c0jHOYiLDg5JOFLXlp8C0gkn0NlCU3hWqhnHIOXlTrSj1LTFIDHAA8phw4X4KtGr6
H8AfjxNsmg7WFyTriSQHOXE7icOUYYQqOeCcY1iCCPrA1AgdPq47NXM/F+wmNYnNMwIFJDjrFH4R
uSDnArCBBAHEediZXx6TpIXQKKkwfEHz2EcS6ysLctLlPHGi4/sCmJdjbnHOFbwvhCbixEgvZJ26
IF69VaTaYAmd4Vz8w2YP/1OfV+eGkya/QRoGGHLEfRg3iZpLkTmYdyg/r9V6AuT6aGX/Bu4QQWBL
l41MICmT3IIzgLVt1Qr3bt4rf37xN4SAKFtVzIc+YUAOqh/Im2X9SbEHnJemWay+olUE6bkz7Liu
oA6cx4mOMBrjcgyBVob1o4H4TBYRkjJF3C0lo/wdJ412WK6WXhSDb6gMGtfLWumYnz06DD9yvxBp
bS/R/BzJhYcQBadwGt75ICnjGxcKQHJxhvsLguRvU5ub0vZm8o6n+stvuKTUGTttiz+6hinmGKe/
PuTGK0KIgWBiu6RPxNXKtas2izawChSEHuJgIpgAW08kXy9fe7xZoUmsy4Ccep43+XsZyOFQtWCi
qjVNEYFTrUG6+lEfyFheyk2mGY7mLBnh3TImvKZ48Jz72VmG/GifeiyreUHG3nJ30cYJt1kVytx7
fwcXdhDWZdkYDs9ilPkfFPoZB2joNmtwvSavZPPaTnm/lmnJdvzK3NYDHVIjC+ve1z5U8ZbalWSq
eXKzonhexoP4yqeo7iV8Y+QDcdEsrs/anp8Rm0gvdmmMmATf38QQjapOSKjYoRQAYvtdbkBt9B9Q
8a699XLQQIfU+zdDNGmgVxBsryUfH9WpZZvdvZ29mWV7e+NBkFYPcHqmFypHGZOysVIWWMWIUFzx
sN+vX2OKsFCC71uY+CbcPM356W/nRP0+aO/FMJqe0yepguZs6qnwbQ5h8p3+l1th684SvdqWeMgP
UJz0nkwTTbPP+aojgy1SMpsiiyCYpeWoAosUWIScArb8iZTGzFxDn+U54di9AZmD6mXOvI/YH/fD
ak7QRuPJL38EVTuQhhrqMfVONzkG3sh7XitP5NL2fXCywIWPhLgqT4iSWBwAZipdrnCYmt7OL7Yc
moIFufgtA2PozeYLVLwPfaWLZaOIgi0tPe7PW7xP6XER9noi80Q3uMJz6GX9T4323LdxuRGdw2tB
55m/dwpTjF/trlxrYSy91OtWZKD/IBghTzCyXtWnFL3jdDau6k20Acpb+hkg4r0NQsN7Fe4kH7my
+0VcC0NbxjeVnELipLtv9iioic/T3EXky71dLSa8QEZtyU+59ToCc7/2VZwBnEf6+XlXHt2eJZNU
C512/H1lqMmAvObIEnJUW9yUJ/Lw4cpjwU0YK1BJ1v2C0+/5X+4qJtHhQd+hKfrtX5zdMCDnGDrm
YaZvovyBtifwu/RK8X70fV3b6DsIq80YWzhP6Cj004cvcExZ8MC0FVZDi0HgqNuGSX9BmSDnGbjG
nIa1KXLsY2YIKMqWqQUsKjrW+KeFSbWkgT0NExstMILmau4SyAWbgMsiIOFEq+6irx20jeBFW+u+
fX8OYpAw6H7nRkEp+LcmAnWaLJ6kNLBkromNagT4JMSMcTqeYUgkdxBnA1BlyPWOgmoO7BqPKyEf
3SdK88b+O/QKWSgS4BcRWnerHY2jtgqZJtmsRJFUFujVdRxzc2WuGcgf3lZwGb5U8IBz+ZP0npra
UCQXM5wskcjztFVgur3xZonmRpI6FdVap99BgtA8pfamFPaxHwRGiguhAHgLLlhYBQaF0Y1eiGsc
oRyi8Cc4StT6G2GbMe30hMXLKVlhwXnN/vvFyjkxxElJ7CZ6yOmkUfZGt5tqNqvbFNM9JiS7GqZv
9K+qix1KzYGeo1hdKQvLB8VO4qZ0JTo97l05Hyga88apcsxt+hfswjwv5jaoLdqUkZXRXaS+YpLK
QjbeDFwOBZXD75/JLpnpt0zGiUbLOJ25WIRSwyzP47tYH8QKRD7TbLn37TOboARF227M5xVHkDNd
TwmhaRihypJgCA3oi/NZRUnf5ioDFuDLphY1Z33f1mUdz3ScwLGabJ7ZpPeEysF8n/JQcCvbHJhD
eZMZLgKAa3XM3IOo2dCIThSjwch+TNOTppq1pdkYI4fGdkVA0RKaYQHGGZo2qeD2UFW/EW6GnkO5
QlBjVFyepEmAQtGWIwxS3PouQL8pc7Ml8UyVYDY1pyl+vyYyjYFlWaQJDqDHBNZoUDqE7Do6UHL+
wOYf9f3pdFUVIZKThHVDJsN3L02Wa/xkw/HKdbu7hhazsOuBVFyTmgApbgsgUP5e4eycTWIQoWro
2ro12atvt3lGIqifMki9U1+DGLS0YBS95+hxPFgIS6ZHWMSHY7gkqOJZtmiHbqVrfAzqeZ96HNND
djXcUmfDSbSt3fC2598qL/USsSW24DtUotJ156LQrhqlba3ywwxHtKIsZ43hIlLt1e9aQEh9ocUc
NR4uTKeiTysVk2DKIVwdOxq6Gk/W73dcJkSHmTlbHjrWL8Gp3n9UIbxhiGv3CIJFxXP+v9+akRdH
rJn3UM0bNpSREjWn13bqgaWGbWR/Q/YM82tmOn8vEWBeHQeoAaM1Z7Shih3Nk5m2Oge/MvRz8KMW
W4IhTZyqJ93TeENcsO0v6ES20JhBTj4Gw3JfZQz/ddFRo16wcy/xH9T+h2kznkY/XfCfcLKTRScw
jxa5o5fz10I12wM79/f+H9u3h8FqnSVcSS034qIrqvsd4GOfBfelhS/X8jtLKFAUY022Sgtojsfv
M3X9lhdlyM9VQdLhMzM1QNTNBJA4A9RO2JfR+UvU1HkWub9fqqMRk1LMLq+cLbo4WY6gJ6dnn9Y+
wW/nDGy5eLPjSyUxij3ELbegyCrX3FmRdeZbBE0zIhMPGoGgLhWjkjUYeaosIUUg6jq7WUoWYM4T
W5mZm+H56CCJP5n34MzReRt1pFCLLIG2AZ+12de02FIcvvauBuvpNjnlxcfxQq/rH1Zf1U3yjBu6
pPVMDDutII2Zn65ZEuvWJnv4+lIMElf27k70dmM1bObXLoTipr69+eVPMeLW7hQ2L71oPxvP/WzS
lLjDr3Zvu4OYoPC4Ttgw/epFvFYZQgyh7Hv+GRm6ltMeyPZVDWwJ9h9btjS2FSToJPU/sE3ZVmBU
tUmPWfah1ilfhNm9xd/1QiyZoeL26nZYXmo7RLE+O9ky7n4N2HWTfMSWzyiZtQBtrQqEvdWidOQn
fYxB1c7a3tq71MV5oN4Rdllzn+0no6slu34q9b+Md/Nz2C7EpIFKg5vsOLfFayCSLrEB1wJ4o+GQ
7C8lZosk+4E8cmNNENxYfZBgvYmaKrijh7CeDjKmjdqFbhfE1iWaHRycdeXLZtBgHML8I7m4WsW2
y8cPR0pw/cySkf96MhpIH8zJLEKKsqLyryhTN7ruWMDc+defrKeZDGatlAavR/Kv87v/SiFDRC4w
c+nmZDBuzDwd71REMLfzJOotZu8PKgR+SEkmPuavGNH067XAJG3cdXNFrFAE4f6rpmsnZPM5WH2/
JuKLkUBM1/awLDkFKp5WxgJ/hPlF5zgZPlJFL/hnlFuh8OaGbcOF8tY5CWzsEgERq4ZVmqP8ohmB
ysLSadIjjXxT9UiZ+V4NqqVAD2XZc96GpiSHStgSkYm8q3r2qNRuNQ/PsmgnkbGaHqRa23OMsmMD
SbDe3/9XuryLbo8f7yyQcgJ18HaxbIbe5r38m7V8HMSxznIosR3PQHozRKgnjqrat41TAmmXoquy
d9OLyyT0dKa15MYrGIBU/N6C3KNLHJsqViC1L867d2ERVjwr0wRR8DipcTqFBBhuKfsLzXdD5oNB
wgkN/wsCucz7gWytXhQG9Xp81Fu8bOj9kpzLcSrTiuxjGZjAyiH4zsFNzIOEATO+exPUjPRUoIma
4Ch8oMQwRP6iz6BUNz3TRbw9PTfCMEULgUz96FQ8BTjlzvL/AbA8dn9ykFjawN7VciwLviQRp4Ei
iinL8Qgzg+n4LxOHxvGgLsO8krKitKgKa9nFCFn0Keuvrk9fQNQePd/6u53zR2d76YbrCFmi/xeP
wHw4rmC1Ap0o9h+5XaFdMrKJEYIqAAC2Q1z2NvNjPXuSxOw3FIp8R9v8GqZ3hSS6c3aM9vuEtVjh
zayG09dJeeRYvmGX6IUsbBueL+hLJS1KovhsaE1LxUrZmlr7iQxVxdUQJyCVmCzi8d43zMpmmSus
psnwnuIUnTCfrd9ct9kFZD4sZCw9oOy59aW7txNOHMw4tNP6xIXlMeTqURUEhrqckaF+3Q+QQ52m
oEIgbVXdnOiI2Kz0XPMLQYYTR9IxpsL/EsoEXky32trtPsCkS32h2rOn1JrwBWPkq9DbM44827SD
sns6cSMgKj/oWn5LF5ZHWba652w03QL8sO/5aCLTSFCapXK98mP8eOtTsxXKHiNgGrrT78fvw7mr
BKpT4N9UfHvn8c+Jw7sIrgnM1I63OH+MT8VxWpEq1r9XxCvco//QqaXRbQtdAklJxxl7YW96xJ8L
cnBNWT5OgpdZwQix5G81hUUwqGP7LhVm2JvFD/n37Dfruex3WSjd+gFH6mKvLqKKeanepRmQRKS5
DB9VXcqux0krb9DmacYGFt4FFiaM/jtpa8OCkOjyqw3dB3gfsPzTV/xTdmFfVu0QPzKpNkE5P0v9
GyCdUtBXLdX7VQXWOlRIGsO07hxCLc5x6MiDQNzuM1Fw7WsgS8DBCdEdLtGNo+5h1R4sZYyTNyWG
IF9ZFB/qZhnQJp+p2uFLX+FnvoIRKLJW3en+3APq5VSHEfrJRxU0LGzfnA2eRfJxGBp+YawOJ52n
NKXBtIydWzybm7qxrUjacfvAODzvWlTYnUBB+7aIu0mo7nZQxYh8l+iupSQOys53qI44nMdRRk3h
CQJ+cBb4G47DRK/A7mYMO3Z1y+yJV/1O1jRxTCZNqpLOAqoBKXkAFmk2dkZ0yfnJCLbyhxK5HYaR
IosMHvkMPdbaySkJIZ62A9N/RDnp8SPeftMGzW5NOhqOPJ9+CwmXDlkU2jXNx7BGkc7WQGXPIVw2
L6FXNvz0pHd8zWRZ3p4WV3oOlwblqPGkBzCqyB8Aj6DVMCdnW11GLqr/tupClHsSQoLzdf9BEXJe
oqfRNzyjiyRPGAULJap3dOmF5TpkMzCSDoJ6ZLjA6bkcl3C5cSWYBrH3m2QUn2zWDhEOBCMFfpqG
xj3s6fgL9ZcLQb7kL+a1W8CGOVYaFi+GfhveLTAEUR+/CkozZzGBdFj/G4ijsuyde7eleAcDnRBu
6rbDcMoUlm7LmAGym5/52uFTyQSekjg4GR8ZGAzc0zWDzIH8eYIGzgEP5Spo9GlOvsqJFnLbJhQB
VWxVRlAa8dvMUobnSqLf/d35Gu17GaB2ixo60ixZIhvB7QIQyuaEm+72sB6njZvHPtRUIKC6AoAs
z753oL398CnLFj3KmAa9WKu3ziLcsyhoZaenyikoerhJGQ9BmFprmGBHjFvrQRWDNZ+/z+2JC9Mi
3AKb+sYnndPWAGIjy+0tkBSm2Ik9Ziix1tg1mhlZe5ioSYNN2Ok47ei5IxGBUfMMeL/0R8pr4YC8
mH72Mx47tvtJ148ATXQZCAAaZiqVzD+0hwBwNn/WjhvzdBbWvKGdmWXIuaSOMvhYQRb5/Q0XOqcz
ilvFjOCDCPolnYYLyp4RClitMx912NLQ+SDB13I3IVDxzRpNvkPDpXEP9lDDWo6nSLbaGgLjWx1e
XKLfSwhNl9ya9itvQkWwoQu2+aH0Y5lKU6KGzaoyQbfN+EuqkEkASZNQteR3gSe6bMajEUhJErPf
yDWgewvSSuQoXayBTcylkEDMLKsXUgBTqs3mEpYoeCEUpyLJs6DpEvSI2+fXudrvAmYXOKuPGPVJ
mGygIZ2lmVCB2ApjlL3uEsY4uTCuu1+TWXNuS+tzopC6+AE4Dz/XbgvidIhDLhxecFMVuEZs3aX8
LJ2293dlPVs5x1b64GNTojAvQ5MYNL/9iX1jzEpo3hDgmK6leA/sN+RXvgHXq7npVsG48GrJhkYM
g4OWDrtOLGQ6p4ISKIG7dM0zjDtFILjig+q2HYLAZHrqSCrnrtHPD7vZwG97gVANebMukeuSJcmF
Cd0JAfDsIuty0IpEXACVZuBhp8k78GGhQT4da1PA/fZJcOs5iBA9K5Mw97KK5py7KpvxmUR06qkq
kC2QLvlyHlbQRFdg1FfaGWqCY9l+B9OMpoeOxj84WqGHq/TsqW4uXl6/ttAi855SWpezAsjEaBrU
YGzxk2CFuX7kcIL1qsKkTagxR7+FqpKnbHPiD0fPXPZLrI+B2ecQ/0qJj9HqmRkl0QcQyMs7Bs3P
llWEi0Oa+Arlk2RYWEJIq7sdc4QXD7/QfjNTNrgTEihJCt5cHYQc2SxNv9MITym8g3AwxoGiLsgq
1j9KVqhdg52dbeJfmyBY2PCIRUm+GAAsungiBnlVYjnl9uA5szhHpnZsZFG6Wvcy7SPZV6M6IiDY
c6IUaFzDc6OpSwcG0dEtljHbv9J2ClJavYh0MGW1goXIdh3MQ2LPzLZH4M5uDKSgQieFi89TpSKj
HPAuBTK3d7uumgWko/tIxIiJuELJqk4DJcli+I1+JyKi0QPzYCvjOY9M8kZoeNbSUJVK6UWoDAY9
Mz4QF9UpDCsxJXUqsbN5Sem1/YjvDfP0ayrugEWdJLu8I5yJ/ehCJ5kBWJpceoSwIKmiedmyL/tR
fpgUHBKiDubeefmg++667vO5nbeVhEcwtVi/yZWo4+Qhb7vqitqsv71DXGCrco6gj8KAashLIHVC
bwEMKUzkaipR9jAgtKlko+GX5ljH2Em6iYgqrxAGZeGg+GPomtX++dNJkqwKrMvyup/e4C6awCGT
57O9PNmxVXfUdFdD61NMz+djawws0x5jsZBAMg6X43t9CrxrwJbRJMKfRhX4y3Ghz//bhCVvrSC1
Stz0qanZsBDDmpgmp2KwAogA2/nHkzSmlNOVmfDNMfOYFKzJlwqUvnYIxSp1wky5614Ab4xrDOPF
iDOnQHl5MypYCa358mz7DoGBWxql1mv0AieSh2C+YLF7kOZrd49E7RKR49+SVPHTJn6HjoW1BiMx
9+gNBNHczLb4tI1ms8OxBdgf/xRh5kQfCgfSgzU2pb7B3jP62aNeINV/NCwN76FYVclcXSQ4vxZT
AYMTMR+iAlglOZ+m3xffVFOSor/CS2gyN8KIlSAB9kJ65tBOlHjegwpc7njtyomTF3E8C83CFdBr
WmAZ6Vzsy9UeSptZNujlGHWpyNafuR8f6gCewR2YImHM7qt2Tij3lPotEV/hcUv76BCjX1vhCKTk
3InN3WpQEKm8MiSEMauXtOjugAIxaenz91nUQPjW7Uhdv/8mByNbGfJ3CWKt6Yq06BTZ6CfBInPr
aX7QRKn5JHKAAPvCewxxPmlTQRvNvsV1Yjm++GejEd4NJj5hx73xk4eRaXy2PBH1CWKxHLnnAzve
JDfjK/duMIDCBVcBp8AOZ2cSGxPXD4q3LSE16qGPboTFAkJsolF5geJf5aDJsDQcfCjMKCn+ggSv
un2S1X0vMRXnC+NQfQVvvJj2Z2P9dS6fiU9O6s7w2Alnnlc7y9+KqI0k7g8wwVai6KozpoA0FcgB
cFIuSMYWFWqpuDXkU00v4WdZPWvnjsGUUBPZvTKl2AzLhxHRgfd4J7fTtAhwqQPjCG5rdlhVkKan
maIkfby+xXGq1SrxIbykq1uSVgHIMcsOzV0wpl+xjFwA0Q4V/CkTRjz66Ic4ZJehGfVvNylU14Zw
GMSHbEaIgmH420qLpqApzpg8Pmx46Zem704OyXSB1g9aQ5Ghjo6Qcp/8WnxcPjDJ2sUqPAyy2fqk
V2XorvsPDK83q2pkI892CuuEQYiN6ZXaRTHo2wv2YfrAAf8YxyjyHrsYVA+0eETkbgCimhUbbunW
T/LegKVI70PM0yW+jJURKk+uRiVsE+Kb6QYazOKC/IFBtmMGNr6es4qzhND163TKoOPX2B60roYv
CmArm8fPyRxWzICpU2yjdJZ/veWGpQg2aOufCdDcgTroMPzcC/GEXd4WelnD4pCrIBSUXjCx13Ar
Y1siq+Xn6JwSqu7L1Ag9poZcyeZL7LmZ3+5CKtGPA7NeAZmdbc1laX/s/m9jc5z5Zp9WI7mNFaBL
L1Fi3kEUNAfG6azKf0z4okZwXivKNkK+bR3mHrKaUYsvTmBwaX5fmfJCgBIfau59YJ8g+D2WeU1X
Cu6GpfKNCGXDSKOUUTsyw3H6IbA8XyPrakewA4byJ7rfXA6jF/Z5B2QM3afyKMqU4kf5zqXJ0Yxz
YTtXQ7d6rkhVy4+2aYokgtdp/m4AE1FaGHCB2LafhMPSD6KHqTLe4xQuB86KDIx/ovh7pdo9Gmb+
+0Fz10rGOme6fdOmOlg3stBOu7w2aAvupx49utz1PYBaHFcCwOxzgnOsqt5cjflevgfPVcrplqZE
1I4x/cwYScszoaG1t0n1bxxe0I8MaZzmQGwPPAivdOs37Sv67maM5Q9LaliMKIo34U7IXNP0hMac
M9MCnmk0nLzwhUAKMG7buwGALhfU9i/Tb/v0rCU/RPtNq7z/Vb1xlCCdEG//DG8NYDIU5pvvCdgU
BPOFje1F7JEDYpzR/MXIqhe8JIk9G2QNm2PL2RG6C3Ihf1lxSSNIHY2xx26hYGb12laIK+gCeR4n
a1xsemGQCSnUA8TDvVGu5Lf9qvbXG1bRUEjOBPFuIGNuwcIKmvK1h7sTMAuoRuKzdII5z2/uqxdo
/4H9zfmsD6HhVIb62NA+7gmmOvPXYpfj4BFG6I7U5YkbOkFwFh6IB9VOMkV7WM3rXuZY3Pr2cmoV
Rdl/n3b59w4EBF3ioSQGRgVeRp0ok84p9Yb8KDOV7plE83wnWqjBvrI2QW0A2djedm/BsoNRnXyK
WYrlaVfED3tuHm3UcwvIKsglRSgboDCcCh62KiOKIde5sNqeck+93NdEGnCFHXp48mTVwm6VpQTC
BDIXPujSbGoGcdITKzYAyQYm6VZUSBYyo6/2h/tiY+i/aVwvqB66wz6yjh1/rGHDNP12eaeyyv+w
YNGVygqWWyNkKk25P7fD9LrnATHMzwpAgROzbW37jYAqeWl3wkCSy1Aw3abe74Izcv39LbSs8vuH
z8GVFBkHIpi0eZrInnRQGhWTsDuwuphcO+qrShTdsGRRSjc6WGNAvsbMsy3rGhS9kUmylWdLriNN
afDS48CHzPPtfZF4Ed+GG7FJuuuZrpVUJiOFiRp3cecBu1kQkoUGCsxFM1JtG6GtpNDL+P/gD/Xy
EVi5LPohzSb5KCU64ODwtk9+WViv81wvewqIRhBeoxMU6qCzDCz9DN4FK4qlBSPkTFS26bN+mmp1
/YPwDb8DDrLWSKWu3YcLeCoGaeiJRZNGqiHsUCeaNSrsuooop3D5pXi0qBd6GGGPqjhWo8Fba6y1
nrXNtNIhd/JT2LIfTq51p+T2rYT29KtODhx0tT5v0qUckivhe8DUQnXfDfqLLdV5n1i62OnexYjK
yNptnmi+bYFqF++5VIFUSDDEGH3ZkXqx9RlDR0odaz0y1/WAHLCwKM4JQvfq5upRFH7ij8J1chtB
d9ZsIB7ZtLm457M9dzm6cKKRtuA6o2+tHnmCu4i4ec878MwfuUzEWEuwG33JGTtIu9VYbHUxQyz8
wnIH9I+YmMwAFsf++F0Dz2m9Bmyw0ho9kBT++us+09WNn3Y0c2kX3S1t+Ut2173DXMXrAMgvh1sU
QpnqWEzmziSGaVQjd0UQUWEFwVwJtCYALEW91RtOJgfCKW7mSvtziPaanPf1Zt49LW56b29z4ORA
i7YDSG4lK/NjTfPUJfCdRlWdJvTUJJ/fwM5OEWAAJQyo7irDwPzY5Eod25sAOgJ7mIEhCbRv1u7O
0VIe3j7zijxsLOjq8GTh159IKqfdKmYDD1wATpYJsLk1mlRUtzl+86Zc49Y7j7pjuon4MDimr4TH
V2e3lD3R/FbunIYBRimqTcqm1fCraTqHGiI5i4skpTwHczCy+Cc1CiF6arWfniT5TK1KAU3I7TY4
Rk8+V/JL9/5EAhqMZJe5BYvRb6IZxAD62yxxVzANJ+8RUJhm0e43IY2dLjQ/TM5v7cANR5HPsP8z
PAX18gXqB+QXz03ObrWW9bCBFwVakeN+WxQt/bT+83zuNTWdKR+B2xQroY+MR+9q+qTyorpVM/21
QmPzFGSFqnHF0chcM8uoTh+UaxUkHrNb50YtHYhmvnzNrCa0nTosFZU0Z+o/VnG4Oo8JZ9qntwAX
Qlbp/Q91L8ADa23uAKjHleJOUKaFKW5ZCq/WvdQnMWq5ZV0eqMeoHMcBCrKARu+O6xVVBB1yZNnQ
l0znAkGnJe7NNpGJtE3H2X68jU197cByYWpdXIiCAjLrJ66AuxMb0YaB4pgIEPaRavH1sSc8rsVs
Nh3BJ91QNN73ZQoazM7HMEwdhTraFToXdFE0PatQNzUURq54VB5endbGQgO5BehuUV9dw0XAQD8E
+P6j+KjrvyyxnGvkF3ihJU3xppg3RPeM4XXlw0XlbTDjy5J9tJ8emyGLKycFnM5b2Iv/ih1BlWGt
LXiPP2o0vbTiMPvU9mCz8opfU4BBs+Bwic/QCmgfuVqlxemc+1oR7F52nObos/jbIfjU8qZyTv/7
yv9AreB+WZFPypF2kqoxgRGaU7ICAMe7lHMdHJwav/8DFD7qfd9B+W3qereTq0N0Sm9X4KK9Kg3C
APbWzSMKtT8vXVCfedRARlFY4YgL1zyzHDIVpgtkgEaXRBgrx9cfF+JYoiGcang+blJFEywvxlP1
jeVQg3eUq5n7cxXZ1fYMXlUYdQriifglpgibS9Sumgaw7qliJUJgZNmwZdsQnBeBc4yPKDzs6NUp
RMQpSpfl87Mj7zbRrzswWuEwklGh+PtSXWEGHDBApSebM0KpOFbXaAK9dLsBOOljZIAqnK+IcJtX
5AbY2fKTi1jsE4ZQt0adi8BAbx6JMxl4iPIxQcYjuwr7iRnotSVfuvvre6C7w48tk4eysNv7YL/K
XnRvuboC9wwNFwr+CeDEElYDOsBdeEXP97ynYjY/N0uavhQY7I6kvq4DD2OLLM4uCVXGzxnYrtgv
KNyJid8xcROywQfChgGwlnqgr0rp/pASEzpPd/rr9Lzp7eWMluuOcl7BdV88DFGFe+1x99jBWtqn
7bGkanTYcFShpQjQ0kJSMDCV5kSC/Sc0FqyjnUQ87bxWKuSGn88mGOF3fUoLhUHzAf+0jeE3EsCS
/YDzghg2rIW9wvuNj4MNVADcZUKQfORT4IpL0NTwLrZU9nBafSVWGaZn1z58p+jfuYr/LqsgfgK4
3jDsOECP9aErxTcYWQpJra9va1tlaf31rxnSqawF0JnR5zYhGHJk5lNhE3rGYKc8T1E7hBWt3BBW
84EajrhTDdtK1LwKVsfPRPp9u9g0iz6V+15GTTFOYkIO2EKzoWylwOWMEvPkrIjbnkeL4h5NnTTn
EoMXScp536+X87ERx6SY0cNS0imcVoZ60ahkTG+FVklDRqz6fRxCeOrEnOmPigLij8j9rKT0LOVg
9DlIQiAt9XulZkOLvGELU2S4RckIJsx6xVtJWh5DNJoBjTvLVO5ZOkYBzraSz3VRv7IlZRMkMBoc
6W/I5vg6HwSMlv4FjxzwY16VZ/jbCyr+T1mJfDDj5yMQhO/fgAF4UWojHrYs6dDoyYxIiYFDaBjj
b5MD7/SIGW5angWUNy8166UporfTxb9CF8na0kSNAlK/nDB/yWVYIE7MkIPl/ljNT6T35wU4b70E
XCpH8H7VwA0TUZm9W+IVcBbWkDjp8MWG0L+AptpsY/DzWjFB3rKpgwBWWvo+E8YL6nYnsYA2GdPm
FgfF/Y2mURWyOCSVG+IO+RJmLWdXk+rNO6N8ENnHVP63npCuRHDh+/JcYKazJxLe/KLU1MocKStd
GHIiL21y9UCN3NsA5izzGxUeX6Dp0mL8k4TXni0DVGPajqUSd/bI4VhvjJ1y/6thkFKZeQERTIJ0
d9n/eexuQVnomfaCfn+jc9mQe252p4x0xJNM79t3uqYm7u09P5qfs+z3X6MVEArOrBy3pDkPNuUL
Ss18dpbMx1ounefqyB/GwGndp8zV2mYy0AgWA3yNNjhXeI28qdwHeU9atkMUIpaCzPGkP7ITJKbk
8Q83PQZZxtWi7DmLDEaCAXTCf55r1BgrzPxCh4WgjxTObS9QjvlM3UM0Hs+eZ4gSdTDHVkWsPEQt
Vmcmehah16mMCUftybBMzGAxVOrgkXbbFYvYr1dYSA5WGGbyCp8cH5jaZBa6TTkcnymFYlN8etwH
o1ZBB1hOlj9wcpk/h5P7oufMXVCub8TA+Iz/DsNkSoPsgZTh82EzZcGxADBcEHoKrv9HhuOsw33M
6BV4/nVXtOiZNX9cmcYUhvt0Wo2nRhP5BINV93o9p8CBZJUxSSQmqyftBSWtqGZ+2plVHt7SRhLw
PS32gBUwpXmB0N26Pl3VWPlEdqQJclH6AKEye/RTT4Hfy5KjTVirf7lZuR6mugW5WxATWJoDfb35
VB8WOtkd8+VamuiYLUiakqIhSYBQL1q9+B9Hi3zJ4deFT0DgETpuO4xs7i7L9SFym5cSpV2b2EH4
vp/83vsMyB9Tue35x3q2CkiB8RNVvHIW0Poo79eNZ/P325OuWApdjIoZo8oBa17eskBGkXZqXJbn
uznPmqQtfL8qJqhXqk6za6gbu2//W5e0QOdZRr86T4SSvOLIj8WKQ5IRDqh9VI0f00on6YNolFsp
FSdY5TdX/zh8oEwyDnGXkf8aqQCsjlf5X8bZMeSGqiOYfiZ02PvvTIEqVSA3EZf9T1POFJ7DRBYB
Ul3Wm1aWCRlOytXQktctf22ExIXaxLEFKv4qE9CP+yJkTAdfwHrPLmhV1N6GsZkiTFnqAUyFQNPF
4ueO+RpDSpiegy15z+fNeM4spAZgD757k5+xtibJz1v85RzEJVTsPKfF9P13e7mZ9agj/sFffAUs
RxaTCUVF5cmUacyzPOOc0MhT+AXL61wt/TQF/oYYjTYjiL+CWapCYzLJDYYdCRuFqc9Ext4dPGud
Os+wBe5sjORVfGbO3SpAu09Ix+jaCNeM6sdfFEkLE+vB5M6+/eWevdLykETGVl7OAH1+S3rmcsBz
lz6xGvcuRQl3VxGY2IsfXqohR52Zals4+1ds7+4WoxnXS1znEJhVkhpo54/W8ntqBUOHjZ51p0eI
aaQbliJ6T6raRvuiNjE6XBBZyIKPz5ktlsRszaXX+OSHLVM8iGYrzG+qHRQ03bc4CQ/isbntO4ZB
Xvdn5ecjGpqe+75oRDPSj6KMEDq9brECjnt5SXmuTWQZtzSwO8GYqgKK/w24YgjMhTlaUnEMQ0O4
2ivxrIIQ7zI2VrENzLa/6uSSRjM5EqnjWSEsNq6SyTicOvbV+V526gF3EgvS8VddFD6/mrcOq4wn
4mLwbOpsWkqOUHxW0y5Pv3PmvKd6uLpzJuel9yISFQzZXL4Ps/1uYdCl1W1hr7apefihba6JIZ5w
CsFUwWU0pR6eyuHwmO6I3aVmuBh7Gp81iT3TOv5Z8Xx/PdnkvU1L0zt5iQHEUvCRQAxg+2xPoV0y
NC4NjHs/pvMY2gPGUnPQSUsj95Pww2faBzphb+ynFPfXAFvkoVc0XcW6xlbznpnh8g0Atl94lLT7
wIY026MOvKRYu2rF0tEK3WKABzxO4danB+98o+GrMlxq0xPpwH2YoiAE5Qr5esYfB4n71pXR8NeH
2YUKObbBYWvcdu5Ov/jpllCjn1slurTD0ryQqnR7HDigbGOWlDd4T2KoewjypxlShV8UumbBmhTC
AmZ5AjbAGv8/dSgVlcRnbRO9KrFoZ0936thc+Q2mKx4w4UyGAqQ/x5/P+AT6MlnNgiz+CHHbzOWU
0UKK6Q06D2OJevSVy+iWa2cRMSLsENVarIrEd3C/grm4u47Nw3TDrcCWhOggGuKpXhQLtXfhYkls
fRP7vP+Wq/ri3Az1hHNDcaKXUDiIbJKg6SIzaBKkbvDlZbsz5U4jllDWEcVFZrIvNRIvx7Z21PV4
JVHVSf2KaSDyrZmr/POUXMyhAw0aUUlk2/wOEbbvEbgwNXyCaF6PmkIQVy72aC+K2Wf20BOCP2VL
GbpuaxXcEllusuGKZOUal5p2sW3598Ee1PifoY6/SylrmyO95x+ISrbJ9D6IwGd+Q/tNIE5SkS+6
Hofui+0irVS18yWrbUnJYnD/SOnnSxhovHncnXHGzHpUyseI3cwo6SCJNCM5btohXMmqDwUzyHzq
dowYfQclnKW2wUNoYCvCWq2shTQVxhzB5At2w4aWlNn8QBKaQ8A7HBOCfTP9TnYa3ulrmW4yxig0
rZ+dhmo4Np4KJ8RKvnNoYLlDdkG5dpFWKAHjuweQkUFRjqVXmP0OET37nRnzaChOfiCDyL3A3Lbg
Tb6YY4xYuNVYdqf9M1YDabdkEa173oyxusfNbL+CXUgv0GL4cytc0Q4rFY1k9hED4w3grtDcAf/x
IpEWd5UIHJGZ4TRKHXAMls0ooIBFaNMJJoqmg6NmDPbuBXrmwVHDn+AZVgDdOkV/lRGjUcGAuAsg
zEfzLpTwEhrfTTRR59H5ZA5js9pzmDQMl1HipSu5Kfv4PujrZvb3A7tOhKXKwNkdX39piyepeknD
JDAkWbtpYETWa9PtKO8IL/maPCpt5Lam0gUajb9eCQD7ASSwo4qVVWs8w4xo+uP/Z1/Zb+fTGci+
+CkDiNyIVxKyrMXfTwx+Y/fXpawS87C7XJECBgcUf1yqyMWyrneLL9RhOkkq92uKuLJM5TxcWJ3B
jyS5cfpEtzW0nBxNC2L5UqzU16Q3Rht6SO0FJIZwcWobPtOldhCBpX3And4MnsshL/HwmzAegCgL
7UJ45V609BKXZhPNo58GRwPamBckX5+AxDkIsEHv7IbIi/0myrYw6mmJQCj5iNDscRfRRPp8k94M
NbmT35aFF7oTMNjOrzhnYIh3lcr2FKf0Ewkdb+nbaqj+xlx0uUdJoD4x7HbFgtuKKSKOH4TIUKuD
sbReCRK7B28g5h/W4dcL+BOzHMCX57aoI5WY/WjBqtjwzxbyzgH7u45BfFXNXqlwrSNuAuCpj91l
6MpxXLTXQ82l53fPJ+1R4eYv9HSwQ3v2jPR4sU54Jki68W7219qTHOKKsKs0b01lIVqRxnhJzgPW
Jn4ui3UsE7qmj797SglXyjZfRBrwgpW5bUIog8QGn7cS70UuzHWD0OpeViRQJnXwUH2PFfMYThW4
3upNs2CXNg7YFlfA1F+GVTz3sCw4nePxBcHSFgNW0MxFaFtAb8W+ZYu2/SvJg+kPrutPprR0tuwK
HhsUjhxtmKkze0HlsbdGXe9S4+UznqGRLEumEokTkxuo+o+WmngOjSsc4N+AT9dRCKmASE8089ll
lvBBFxwVqC9mhKIPjIwctON7xMLjnGNhFitwY11LOaufTe3lrWdifa/hNzYTrhRRHlILnp0tBFkV
/oBdknL1xshtqRY29pe48YvHU9VACcXNJN7/ISDRUI+Ayb/ul+wFR8pX/yG1pSh3R2Lo0N3ZAqco
jSm2ujXvGZfMQ+6ljQxw6+nEIOkjoJyjGXolXZgSHKWxaeMA6VlK3PjcYsvNWi+SYHs1BXbTk18B
7wf+GkVjzn5d3HOVBJMDPUVyQTEo351XFZLdJbXw3IcQ/a6WOm8rb79PcjPFEgrtKl3S/aE6pyxf
o8iui/NKwH3iibUQC/6GTAVtjUPr8vGmyKkYbP8yn3X627yhtJcVVp88+SvdsXZ8bObutwG4IF7O
/37a868xEAjqwYNQgV9H6sB0yGL5sN2twFa/PmhkgsYoTE5KfAYafhfOo9iFCQfuT4nRbd1/UIzq
RvRRQI4HGD8Ve2Fz+N4Ju1hP31szWXtIbjY2i6n97BBv1EO1BOmreXPFA8+RDN9lDxFQlt2Pzk9d
juh10sL9UTBq/ytk6n7t1sx+YuktztNCeLwW3AA4GMODFxekXn3qjd6ELBGAxcK0lvY3uZwZW+UI
mgMV/8YWRXuQpXwx2165kSvl5m8td7z1aN2IJzbn9fz5hkdum7ev50TnNinB1CEGJXLwQHypp+AV
xH1E3w3+QvN80IbYlpNFoKmefH5fq79fYRR+XKyIxIMRTLSmr/NXutsP4cqAsAFhcHxzjb9YHDrv
g680zQf2KQ21xGADIB86UXvw0SxLOi9s4POhzLz0Jlz86UzcwXaTSxNhtSa9AboPVFj43jUsduuq
3GHBH2v0GqTkiqHB30YXNgkxRQDuTSBUxLP1tLe3t0LhsbkzfcIqLksCyCUkIpCi4EUzNDpIAjtT
ZIUWMPXwQMgg0yHXj5Tsl3eE7OWksWSB9IQ7g2CLiuxnmRg7r5+HIajfcg+Lt6P+U8N2E7jBZiwH
ddwKxJfEfONuiu7IM0WwsTqHPEXIFUrHeVugsBLa2yFG9Xe8gZkw0XT+F+xYU1ZqY+VpCntZeMAb
7x1A2JO7KuLF/FSXPni97pjF02p1LAyKEe4cea5onPuSMcB2lSSU3H3gl5fpbwa6Gz2F0HlDqAkn
s3vBXMBjozfYriBzAYZuB0gpbAuGFgItlbm4wXGJ6kVmLZArlxKYRuk++4t6aG/WuBD+vhHDXEIU
/U5fxN3KSpPHehJdLLnu4Y9ffna95F1r4lVehG/uJe0V6KxT186MtSI5tH2YgEVHRuXyCJ9lkpOK
HdW3utCKfi4MG9NwEwTgdih/L5J+DJdAkY6dbg6VWKNv119q1zH0wNoxuKDICcNpxLuw7EycBGkJ
Bx5KmvFs2IyV8MHthjqCn87DaMqmwpj5BooY+cumaRNPAW+VC47rRNpqCkXSt+ntW0sbHUV5IhTk
xIiofxx4QoziucXNI6rBowgQgHMoIuejSQlDeVoHN+qL1chBgnM0fdCh7il83ljZtoMpI+VnUpmm
l0mAGizaRgKb9YuzjgSHWM3SP+rztvpihOFfCAlr/R7+iLDGogM86MxLXjBIaZYyMNGFXRFqmIKK
yOpfjdW6UuKx7lOCU7XnsbC0Cs468GbcdY2uwSxdx2rYuI3AsRsLsma8vLr5Z7OCNmE5yIlRQWap
KltvdIouDBgpDQ8FvVCYBGEnbtHVxcK0rJyavLGO37mazIEcRyIfEuhuhSimTCPzFU09ICLaAgIx
fWTpQ/tjidLd2THeR+fzPi6pQ3uOR/EWv9rxK9BnJ2lWXn4sTe2eyWPCgnSaSwSaePAf4hAdkTmT
TzxSPrJY9MUai5ImpPo5SHOf9mrYTyeGxeAZ83KPyQ/tOV/8KqkHqDh8loLEmiz3PLHvhwoOnsJA
yRyLGie+89cyLHAnLjxx+L66OVh7UigCDuGx1JZK+sQ1w1Uzhc+2sQlFZXb+hSvd3Y2HeRdLSnxU
dvBYVpgYnV7lnxruGeH1phS3atx8LmacTjjCrPvo1cT/2kkPvFum92hk2wV9yEUtbI04Qc8jwZZ3
6KtUyvXLd19EtQ3PKAthWgnoFRBvnZo2prcGbYGSZKwlC0CeHaCKP2GxCbmO+io12MARUmbHqzv9
4H0H8WtGqDbd1IW9tNkCaPsTvBoa3b1Nhf46YxkW/Yp4pRUW6SRAL8nS8oFkfhkn1VrVphLwV6Lm
cGewAS//Nga/oVFNOQ1fR2PiGhRPeyvx9gHDX1/a3UObQYaPdIJPEEQARdbItGkc8RMscIrGsFH2
Fc7R1dLY1GSgTwY+gtDeCEFuOuvlS7/wvECQXDx53a+EnllC4hyC1vQonZXudGRJ6PzzYmlQBg8a
sgYg2pp8YU+7IV/iars7lGqfHY4aWxgSOe1Fo+pyurMKTCYaXvfLxuDPHte/8uuWac9PJk8ut93V
W/o8PmXLiqPHG8OWFUSDA1NYl0g3U//tIvAOLSWFXdtYIPB4hQ5HwQL3YaKLVN4MnjBRp61H6WMO
8MvDb282JF6l4aJhYNp5PdhV9eOlELlQeY0v4ZdNfx1Ks8MKwG9YBX+C7nSqF4ypZBP55kOY97t2
jWgndwfl4Hy5vySMjOlR6mQ7fSlTViCdViXxRLaHeAtB06c4bgPykYQoppr1UF9ZTooZ147GViXI
TIuNeboTA+PCZXgZfGJTwLJZf2qPB7yBaJsCMTYK0yGfJE6qaJ+TFA9kiLWn3/VIQnumrTsv4an1
5Ps7muv6VEbyJZaELAilT1lHoWGFi6DpcSW3QSLWJZ/NBEuHSfMC7OZCepJOhWvjxWVnfp6FfWn2
C+mtVhgzpDGJPXTuIaWKWn9b3g/OKAgXq+xamjkB6McSAODgOZ/x2Y0Xg5N2ElHZv5CM/eOC0XI/
k3jIznCNLGcVGgi+42NaMlYrsG6FZispOpo45EyMIRNJchiE7JhGkBp/JifW8YoKSVRoEyUQGSBl
6Wg6VANR/I5eU6lN7zGPQt5Gl+yi4sSaz/iZgnat/BreFCnPwPM/ZVzAsU3tHPQWjlBjcgGvvUqi
ecnlb3oFoqNMpDaeTPhv6leDAkKVLxudjD2O6Ei2mLSLAu1JFKJSNuroMB/9172EH23w4i4bRbiM
R6Wp2Vd+fvt4CoNjsWQIkb6X+LJrbadpQaMTsbQi+y4XMu59vZsPbdHcZdGtwSdujZ8tl4SRvFeQ
ESmBaPmfPg6ioLa5SqytaFmK2AjuzbMPjulFfPoF5ZrYUxPaWSwFN3Hggh8bAA422KOoHLBVlToL
UAFHpiYKKbxGokojWzbUix6b6TWXE8CFawu5L6Q5Hm8Y2jaSU6jGJnv5GjEdzU7gNSfoL6HuzvfE
c0xGjih1Ft63qndfD56j3fHBhHt+qIT4IPcIXaZWJzT7hswRmufHkY8DLSQr88hXrEUJsFuMJ3Lq
4/ahWXEX/+gCjn0rpMiUT1ep22Iyitkh53T3JFjCbKLeaCvccuvuf3SSxwGWwqnyLmBzAATn25s3
a0zgu5Y/o0lxDViImWH0CpXmyf3DK1KUjuyBfynjvO9c1CWXpY1qWXB2h5df/uZZT7pwKICF5not
ttPEoQssyIiVE17TXRgNwoYEFnUHFmG7c8qBG219YlSnY2+w9oooIoSdQWLQHRuV8OCGogOMVOku
WaHrwdoJVWRGQoYNv2uB/CelMf90chbGP0qdZMJ/QvLdMethpXMqfQg7gmvgratc2Oc72N474Xf5
rsh5iCGkDuehj+H1nNMD0zRhcGQ8AhoiKTaVRKRo2GNUdV51f4xpy61H5DpAlpWU7FjXDdrRTYQy
QYznwopRt3r9tUO6moB7dOSz+tiNbq03YO8g1ndElQOI8aLoFIi/U2VQNHLZgYhFv60ysm0KMbIz
DPxM2aIXimlrXo6PEYi/6TV9Rc8YGKZQU+y48DC8+ATUzj58jfEZUE+aO3X57PNvLn0rlV+0Ssel
PNhMSUHr3ckA4PvWy80KNfAer93ndyfKpoW6GU1pLiytiOeRwTJke6KK0HGNHvTW+XWO6iySmfs8
k1JrWYbkE47moi22Hn+92vi92rmLHQWGborsa5hLhIplG6YH5BybGVuo7M0Xs2L2nSFqAi6ln6ZI
ag4X7FLMC2+4+KINk7xn6x5jsNza7qvzlegAVDx/n02DLY/GV4aj129JAzvZDuJr4Ew8uROzBpUl
W39awP7HsWz9WI7B6nvlMuhbO5U2YZLriFs9tpNUhiJ4YwKDG4Q58TwOTe1d5YWK7j/G3FwnTsPs
l5xoexuQgPAGSs4qtX8Ls0hAmX2CVIEvxshEk6PSFrPO3zGpa3jeVm69kPN/s/P7CvzDG+1DPuWE
gAmSQz3/SO4LaC5PtkrsqUQt91mRVfjQQkyoAM4vnIcBVE0xTkcj/3vda8WjRJV0ppN3k8Gm5CYV
De3r8IsXO8jRRmTneA4gS9mG0W5/b8SHynCGcDDR1oBIuvYkxsVYsIy4bovQXE5Gu8ufMWKjMbP2
dghWN0i7mq/fQx/96Jdws1s3O6TUK4vyeLYd9LBC7IlTjuoDpldBJVpfxXXu4QGhDrIq51IN8yEh
q6DBch/NHHSNsZesiqNA+1T9vANnP080Q5D9YMbGfjq+W4mSf5GLshBaMhVM+p3cOVvXBk/UAAqa
UzQ+D3orzrmKgbHa39qNH7CezjGpIrMlMT0TtVo9GxEmSAZgCBal5fVHgDk1yKAiNQGU3wRNUSiv
C0zasLhyiy/+CSWZ3pmBGjD2AgKgBLIiIUBzshiv+2PTNNIMrpVTvNx+YDybfdifDjLZbgXlFLrQ
PiUDeMAVDINZHLlhB7GMIorZbI01QdBK5dGknFjBt0toi9RPP3Cp2Xkafv6qxe+w2z9xbpSEohhv
+mDNSZiNxqTEUzuV9Lk5+/G/+/njxelXO/Y8jCY/8KXo0CbX+rT4Ty9dNOLikIHmAOkcSy9HYtw3
N892+Yg7GJWIJcKSYlcweV+tfytbMe3ajfriBq3uhYHajJd0vT4jCTgIpin61YGjdhYQ8SEldDQF
cDOL22ov04+qToTCWLsqAOrlr2xQoOt3dsX6wePnx02OfIK1l2kaJjG8ZcAQo8g1PGJte/BF/ClD
WhhfKAB21pwhmp4fcXxUGoHCQ0neiAnHND3ZmkDJstlROdX407Ymq0PSx1VWORpm402XGNHH9jCZ
UyBUhNm13Hi+umbMyTSsW4aCRRuSBkU0DhCGVARstYBSuXqCmUsIh/KYj2Qcb2HgkJsCZ7L/5hHa
2EsuphX/y1uO/rB41oRTE2YIMaREoyiCJusgh06RGVodgDWJ7O14PFI2mAb6VFPv30XtjTAc1KjH
aQp6sVrz+zw0tkAulNZFfhyQwUFeN/9WgSODJ3QpseEblVdTTO4tbL6htzrnECvXjuNYGHuhu93o
WPyhlibC8SogTb/WIpuFZk5l0nrdkIenqXpXynoL761BLmy/tBtIHpYjbJ4E/Cn93FTgPQYN0qpS
AW6RT29qbTw80Iss3h2E70KJynZkMKwZ9t6zEj4XizrXcXghl/GtZDA4xvD/gF/Qv2W9HnChYETZ
qq28znzZ6WIPxWSw73MvmjN6HTMbkhkdt6yZdxrImdwWVrkeIwYMgQKo2CHqSpBsLtJZb2/XMELC
JPjUJv4h8D64I1gldCkFKy6tOUCUNd2S69+zy89ibibBzakWe399lR+9C6+IPhgM1Vv0i+lbhsi/
t/wRLC6198s4mVN8dTTO7ZSUJQi6IqiRx5Hpt4dUeCWOknsteYq0yCb59S7ma/2wTxv6B889uxdY
136ozgBmmc/yKJKnbep9RQDtFnyZjKeNoLXfrOaTUaHEVSp8YKzLbfwpoz1UCpO1fMUJkcugJp2s
abXAoogFQGrcT6IJLhm0s2X1Zetl6F7hJfQMWhhsFjmys2NTZizvctB+ZHjtDNvKjojYO2Qn3zak
UBe7DfhiNr5sz+k3aJnajg7XX7otvzlM66a7BHYdwA11kfduUmNe7alMHfduHhU0R9XDZsg99TPT
W68M3u0j3YCI0RQEhnV9vNA/+mRitwucDDqKBvvMYITmjLLCj3QNRznKpSpRqxP8T+/6Wqt9t73U
b8WSzWY2gp8/U+VnUs+5OmraMd7pGxNau7MuML+GJA/mqjCo299yyocezU7twFkhV0OzgAt3GU3Y
7rltmNTSaOykjHTq15rPz5fEHbmSw7SBE+6j1fDpk5l5nZtYnmoQOU8Vz/2+H/nm9NVzRUVI/yJv
pOf651T8RLBVUAEv1U1OiPwd4IqWmMmQB/VLGg3YOAh6Xt6lA2PiJKLmdPiOVV7MguEMdWtqUj+u
9f5tYgLX/u4kFwrPkNGE11HI+LqS27M2QwWXa/NaF6BHscsBaZtePY/Ti3y0y0aQX7m6TzQjTVJl
5XEAX/ua1KEwCaolZg1tKAf0PJ7+tLbANMLG0jAk+I54Liio523o7lvWSqXYff26aFcR033/57Lb
OPNJUDEystFv0kplSCamjN8UqYRR1s63sli/NdHzCe9p1lMQmcHWl56Igs/G0ZY3yOl22fXiLlQ7
Iw3qyDrn/cUQ+fcnhLeAN57qQ3r7uStEMcYK10crX9L0ecELFPTB5l5mWHRAVdW7n5hQBiP9pOHc
Bf6iIJULwZuOVZghOhh1BGisQp4M78skmBjTUJTrtMXifux3D1fa1XCG7QwmoSgU9k6e3geRWb8u
rhTcCY1q2oaI0sMvliOeuCmc2pm6urNFYPv9UgLTpUDavGZ0PMqgEt3qDypokdM3X9k62+R6DOpt
TI+P9WLecoXfTbeZ7vFusM2YkDcpMjHevBQO0lmqam3YUA1K2AFDEa3DVhzA3MHUIpxYThaCLsVJ
MkcZnVeAga3uBKtzgBL+PGvzmlpuwOJa7AMgeDOvfleSYKOJtmLpJ16bFlBWyRlGVqoeWapPbMh9
rs6+OEtT+CLU0DJx8q6mmLhEUBt0jYGcB3H+Tl0b/IFOzGl8/EiBXll0vPYbbDWPQ0pY/CzenAYU
nnOSLrhrXXccmlAGiYHrXw0SIjdS6nKobXwmtL1JZd6G7E1PxpYYqSna97sAb/Rhk++CyoQVeISP
MdQYG+VXkbvq7KR/OllV7xa8a2jKAQG/qK2zmMs4vGuNVCrqMnZ4ctnTY3Nhb+qSyjqC+LUo/NSp
5yykipgvDS+Et6AkVSCF6HjyYz1bOS5wO98lM9VLhClVfw0S0nGrs+8v7T/JuLS8BbzF5VzLM10n
0Kdi7n9M8VCmMlBUyp4oIJA1hmJzXm9gJ76Bf3JGc00mHYytbld0GJtc8hz7E9uINuS142GhGnRq
fTgQsOwxj+d9moissBtz87kLmfzoC8imbpBmYLvTdZYCgnTFDLQq1Hcvor2U0Bk71QFEMCNnz2V8
XnS1OLPxXqyw06kuPyTln/0iH9HAqS/BJ83T3rRPPASqC8FDWOwnmWsb4iIQAt6x8p3P+UyPUrHk
K1GXBR3pVrzWWPsG4KCb4liK2QGKqerukyDBemwKap+1VNz43w8p6rp7JMZa2QcByRwN5HLqnPQ+
dmRrqQUsgspPyiTXa7GbvJsTyZZDliG9de2f69zToNFZQcWcybqZYXOCmEnKxsIO3Kxx3LmqaBOL
tbc4gZQHRmYK5roFQkNaGGr9KrR0XkFOBbwiZroEGNJimWLymr1qnj7PqTW4ul8eSs7yxEmHkgVF
7CSlArigLVsbsoMNBMXQPrEoOORxp44X/exsNj0ZwdP8qXDr+DJGe3jG5ITTgTAjSlXIKnI++94k
t9LBxtrFp3xO1tTLNWp2FAwo0we2RkKzsKzLM3MffNhhiOI52KB8l9d265h3h2sIExKfDUkGbra5
xiANmMemCze3hLeovD4xO5eSft+yjhtbbI8ZBML8plVWx1nInn7CukH/ou37k1+rnrlQaZr5q+a8
dNZ98AOCmwUEexHLFNBIYMrdNVb0XVtufqfYkX9TxICokKmYzfNXNSUQ2iL72o5BWW4IdSjk3u6u
2ZDajFSdUKoJcauRYmgzrvBfwWLr2uUb+vXpbd6xwEDMCpOUqIACfxA717jyzJlcMq6LV4sPOS63
9j1/f8VYzjyEEuY0lRqVf0SvRTk0VbOO0B4x3xH1ZiZQY3L3jq9Vm8kcpaLZiZPf1yNEdlnRTQrg
R/pMmNZ4ZrQLn+5FDgSB4yoiw9p9tiONmxk3JfxWmEVBNwsEOKRvr1DAlJikRUqUJCTZSY8ldFxq
Tsb9eon+/eM2xURViG53nxwjmsGWTtusHzetQ3c67fh/2ab2T5TAVJK1HNuRlwsXzxUP9Z0SY7wI
vBNRtm++PtQvH9XZ7IylpeMI68ANT/PFTeYF5B9UD4mj+i7Kd8de+Flejazz8XZEg3uvhRaTe9++
1WkF1rLKuAhQi+NJib5kwSyzNI9rLXTuE4tkRO2qzq+ntCG0t4QSlkAnoBbSl0xnAVfs55GmGzoI
drKEnT6KI5yQD+pDP2tHY7IcuN8AgghWmW8HLAgKa08B9HKetH48ZIA0IdHx+ToZgXcpt47I6+HM
19IK3Mwl7dNRpFHtk2+GwrYBAfKBgEXuRZSa/UqXDYEe1Ku38yKqYCnAtEE4NoTNHhTdBLjUgHa/
0RJw+eTCUy2cGH+l+dH5DiYP8A/X89R/fS6qdgArmtHSKaWDibGPzUDqJaieV39kn8HtqGCTMI3M
Xw/oUfx3oDxsjA0P43fE5ISb4bSNCqcrd+wMoMFjwj0QY/WpVv3jLqKazHqsg2STCs8SyjcXaj3K
h+xu4WrFxitp520WHFHjzYYtdfabVMBI7qnZUGRlFQPYp+kKEwMNC2bMRuIYNHUhDa1cFM0BU7Q+
Cnzuq6/u7RJqweeHlYMzeHXOXcRKdJt7fkTlmBSt4rMqesHX+UYWpm6zDVq8NM76fyqY3BO5XZE2
khZXiMZYl0P9Nnwen0pcEyH3RWnuCskT7FWyKU83EN8aNCfxB2A/HBcX2Q+PICNMhyaZD2svfe9e
rDgE6DSkzj0VmKccV0gOdYGz+NbGTePzzd7UvvZsySlJsIZqtpHp9dY/FbvBLH8MWCXOdNt7ucGz
F99AN0YDI0gJsPYmLpSiBQoZZckx5QmCZlLJCte9aA50v3sKdF8meN5QiNDylXaZCMQ3ex3GFOAB
MiFrfFur8VC5YwttcMdd6KnxyLXYaAQ9iODCNHbO+r/7eD565qgjE0hAHfqTisOTq/fCMFeGgqU9
GlXRudf1iOF0p1oiWn1Ew2bg76RaC9/HApYK2T6j92SLz5dZ3OiV1KMTWRQ7iYveQQknGsApGKKs
4nrl02GzfUOa6NkLhiSE3M0h9lS5XQePU3KAIvJqwXzx9UhP6sgmgE/18xwO0c5Xy+lzkFKLOhPn
XHH3efveHVrR7PyqeZSn+Ft9xBodLRfuReUM/xVrOxXPmWYt8eNT9gPfeFA+e0/3YlMsdZWT5+Eg
lvPH/sfVXZAz/2FCvo58KjzQqRT7Dx4GM2/RF36Yb6OZe6BIADmmQiM5T1CKomkZLrvy+PSKV+h3
oE9ykN0rIA7+gBFQDyIJEge40lav1p3SQFVPGFcyeEM2FDlcGO5kdz2zofU9T1rL0zUog3u/oiTk
LmO3ps/HmMmqhTc29EkCr3hAUAx/H5z5WOV8awlRdJ6My9Gq8K0hZo/JMBw6GYWI5WA6SoErUlb7
h+Qq2aTNrU1GLEbaWqh2UBkh7sJJchOQo5rYElQZ5aTjx136rBqDN38yBpLOvaM1HgM/cDUZwoKK
OH2cfb94eaoocsg+fL2CjxlRwuLhvcQwbp8DzwZX/6k7P4NXFmBvsdFmtf7Bk/8FoQf6NJ1sKt1o
3zugWW61NPO3wxPW86KCaDCEPUbVwKoEIQ/8t+qSu66xAhKgp5vMq5xdZTE2Ts/PbHeXQwEw/ifJ
IR2asSbrXLmVPhwLRi4nk4gK1khqYpnwasyZ4SH17NIxF7s85Z+oGgaThlFtI//8E8aoo2goO8DC
g1rhIF1yK7JsGVG1em1cFVFWbl2BlQfeocoE92BkpviQ7fBazdbnaSqtr0eCwIatiu2biVK6X5zF
Cqj7nQPkCystdZrLFI5UeGv0mGh7Lbk8MqVCaTDxAHMOZUTPN/BlxqMh6eUCjiAAASWrkWAmVsmR
6CPj95dmOkurTdN23zIb+hSYwsgnTE8GckhreYFob58/xDQ3tLIwVe1x8Bf63zWDVmlTrU2L5tYE
at/qe05dYZCEwK+NYt3NMpbiL602MYSt2eQT6arki4VohITAiGCnS3i3kJhImhnfRifpye4ZPMiq
6JWXxM9gxJR9IiH5I3LV/KDNYRtdDL9cYN9IwsxNwMEGFlx8oaJ3moSf+/z4A0fBwp+SGFoIpcvQ
Pv4JMLFZFB6VMhGOD5YjUmI+MFwFqbCkVbnbvkMRMxfxLAcvvy6UiZC7yh/xSb3mvQfhsrxExS8z
OP2aKP5UgsAMyjDvV22hRJQ3BAHkp0gIEKYdKkbXuTVkBzjhJHmC5Bplak1A4UFL9WaktbkXvdAD
ni8pwb0jB9XsqUl7D0X6pm8vE4ixolaQccNY0aoK3X1kD+VQmp1yFjmLPyyVc8Inr5Zsw+ytUgNz
61swt3CULhwrtcavMi7ovrX1/nEzob8FgO3yGvvj3jwyQhuqWZXYKL83J1VVWcoZZjPFWK0s4VTn
9ummPKhBPbjjQ9V91Nr2W/WarKmASNr81lIbS+/T2XbNgY/i9BXaEJpWJarsz28Yt9h1lFZ9j9AC
dysKdyw40/el8tvh0Dq98ekFovNjlozHwpKr2zJRbzFPu2G81vi0t4O4POwO4Rkk9ZYLrE0dIt1h
2xgfIPsX7fSC/6J5hINZqHWEDxD/v+KZB1LxW9x6VJSp7OkRe1pAguUZuFBTI37TxEhrRd36hBXw
HUa+H+IN20I51i2vXC5I2UR8iMA4El6pl1nzRNXcch26AXRbNzDHK6+WrkMDvM5rURmbcHEd/Cif
kS7IkB1ns83Qhmz08EYwpG94Y7HYJSb05VcFf2O/xrYWsDOYFDE6j86HvRwK7wjqgUr4cKlTpMht
3+g38tv7PnCwfaxmh3UpWq0VN5DVGLs2CxU0TeWfg9uje5mlrN+TZ8nOfusLPaU0fVQpuvXORQkc
uylIs7lhao6ddxwLxGssYGxCFEdp0CmMZCWfsGM2wY1nIIHqFi+jUagMacNKzw9ilCdrzP+ZEk5C
yQlrVH2lr0phUpkrp5CxLcxJuHTdH2ZTUuJEFRDwKOh27//yXB5bNpU5iVPEROkRcKjIqFx9ZBnI
O1UlSwQbPdkzCN2CN5xTST9pWMIl4B33jxyUlDGTFGNp9AFIkcQHaIKXunmUtQZbmG025Twlzgk3
4MgBZmC/3loHtAAReIhyaCBqD2CyComPca5Bt6i6y2YS485izxCuMpE1YEf3REpbGxlkrSLrpT1p
KPe1OuLrt6j1KV71wSpZ23DJjVkkSeRMr4PHmh0sRLHtXvhaG3fUjNFEUzTUzQupGTJUm+S5kZ1i
hzYHtP72V0iIijJ5/ac/yUN9jmx8vpLCByfv1lIIZ5OziR2ESXWpzrnWS49CDy9YvH/HXQl434If
n6YCk8ZaC2Fpj3ouG0EKdzSMaaFxThY0I+MrTnYJS15+LJ8v1Aoi3eEqogzFiqrduCUrQKjoLbTk
FT2fTAsouCO/mHDNnjbXN9Oaomg1N/0jMT82fT5I5JsT4g/VTyoIe399BygrXEJcdPKQMnE9FKw1
+Dem4GTWscJV5ESZlWteAEkSOFB3rIrVqrgAooIzV4sTbx1h0XOKpdswJu0Jj5YgXcYsijFpHT4S
B47aEHyxUkR9p7K6eL3I6Hpl7FbdIKgE1N7gDOfJJTpWNf+hYl+3RbnESeqNqJ0uDlihItZefhVV
DgvUZVhC6QU6hN0uDNYgSRrep0SGLhoGsm4BPcGcpaWnxPFOUp6KkFLGI7wJ89Y7QG5WwILc1T4G
fZ0x7TziOPu9FS1RfywCPvRex0twLkCQfGjXVc3QUev8h3gz3H+SWwd6yJ8mf47cpYyYVdbKk40d
WT4pXz3aSiDMQlBNnQfIIMpsIExUloV01LCxOFS3878mit+cygJbeEvWVkslV1ZL0FjmEIqvcujm
EssoAfddhcvPlGXXF1R/zfUGGApCKKy3GHTGl6t1cZRx+IynISYkZRsf9WbYwGio6O/h+z+3fsHQ
vJP0SYomNaA3cgTZd5iCfYDwIBp9hCkDNmcs9PiFTPoQmdDvZkKo4T/9kWC2q3Q0OMHqTn65/z7o
FFR+CnfM6Cxu75ReLwj58wYWd4OftfJYE9lwFmjt/KCVYUht+kiB56b2ksGtpTlK5bG4CLlVITUD
D7PcI3C3qWjgjpWKzxUp8LI3vIARqGfIFXGD60iSfTjocVFWNp3jpfGFcIR72vEjwEA9IX92aS+9
tzP8plhVZc1z1mRWBJu8dv74r5FbordtxIj5qfUVYhOPCQFbvhM1A53gPxOLsP019blh6xDr/qUo
AB7ENCfifBnLBu9A2ucK6cXTYjvNgO2Iftt5gSBu5W9NyQADhSQGx6g/Y++DLQiHLDsrzg6DP2qz
wXuo1IQjnfbVfY1OJDmCKCZRxztC7Ta/II0vMH0PmO5WjEOSEuYSxprZqe5t50GSOPZ20VQrDX7u
gMBFeg959W7ImtagRbsq8ynrp93pZAEJyeYyzaGUuNS3dcrEmut/0RZrHFWEYi1RmDYvE0y2jcCw
SCwQCRlxf0OYda4oYQcP2rDmzVOYgt2G7uAJVnFZZPmpTjx7QtFGJvlBROOwAtY4VKRiUqxETgvA
foJX6v2gTptD32v8glHn0h9RCDkhPLVMUEIBd/Y8X0oArSXqsqu8bRfxep9gXSyyir7rmRhn87eK
aBuQceukKW55VLAvBIsEbzu5LsXe7rzedFUnvH4E2P0BOnwN4SMfyY7+zeOsEIu3VmfsVSgDKmoc
566PMlRQtcTb7gm4egT4/j12fShZshkAzc7QkRPSWBm1lFL2Y0JzkVRFFuFQ836AlT2fdXerA42/
Q4DSSCzyQpH3QiQiyPy7eyQUE/iC06wQizWNMR/gngXV2jOoX00T9xKkm7+pLQ7QnY2NL65DY7nJ
mVXoqPflYPPFsLGVO65bq0R3yy6KCzW5Ql2fgFK9IpJeXuBS3BMnJ4ZO3fdSYQVIZ+hAkxQKn4Q5
lDNklq69byKn3ygmrLZBYaz6PrPDg0KkNulnodZUkbiPmUSx4U+/X1LYFGNx43lwS5exp0EnBCsU
xt2hURDheXMH2meGaRkNJA9R6fwbXwnFL80LY7Cy+7yh9lqsQ0tFCrknMrPeAyagtkkMRDN2/+r/
lJb+qsKhEPtcZLASXztqOFBR1bcdiP+PIOEIU1PgEDfIizJW2NzOaS1qCzeEtQbQjVTp6ADBjUFs
gUIcNz14mBI2psGE67s9M7H0ndbgsNb66VkdEOK+dURKAetkQdNTIln6aT9eWSPe0Pf1d/YLpEgK
hveHgLVLWZpO0auJnziBdFtJEdw4Ndv74slVzDmJaRk6UUHZAnC0bkXffX85WkAeV780XNDMSk0F
EXCjQcwATvYUbQHvJCY7W7BanB+SZtFvqL9YPhpSuDRk5R0MaqqCljotXWnhPHw3N3eQH1XzCsr9
6/dOMRmwe2rYBGO5svUlPaZHrtqsSK/iB9DYQCaTJuOViiSB5o69d13O3moGv0FJosFJ6Mx9KM8j
lgydTxeMTJrSoilFfLsE6Qg08DULxSmjuCZhIHSgWk3zYyEqBUG4dBaong7OGS1yV9g3wa4B1b+g
q5vKgLjLmCbRc6ynWZRD4AEtUDDte186Al0X+hEQP9GRf0h0tvlkfAmWSlSS3JuIP6XarpRXj5E9
NNobgDAy1KoNGkj8ax6/PxeLno1ux2Il8q2uQlyaHFzfc9i6uwfDXlYdMvdrON1yBhHMNwFhd2bH
Kwnfi/IQHZhFZrlRCupaFCty9QtRZFnbQdoacfSXDaN1WBHfhrmzss0g+HEZXZy3F+5FCkgKdVyg
e3gnpIJy+q/EpbEyyqNnLODlb1/AqbbCKYspRHFCBcB4BNSt3z59X0vIF3NDMtFJpuU5qg0U3X0Q
28sVLbJOBulBuNrcGb6+E7bfG2dKeSKZzjGPriA8WlP3aihAsPMr0F2Ev4QyG3CEe4KbG66ykTOZ
fj6+ksuimmzjDYHtOBjGnMY/6rX2tB/iSwjow898xasICRXkWIuP/vq/5id6G4UTCqMyO5qsKV89
gTvnjYc6BqG0wm8zSs2zKpNhZcAkW+vuGMPo2Nyya+yseYO3CIswpMgbxcFqq6lQraCqvEa6zq8W
IgMWvzKm43aEPnOUa3fmusJIhvKIRDhoKDHWL9350J4V3YG1LDGbvnbEGNHciEZypRyBBg6rg9zt
QAZTDAdKDtIWjFUAd0tl0psfHwoGpuY8INlnKluVqXyRzlbdbL79hV4zA36DpsxRWwh42tA6qyY6
hI2ohcx9FidS9gk1J6YHo1/6PzsivXcISN7eyQtrZJPWB+ikBuVPh1NgOkJSJT/hdc2G1ZN9FuU8
6lUOOMZR0gKkNTYgM2yDFvn7oYHbeCKKc+OHbSyJgaK/Z5Oo5N5weHMMSf6kaorBZS1APuRDHa7C
+H6e08DcmgKIAxM5Upz8L+MMGk2fTPScGMexYPmB8Ja0+5tQnH/+A7BoqU+hU2H7asstbQaV6QIv
L+qk+SI0rz+wbN5oPlfQtgQTNXmcpjT2WCisVMAuKH96Awf9WWaocVpPixKOcJGYsE2Zo2FSCNY8
urS2iCWHtA3dxLL7erdMQ/g5Q9/7PnySgGRSo7W+KGjzQDz0eGcQHGiLK89N4YNslgrGrLl95C4n
Bo4faLHtdcxtuea1o1dpSEqUXrjibz/VtxtAeuk2Ejh533isRpNBKT2hHeKKtzzNl74feFB/9A5p
sJYH7VtSGDYOw9eHJ3sBFUZOyBMxgmBtyTUHOlDDTedY1puc6uJkDzFC9Mj95iPJwO9Yh2ZsPSeD
PbYd43fJ4aJ29bBktkmwjnzqnGpuqlYoNjZfixU7rLl2tBf/DI5x+IBdRjP1YOGucetGf/g7ZtNn
vBG47rptV0F3bQNidbPdqcumDxTT/hr0H1IQSkTLFbrpW+g+Aj8otQTXPxdjXMy/niAKQMd7P//J
OtDtZM2KvCSktj488jrRcBErRwTrcpBw8MR39aGPLPruKegooA3SqeCZITS3MrsaMCeHTnBJauXb
xqX7JFP8MJOd3HBPwrb0DWedM8tfFw3c7zfiZ7cOO214CSLi4aUv0cNCn3LwJQ0PB4kg47+qI2V3
qvatC35tWlGTETAS5xf3GPOucxgxhEld9uieHVIHEI+TXgiNjYw9Bn2IUkLyWhDdsbMExmbZm2s5
/35d85h/M3Miyp6+NhJ9XOeBWkD6/KYeUgRpAguY5eQvPwvU/d7k80x51Lm2FwD/2Qb+FEvvg53j
LcbZhYWJniU/rIvrwiK1GHleyHC5c5sDtDkmCiJjtrEUCrHdNa3fYBbWLRKkAWpOg73CkGpucGUN
WEH6n2OdpKKhWJLKcuWPZM/lXOSKdFvB2paOZKE5eT1rcu4wCMSi1m81ZMcMB0/2tPrxMAB6IIcG
KzE1ZqbP1KqIZTLB/SjfyS0ulINCb6Pmdc1bbH7D6A6sJYX6psCH/3CDbG+ZTEWgYjaqPz+jMwee
txAjD98nlMdo4lFVr6aRFDIe+zghemooZBP/IFqU0PmP02Ldcu1pG7dfmy+gc+ZfgzWcKphmrD6H
zxO3YZHzWEAhIXrm9EeqdhPCYWdqWBQbzNaAY5HCD7jPpiMNfN560KvhwauhHLbDOUgKqfsx5paB
YAP+fykOR0Vtqaw3XS7WuXgbQoXnLI6PD/7wdp5/cp2T2T3mvG1gfpEpwQ+cPP0glfDFsfJ6KYSu
i+AXmEkJyKONlEhwLzWmu//AWD5o9w3AYpS3l8kXJg7oibnIChUlzKK4XtUSP5x/tmDrmuhs9E6e
aLSE1c1EgpUDJOo0NBlFTbktqmisKBAPinLrjct8x/YtP9GUgM1npz/zh1YH4fuHivkCc5KZ7A/b
kgy/rswrcEcf9SXYFsJgCHzLdKTPYJxARgJ0sAwhOQ1LM5SZGhXiHMnchoerXdepL/u1XskoVhlC
Cuil09QN42afw1stNtQRPYgInM8IY8N8C36ENxtMeG0O44+ZrRkDAcd2iYEuD9RmQYj3gCIja9jq
GYPEIVWs8xDO/hjL++3LeqgrYVyEQbptyqHwiYCnaPe0DohA98kaEzewTSr9OnC/RXRtC+RjtbM/
aJzgsyH7gXL4Bnb6/PcYq0EP4oPclgiKHhhUlFQ+qzWGBkNaXps/O5OaRgJwGgjiY9n0ToHtFvQS
AEgJ3H3yxNb5QWFlS8JYMDhPgcFOZYqKLEAPimTa4TyG1CAgjHrlPipl15pbQ6qIiPmMojcExeyH
hSl/0AC3jxB5dwaHmk4YLCPeSeCs1Ja996Zl45SzODoCodcZfIr3IEDPJuFlm1jhMdtlpR0tor5z
a/tolXvPOKOBZOb0ZDaw0CAC3dwOnvPUPTtq2ls4zPB7+VVg93fv9jYIxz28EOp4ddVuKlnsJKCU
+cLu49ZinV6rBWvpPlh17oJpbkW9HtWt3FxB+LFu8/0/dup1+D/6P42sZ0Xjuf1pKHivAHHoLv1m
gJGrTQ8XI13lkRnTaen675gH9yktX7A3SPAhop8osWJvqY3nPrC1BO7OKTA+0s7wkmCUMZOB5vtX
B1cF5MfmuDZsTaeNgWU+JLUBKw/uZtryvsNQgaf4fcktEue7tvdcNF2Fdu7B33nt8Vdgb6d7fhtG
suQT6A72cz8QYdTT0EY5HZldoFzzAhmL5YuCcvwbK+5yuUoR64AuTf2hkhS5YKHJBnw7oszmUOX5
xpvNDEMK+Or05tBE+SODJTzuHymi2+aP0T8KtYTNBhccfk61fqW3phBXOj6aK3gAvxbK8uOCNAc7
bBGTgloUbH2KB/7eT3oogmj1QkUGR7cJmpeyVCBNaF4G1fmPieuVpRUY+Nw7l6wS8eXFoQIrf1qr
3GKbN3DL4oqQQnTraWBoOWlHvfl9/fDZaVnoM/lfO0B0N+UoM791vZJD23xa3+efWiZ6H6LpdkaY
X+g3EuLbZht0WKPI0CTXrTVMgV2zZxfkyRpWYTfSSSfzY2PzaZpWSU6c9yWuifkhadytx6nYbfJ6
SeuCd5Hl+f9QQEZUPZqPzQ+qkEfQeM6J834kJnbWUEcdoVKt32L6Ux0PMMO7f4DayQSMB2Bjujed
yU4dt1ZePomtj1UJYfUW2Pp9ihDTEfxFNCdJSwZ4kS/sdbmhc+/YmA6zGqLNGhh5BoTLhE+KIlTm
8iSa/uPfQ/O7hViBdOl0R0hJzY6Nz6SQci28gR6xQu7xB6xrIZgEDap5Cj0EgvUyk6X7INY1l+j3
qpoZFoyoP0WKMJhmNMCk1NOoRcA36klQdeXwrazXVnkehj0oqqHOmdC7G2qtHLB9JVpomXzYMsVW
WhtcWwq9Gu3lWoCHe/VlGQVNqc/ACG0tW0wD4LWnopOoVaOKqW98mlFwOM6LitOzwidhtqu3eU5j
TaNA9bIHR4exAfRXW08ZoSmwyyHLxVu0Pa8j9oqQPMCzkgNAxK4UJiXNTcLgSjO1MBAmPFWpc1Bg
3StJIzzXhwqblb2AGsMaaGPEFyuNS++I9Iv+v3YrD0JmysZ56fcBxjE3FunjnxziKp70Q9ynaJLQ
32OvA7Aw6gm5OLG88AQWe4lfjk7Px/T9QNrqc3LbcdRyels2E95cJwEHMvbhfTLQXaC85DAaZC8G
Gi5elnuiV0BNi2Pj/xJtMLUc4OtuhruZesw46ame7dixLzZ5pUKdCSUe1F95eYNpVUAN0i3LdTOL
GYe0uVXOroqPVEHDMHofd/DpwS27sBo0+l/KxxPCz96neLN8gM4Vt60mxBHGN4LjKoZb1Mm71N5t
J5Y5PsJvx1La2lKHCF7Jl4TEN9keWfOp4sOJdgDCyGCSpRd8/1jggp1c4lrY1kxcJRoIF40byy51
DYjfNvoYsfDyKQ1U4zx4Vnz2lwwuPbRc0S/swJ/0YxXtv78yMa7enikKeVPgsbcJZz7iu9Q2f4F6
9Erd2cDa3+Hs4AfZEKYh1zpN5ezCmIkU+K3UqyVi0mkKExBOSYR8iaL2VZP5wuRaKbvRTtb6YaSy
DzHb3DmXY0EfCrp2ZSic0eMIG0hYpFo86mgX2ZL8fZ9L4Hs0AGKC9A/pfIPB4uTsX0xbkDuO5Wg6
cOfnbnZPEQZYzvIFK6ayhr4jqwpg6y0U6cIzzBezdR9wnbiBNWgp3Qs8WtomhDdjGnTbp+RU0Twq
EQjq8PfWagKg+U5nkWB3XtXxtmqHDml6C5w3aeSB+KC703cR8lFq/sbxT1M2yqED2RA5KW5+l8Xm
zonA0zV8AUQ9UWDoPFgxSBE0jOoQBBaGVh1avco/InY+LsHrtrOy3Dpmbqe/yL9szMcZqgsBFxjm
MhpJfPiBwE8NrW0PXH93N7iUaF1bn0IlAMOpHMWWEAudIEg0a3t3wLMwcryeQbVJ/F4ug3VW4mo8
tLYCU7ibrUTu+p7ygXtSpXJTc2nsxeTSZU3XabjJCS080+G4fn8pvKCSfzlFLmwNLEPYXuyWCPOm
Rk1/2h9GCeVDRDEiEH5bLPxlT3NdyiZcut+Zx/OyPzz0gQ0zoIT/ahkZyZE3JVfMkdM9GXRdpATC
EY/6Q82D6fYXQAM6cqCSHrKz9bh+PHJzFGFBrimCM6aTfLP912kK49fyBi6ayQGGCyOvtpyslkUe
RL4R12AJi07PO3VDCJkMXF1JXqphUY610Ato4ALrZI3WDdXoZ5HIDCr7/LZt7TK9pw/ZMVeq6Vev
DWobw4LocGeSzj5r8Z68QJ1yofx7CQpgxNu9CQjfu6w24qhiNjGoNoenY0Tq2loe/5+Mu+8ckJpj
NmX9NpvCxKMmS9wtSk4zFnU5dhZmMZbFhLOsTbGmoA3fTHSYBcG3c1RF5QZY7qQR5wa69VbaH7mp
vwx0+frbD5tGqE//uuMWiDQ3nDcHRkvSnUh1uqCIr0rLnOaE6q/omrFNF2eBRdmWz7+XsvHRwRuP
0t4eYZIQy/8qmSL+J64tlZhqMlzlZuSvhNlRJ/q1nUt3w8tote3Y9MLhlKZbG0YoM0lJ47ZmdSL4
dj1O1mUNL0FP54dhBtSNJSrI4XIIEl0bStwcBWV9DhhoPivMan9XNsLcOEmw6VPcM5+vzNuGYrgn
KIgcdYO0YNhM2931c3PxePiuxRauuShaf1KLMJjHP9By/mYhl70C4ypCyU+aC+GX5OrfG2HMFGXd
IvGd6UsTS9P36xZx8KiY9u29O2PHUpBJrA/sddZ1GIHKo35b9/QE0m9tvkt0Hq5dyyasTLIsxbuA
4+w7cAv0KQIlNUwwID1sMcddHJ9Xac1CMcZyKzMhSsNUAmesS044khEtp8KDPzktkMSWW7KOHrJL
kLAHe9vAj79ISUDIroPEvfbIygI32i/fyrzzJMlq9jMmZ1g0Ic2uDuOEsK55W57E2WU4tnInC+Q4
gJIFk/q9Uf9MyqEcH64fwT2oyqaNpGMeUbihKSz6jRhLkyWM1jMUh+/wwDMUNvokLhwhLIuJtFO6
D7A7h1j/EmeQcAwhXA8CcLHAn24SQGrVjZZgx7+pTLJW3rffjLi797daPbZZ3PtjA/pYCfOQfKZR
u1CQS2Q9c9t6cTs/3FqIoakq4ENCPGE+t0yYyOi8F1jy6SH26LDegPFXEVM8lhkxj+enrktZDnjz
Ft+TQ0mckzjB0bYuFuRJMaQ8ug/Bs5x0809EZSeve3jzq1rVo/4HVGUsFgnHBue/8SSZY5G7At/3
99ZDPuA4uWWJ1H81uTzIrrWhskgNLonZJ+uhI9xjN6YdkmaHPsWLauewzWTeKdeNXJPfmrP/fVLr
6d6AfeTXW2JNK9W5iedWYvaq0OpuQyNSoSZJk0uGaaRI9zxnnEtB52pN6kYhUkWVRWI2GerUu4oi
ftbWwTq6gYc07GkK43Ung4vcD6wvghGXm3hA3Z+xQVbmPCmGKa47s4DWNI4Bldo5WpAnOVZgH6TE
eYCsjxdF9kNnhdC41/qWmaQ+Lstow7ygQ+HRevjPvwL00Y4d38V+SFMjoORtmfKqOhh8d+Z6oXL2
Pj4w2/2hYDnCTLq0uVTnOAy6zojWmEL6wNiRIr5eA4J8BhmnhmxgSCCULFH00Dyxs+pKPXpqpVmW
P9s5lcCFZ6fxi1MyKGEFDYZjWvPuGLjDHVZMvrk5vdN6HMbZAsPPkGgCmIJYwRoKLqG8CQrinq62
m0bfmIJVMq9ppIM22kKjXA+GDYHmJ83/uAD+R53ISkT+cwarGa6VHe7Ho90GojfjO4Coh0Set4k3
fnMzTvUgmumjGLRN3gzJjnYDqFUQWY+Twg8Fj+Fv4Gn/EI1gtIZRtfUaCS2LvQEUru8XpNV3vkwC
BJ9+20ACrADkxwoxOqtc0BAiKbHSgJzFfUx4Jc9CYPzb8CnWTjiUDcMAj1GE5FI8GMY0E3PHvggb
aZC7qrDuealOSpJYxsp/5ztWAPAoYymhDFDuMZ36TVu9tN1/gkBluPOv+p+LB0OIjD819/4mluxf
RJnvX3T22QgZSuljsSZpZuyOEVTAetQy27Z36XTK1J1O3dPK9M/rdcJvV+SMY8i+7qez04YhA3xm
DKVSxKrYulctNIMy54uodp44II+ab4197bC5TEbypJF06eeV4vxK547FkUOJQAfUSjYjTYMTpDbJ
KqnHpni1A1b+wfhm2+DKEoo0GL3AgkwN0vNpdT+JLXRhygKl4HH3fv3fAwDXhDgwEBbKuAy8HmRX
rLSW/ToQRR/BVnnE8+jpXcivrt2BSPy/rXXvDtK0ayjLRTguwnFrLZHZoyEfK+izXCQjKyWIKPqO
u5ROpdX3SbKdIO6N5FeE211YXohmHXP8yGEsgCrE0zBVbygzfTjQaPiO7/S29rTIM5ValAGZJsyH
Ft8m7Tr8obkieuh7GqeIvh5Z1pM9ubj2joauKeEwIy3DJC8JBx1NkIjoZkKtRoXODgbfUqdBWhQq
ZIAJ7pepICItneydDpJ0gtXWdYDovQH2MEk2UddMiEoBBG6h4/NB6tyKoIKyycOJkJ1N3Of1u2T9
e6Pk7H11/F5YHqjaR+ppJK2LEoAbUohiw7cJqomJqLRsoMg2+OySVkKDJh72f++L0hAcNj3VcZaz
YrNHkyLc0X7DGZ3GlJyp0SHwEjEZ+4IHuXYb5OuEPqpldgH4lKwCEUPFh6zn+b78YD/0WIfIK4gG
0qLijPHlmVUnicvpNfcbb9y9yOIswGiguAO+VoraWxCteWjD/5vlYg93wJIcbYX2yagrriOUXwZ/
YEptgU4/HJw4uLkvWVQlBWdFeC8bvMwX/IBkEvTMuaKmRRVH1X5z1CK7WEiq2lYdvhnlK1NEfGAW
XsXQsqGhhqz/QEHc/+5MDNUMZ9nn2Qm+fv9NQlVOrd4K49stT+CExSpojk1Yrk+k/MPVdjD750L2
nOKeDBYCH3noiolxYFw6V096jloK0ZZs0Na+1BE+7aeHyZj8pM+klXsWcKjeWWe57U4sVx5h/lxA
wHBD1KYROTKL5GOeoudNSE1+PfcFPI94qbK1J5+rzMH71fjPrbF3xWp31NaDYZ1BGv2GA4xqekaJ
GVjUrg71FuCZfxl8i0FrFSht79sVN1lnE7poRkfIsBuqIPWx6IowFAo9DQ+Hyx8c6mD/EijOnwYz
g4TXnNXRBihKfnJELm9n5n6ifN6ukqRPoJn0cGhUJGF+AwSzWVcRJpxjVwPM+Rmib/WQx5IonJbx
PD+ONH23I7kxLaocOHeFHUZGCpx9oOrWbDCwfoxDkYJBMsaYZkXVjURZ4XZwXSYl4nN9B89WuNIz
rOAH65nFh/GYdz+UveOzenMMVw5QKHMRyXGg2efawwroK/KgkN5sPoa86ijH8ZLamXdYy+S3pD+V
TLlHycKCsphJlmMkKriLQXCBpQicOTyYyCKa75ep2aqx/aRvyNXrg1jdYNIBk4QqCc20ftYZqb06
mj0ssBcjbHljdZZ9E0D/1T4CyRLTgDEKfpuyF8QQBgI8fjm4lFc898iSSdOWsaYWDwDNgZacOcLR
7c9pzFEOlPtjpUdL98L2qpyCsoM1jq6N1XdsEp7Spvczs13wqQbBZpVPVLIfY9LSoKWItT5PvWGG
A/zNyG8gzyaQ8Zk9dhjA84SDb0ThPhpS8LNyS6mofXvL01Y4d7gMBjRrkg7sotrEqoeZZHJYoWhs
9lD0yRNqH0KzSnUue+hAZrWKB+BVd/lQ87vvlqAtd7EhK3JinVLsOhN/fHj28h7/NlEhhUOthl9g
tYIkYH1B94okge6fkhJ1VKSjGdsnxOxG+tQHScAgqomhYLBOD4JPth+nzK0MRPCUGQWQhoiZLc4j
1YihPHYJ4s6cSn97aRiEGugLlN0AerOtbwFIjCy1zOEc5470YjUNJnj0Lq7kONnp/RLuQ5PJr1rX
gjxZwQ/+YoIIboc9ZX22oeQ8Z87P/Hx+6QtiEtPz0MKXsGWGbQtRTzXll8qzFGBmvrWsHkmRspBx
IPwp2gwAY8VxiWjPc4fP0bQXIZ6ZnhyUTc0CuMF6dlC/fXh1XK95RXL6e3ow0iMQ1DQ5hNez5jJ5
tlClC4wOmPMPCNgWanPv7Dd1B6FL/yMmHkYr7MPbxnyAxfjsuSHJH6XJ3724dOJ9ORVgaxfHt/uW
S2fPaojkITtTcfWcyjFvNW1zY4tFUrIRiCIUEc5uoYrANp0cEPkKdpdAqFkBOZ6fgBEVwdLUqDaK
XER9VNFDhZGnUz1d8ijPvBFa6k137DYh4S5ohHdd4oDjUFiB7T7TCreNbTc1GLeg7Pw7xDZXGvfh
a5lcSpC0MOZ2+qrxFuUTvtCKGLxWPu8G8eqXEIGemVii4RS9BPj+d41Vu9lq/SMRKHEJEg5mrCdd
JWSbtadGoYTocZsbokGWAlTaFCpqkNy0o6DkCpuFWeM1ZNhZh+uX3cJ+iWG1iCz6SV7s0SAIY3dr
DYJQdCAGolX6numCS9yVK1p92lnW03w4OZa6m6DO4q7Y+knih9TuUG1f20dOn8LZyDAAorPyjLLF
t3kjliS22CJ7jWqMMH0/rJWC7sVoncJvuzIwDJtxfzISp649KQ0cih2PddxmtszUZiOj6Pwc+Wtl
to6Z1zhlS/U7Cu7Y0P7wvpZDPk4Bb53DMkmCSA7lxQMjGkEyunOlmGnCvaleBmzZumjA/5TSaZcJ
fKbfcZnue+pLhtlfZ4bvbv/510lQedLUtoI/DurYNDOsKq0RM2fJVdv2dbkRQITibjiAkYknM+iS
hhg7Uv9GUP9VlJnE0UdB845xSSaYJ0NSlQr+jFayvInu7RlsZCKuT9fW4U5NcxVQlI4YNaCkPeEC
M+Hd+7aj8NTXia3VNCCzeMnokAmz8eqR29E6LhSKnAFks4RIkV91yvv4V6VoYr7pXFqpEkhBdDiw
oWYV1GB9Ee94l74uIF2fK0/2WagEag4zUbditSYtO7U5oc4xinDaOBa2i/71VGS8hsB30rCkrBcC
PTK8+msgpkNthL2pkkxWeLmcGVTQ9H5IVpISiJvT+iQjc+fGB8obnpTIQdZufxacwTMMiRvPN9l4
LFcoL2P47dXmpNFHlXQFWDOlP8FypOwb7JE0YRRAR50lQdIQ00wlFkBcEQB4Ljdcva6sRuTlPMo0
IucZze1c6mWOGWZIqGXcYi92b55m77yU+75jOintJLAGHUkt+XLvT52Fordd6T05kPA8cnzJ4eu0
yoIsGK2TJ3zJ5ePF7y+9j4FrW7ZEUniWDGt5dlrXCLsJJqei5sZvlKq3d2fu7Vv+aCRNrHOeAjtr
bXpO80gfaB+di8zK7/8HXPX/tZouELX7A+hCMYZyaMFR2itqkJ2E31BDot2t1IwQQcuOMK9frvaU
zt0yvYrKfaKJdA1ImG6926XpK2r80ZzdLTW0S05OY36hPldu6YnxoAbiAEz5U20zaivMaQWpHzwU
jFsOLfVlh9TiGaTX0o9cVJVu7Jqee2UVDxgvHPlcCZ+f8mWFmF0VJ8GDx2N/tVFB9vUXHDZUkqMK
Sdr8iD5f5i0Ol/1GmLCgEBy6AVpWlBZHiuFR/mJdoBXQI5XEoH4xynWbAaC+/rhv+ETbSRGNWvaC
/z+nTQvT6mST0rF5jXj8YhRRa3bzDURMpjrMtB1k87RQvOj6WJfGuYLQ/vP0FmP45e9b5CoWEJC2
LglD7wWSmUsCTBaBpFspjVjwSeR0+C9Rjsmrl1LQmULOMb99hsVabsVszo7hJYwxdKgHTT8Ch7nX
SPPSh1upSxpXAtK0pHZaWmTsN2hRKPk1J0LbMozciPAzlDFH5z+uw8IcsJUJg2EezmZFy7fPLwOF
ZfskyG5EPGv1fCBaX+ijoYPpU44/pS0QfPmQxnp3HQeX5j/LQ7xR7FhQJ0Bb5c16uzd/dtwBqPj/
tnAjK0YF+g79LRB9+pazUrdmDRufxhAGXcZjIQyG6CoIz/IupcgGcKlElRdkp7B7Srl0E/x9kJjt
d7M7KdaqaM8ZUVagUxJYQy1bkLbNh2YDU5QWCmWjlF3ENpVDXiQTXsd2tchZFigSjldtq8h54WoZ
f6y+/uzMG5LXbPpiyuWRj1+30fk+9iFYLQB9WkIVpzb4kN0/rM6SwvjASDA3mA+SjxlXYonxV7VU
CZTJLXsSmKh9gitrkDCBAnkJ/bTSoebsPpgirgvnFRIKwOLSjj0Q5wKoD4K+sQUvoyb9lJbnufqk
YAszTZW0k8qo6ui5KVcQ/0VzV6T+LY1qUf5qNgueMJS8T7zCSah6jtsgZuFrbJPR5SM7EQW4dEM6
B+nVf+g0pUa0yp4MQsRT4IOGCrn5NWZv8dlFUs2SDL4mmYHn7KNfSMaApLNl0HNsfn1uR4nfGEfa
W1BFs7qU5fvJhWLp4G/UoGbrRBXEvEO/e2rSfZQszy/x5o7bD7Qg4cFsuTny1qeWysmLlFeLq5CZ
VBFnxzCQxRYqvmpt3XCO3fzrnGIpVdVDVlP7GgM7Mk9Y/7oxECBztXgf+0CpzRlQU6anZS0jYoNo
vSwi2RBowL7bjzjTv8AqY01WskjdZIrWUVyQ63Z11UfpYBMw+oYwsLI0P14hG5m0SZiLdbIYAv1L
35xEq0yzeR23H03xhxl8RhrvK29rHj/qsHPVJgBYSKtQdpc3aRnegoIZJRZmepmVPeFuuZs9xlpo
3r0dxBXw7oJESuMIlHa81r5M7gQvuWqorG0qeb3s7b1xW2EGV6Qee7lsjeBnLWng41fd+/ahcxct
Uh14PKCzPKgCTnab52BcYfxo2G+gGr3VKgN0A4Z7MTvrro9Iluym0n7d5XFFpDOC1/+QYo5ONIE7
TSFbnxJYcjCxWciBuNQDdiGVOVnpRMEURrettFcG/A+MY9soXfbZS55tkfdszQNrlYqLofnTUcWt
aLuOch0vaRgwZF6f6V4X23P2RWQiSwKHMFfwqHsCLuVE75Tow23yBB6ApPLnScMzxd5WqwI5IGp6
qNrnXI2ce8sQAZp4jYfhzi+w7SLsw/i8N/ymdHKBMqpH0LPfPiRjpVgopS8wzGhNULx7xgmuTfSI
7Q2PODJPo8G5ip3jMpka6evG+4A2QoDcnqzPL+pWBfgRTI7MiZVcRboLysVnKpzSJhYsrUJpZoCO
rj0l7j38tOjezR6kBIeURXIRLjmj53tdgMGl6ZN50NFAOP+0OEByiFG4mez2Teta5N9PYs1d9KO3
6UUemKP4AhJol8nHzT5VoqmuAro9aBp0r33HANjkLiC0vynXWYT/9o0hTnYnfhvTQcaFZFEZuG8c
f+KrBxloozlXkavGWYYrIIRYgRPlua/N6EtoiuVwY1JUDAgmo2dXeb73Vfxt5HjMZIq87XVeV+GR
tyfXBwF9GyN5bTiql6VIW21C7LnXVpHpS57ndzJLPjPDLU5RNDxpZCuLLQhprZcSFClG0hFbU/G3
BUmRc17RMRD54sXUw76dn0glYw7DprICmnZ3a7G9gNf/9lspE5IsId96xItEBEpiiVoNA1x532KZ
JiJubHkmylKt492OI/OFYEFHBk461q2DDWoWGczc52Q64Z7E7Xuju3PEtOrFg6TOLiBN0UL7WEBW
14CCvGcjZ30fcJolisYNO3qWmJfD3Pjb0rXXrhM2ERa92Pbbc3PyAEHLc7h6C4nK+N6gUBvluP85
fzF/rvgEed/rtJYpDwgNLSoenmGm9JJkNUTWfOA1bFTvdGBXXLVkeJXDXg3Y4L2HQ8LqIhmjJhtt
dWMEY3JesOxDDFuXlNkB9ZyaVsDuVrqm3L4TG+NjlAn1h/Q6E28PvePscMU0sAJJkS2qAbeeTpIN
J22XYgOBerre9nFD3D9Tl/0+BYBfvjs8PgZaui4T10Lslb7MeBIXui5R0AlUkEGJPMKJET1h84PA
h770sqq2O8/n7lMKieMenjgUAMkap25PhZGVILAHF9MuSQ45bC/4qdS5IE8oJ8pYGwiLAkIZLYor
vcAqzkU4hQJRcSn53J/gTV/1Zo+LKbPKR9jrWZKLYDCFbm8nRI80OIQhrFH87cTgHC4azfLVXdeg
ZBsZSjEvroCa5zmETbQUa5Bk4okkt9DFrMsdrHqYpm1CTWXjhxqXABWOXuh38DTz9/NHNAmcfLht
wtLTBHj60v48EjTV9YPj8m5I5XChvEKWA93qcmsYw7uB+0xCJzk5xLL9bhhI+sUNoDKC5mV3l//4
ku3sz4m18Tyzv2LwoUenNC8w3kOX40O/CI+KftEumyUnR+2+ZDTYiZXdFn+naSHuejGlHX0mk6sE
hiEIOHeL9ynzyeeeU0hfw6ax8YXsrS0JIthBfccyWKQU8MY8QhZhvbKhFu6u2fMpP7WQPpIMss96
oOI4w0RA7AUdTbmh/D5xBUQmW0EadnEdaqAGMKMtQ6pkOhj2e3D+tvVuXi7AIpLlFWZOw6OYfuqz
U3fGSnnZj5DEIUwXtcAgb4BafmLLTkobGkfrCmI2J2m7nkzvZLECgPEKzPJjioOPLkICXem2ibX5
hBVr3bzox5V+XAK+BV39A07VyT/JZu9qi5iapGcek1P0FKOJMxFpQyxLiQpe01VO5tjoFNIN/1+u
snLE1sf2Jt8GeY+uNoK+g5qSpoXv30q9mn42DdiLNJx95XVEprHYsVPWnK4tHVLazhkzdxBLWFWd
4UEuBy9klMFN/9z+TVnpgYRYXM7vUZiiQxs4f6fTtq451qV5D+zixtFxbuSr7wQxMwv/KTunkAg+
RNMD76MInZnTePPdzng5G8KjDJQLbfcWu1g2Mh3UpOgUT8G0bPfCztdTe6kXOZhoKfGWcsTFS4BC
Eul1zjlFRaJIyR/tIRnV9Eq3iDdRSlI1qNaTcev0oaSMGnDNLtcHkE3oOlkZzaETQCfWUpBxuBJk
t30wT0aTItNzPlifXaNyjTuD8k9CVzdf0Z+G5nojJlIq/SXDqBR4h7vq9Td8BbawnmLA0Bk61djp
vLd030fVElB4Qc4v3DH6uWORgteL4M5CCKNAnH7t9jFm+T2DpDUdHbdoSuL8InsPWxiUTJDA8iLA
vHW1Uov55iCoJ7Wj4QO/2+ze82eTeW92cJZ9VA4CHHB+L7Mnb+1o2Dl1nz/TuoAgyap4msltv7/E
l4hUuYnq/5o8zhmLuMRLLdevf4hXHFgtFVa29cgwkwf44HmTiJzFXAc4BRRrKGnMjTclZYwp5itT
9ugsORSEej1Wf4bpLEciWJDe02/nGuRcrntJawQbYHY4HNhX04r8qLWXGLaIfwG4EPNH1YKs0cS1
KbPCnVFfErl3v2DDbCzn1uXBtvyK/vU+Kq8DGgyAMBykh7EeVXcTE9iLbBGyx5KLEQ5K7XJAA5cn
UXPPy3gz+t5xW933GfAOKPkLSuLTM760Jf7eMWznUX/NBFHvQVV6XkutXzLVYu6Wj2DLwXy3r1hQ
NbKcIzi3WmPUfzL8R2cV/yesN2oIaRd0KsM8ExB4Tg7RJnJejxAx+80lUVueAwP+SPPFa6C0Hsye
f99DzTIEHEcMolPNFrKTJJIGB9VKifv2Y41xYyZghX/FZtQs4VfEWA+UMWnrOzinsvMfa2dsn2+1
cWZR4VHQsQC1jAwMtsr2kSLjXaJ3efzzvGzY1eD++uQF9Gmv7lfPaRiqqGDiS48P6bq8a4pBiI+/
En96MkbgjT/Cu6mwnge/ksHWwk3tTmKWZEnaTk1HKNOpaozpzGc6Ah/d31eKUN+N53A25rOBPACJ
4fHBYDM+lm95P17BMQ8iJ6ytr8OV4LX3bo1BGlThNbUeBRFL/16aiNreyAwgqJIS197Dd7JWn7Zg
GUV5Use3TpshBBBkNqP2LqgiLkHlolYN8EXsrpqrhJBuQ3CbkZNZLuSt0jfLbZ5+PSwTOWObI6Rp
MyB9VgtPFmc8eYTRp9XY6ApYazuPiuFGTK9f+zafmlBmhtEiV8fXFsIwsAvkGsV5rwrNa6+pzf1n
/SqxnXMLYVDFLxhnXXkKWCG0x3l8xmRiTB5aAwJ8ZuwRj+1fhIKXCEIUJJzCTatkLELQHDPECWR6
XvOAhOM1XkL9CsEZvDxBbx1HT2fMfX2CjRJr12mz9RxtNfkv4RB8zNUQ3XORwQbXmnWDVvEo0JUj
MNgBv8D+0aWTPCdUHSknrrWzrOn3q23oyzalaPYFt3fcg0plsV6+bzPoFEpQ9TJ8zutXtuucNvNM
mXYkvS/cc1vcr8wHnTdHkcnsDrOleHFeWDyb5eKjeGth4HiyqWiw3VtnGr8UJRzvuHsJmhOFxqkW
uRwCqEpxB/WZg9wdGuyKfZVHBuQ+CPwJzBMqr3kJXg/mtTJcODGruND61oFSqta7g5SkAqAj4pnI
hF0qOMItFWL9Ec63mPWC9fsIAxSMs9i4pU015g5rUjralSJsFhYorz0iiY90PfhWm8OH2FyDqqQI
OtHncIPfejbWTHyC2y8ExupnxxZYQd7riFBuUShVUnsNkhU8VXOsoLHZVAoMLwthwO0waoGwMqfH
NC1W/QrXjStyKs9DCHMYIEac9QHUyaOz2GIW+B4CdEJl1M2s//d2PQ83vPxHor1r4GR57W8RIBIh
O8y7itxEvbgCa1CF9yH3tMdf0i4x0GnDi8HjQwKpkxXLMbq12Z2sr+sM4B5mETtKpN6s3HEgxM4Z
CfrFSdhzmoKb6zy7lSTbT1yQIOnyE0Y4Di3DkLbRcvzhas/NrLZADf4ZpBN5NGPP0EwfCsa24bJc
egR6c1SAz8x9V6cCt6svrEN2rqW/8jW1T9wTTKq/8OBW1SIDmb13+pwmvVtdzzZ1eu17z0hqToin
IzPGmnknvI+6qp4FjXydWupC6VitVzqqlEdUXyleODTL8wAJl31eTlJAo6WKnieyQ2CB3v/G8nYo
WKGtUkT8Vk25K/uEJmVt7758xCt1uhPyfbQUTGQtva02lA1gRBb4EpGZ3NgK7h7AcQTJxyrGZf5E
2yBs2V0hGX24lc1omMPXMygQb4RVwLx8p0xl1aXg81pSBRyA4DudBDr38KuWaOSSNttvCfD4TGuk
EjAHXTLloC2plqrdRJ0Nj+YZMi6it2YR1NXXMo50P60NHmOfnZthLE7rO3klxcNOIoQo502YeFyd
JL6qGz7jHGdILS7ZmK6wpVBU0Z6VkxgWhOYzt8TbLFJI8+ZxJQozLpVyvrW5Ehv95M2Hx/aVLgr4
tLhetEA7Zf+EQQAiUYUlYQ8ikIrwLFXfqKDQtPqoF4EbgQpGVPUw0vOwXehzCqfBPiagRVnKHtQe
f9sZR6dyJbrzhMnY4kZEDsq5Y0YMCyM8xu/afSWu0QdpnPdN0VizcdZToH/dUoBG2Ja/8vjtpvHo
xqbhYNviWgpbN9s+GXEWjHVBg58JkjrW4elRwk6/X/ENSCZzGVRtoBjkbElNj2ja9chCSeZfLfYa
WcsVjCeef6LrGHIgyUQWupDNAnzE6lgnvl2w1/Mk10JA7wIUCmHV5z+O4ZyoJGfW8wLjVm3Zn2Xe
hT87qN4tMblRPKRhXva6IC7vJWqhd7d1wm3G96Um5MzSuVSALfD0ZuUJxvFdHsk3ZKMaha+kGK1e
RjBzJZcTDDpXy/+uFMoyCjmY9pVum+pWhexG0CvR2LFeuBdyjgxAj3MHeIuRb4MINo9rFfU/SsuT
3iJDpgpdRKi7QHjvktXilCxbU3DJwx+2yjb6PsAPzjT3C1PR5AwB9OzsjTygfJtjV3RkrTGEB/IR
PfTaMdRoNkHPJaX4wZJUjON5dyYcYVntjfUAka3wHXtCpQHoi91+Vnq+7hBtTfvmK1wENnRuEowi
C3LyOMouHPTsaq36dpWX3W4eNqIBaCBTunLOb0aZF3MzfT/kZmiHq4rYA5nwR7gqDg7JUzqQiEgK
Oe1QuAj3IOYwv+QCfuWGvD2Why6UKY7mwcKgLtiEWj/P78/h0AZTAVBj/+yNzY9XJkI9z58JIZBk
IbLxpzMt5Xrrk8RNJ8xTQ4nAs3N1HvTGoLR6k1EmkOPefGr9+2CppD1jr627Ue1z9tCMaRiN8Oqr
o7C5Pdi11UE37SR6LwL9t2WPXuXVBcI0vuPFXx7Hm/i11kvxvFtP/P9nU9OfDvrTq13aJgIUKTu7
xf6PG9K1/A0adNi8bG+3DtJOQnNBJKsmR+Gc3UvIJHhrRXuCnaPlukUXVp8DDb98gmwDJDNOsw5q
WokSiSsS0yBSuAlJxIZFuqjicbhXIlHFVGKHBNHV2IS8sgP7xqEO7EGuDgVAl0a9/htbpi/7mdZC
7D6Uz1hIdC0ty+/LOUwTMkoYVHzZCApHkZggoL+93uxUl1KA+tMTa11Kg//nLwNlDTyDF7ndMw+T
ai+txfICoFVuToepOrEaWyhp8Q9wpWVpd/JDvkqfMo8HfgOI1JLQWasKtfCe0Uh7zvOhRktvYhU1
W80ZR/cqBbX2vnK2dWP05xALRQjrDEfa+VNBkT6Ekq1sn6lPro7f5fckUlO/nwDlGsyfi/STZXiL
G4RVofOqrvN33YENErs2twexIqDaSSBaBqcpzb3MrYbX0qBNYSEzlb/GNDH3mRXUJ/bXPxSOr00Z
X3Jl7iDDxwLxmedFtRpGu7CVrg7aY5w6TNoPnpXZOBbGN2iHGcrYYiixp39m1LD6Q5MOv8HaOQ02
MtOZLaOdrj4Ce5/twu1OZ1UFtSvO3nGbgRwFJuRRQFboij7SFAIJwPU1eMG9J3oMWCP3TFUGQL2V
kqbv7NINu+ZphKloUom+Io+xwAM1eF9cY4RBdGZQSOxLJiYi0nY5SccIPKPltx+0PvBOqQbFCqWv
IkZhZ1c9uk4UWkhm5cujSE9ML6l4JBFm3MVKplcaR6+8m83FtB3113RVes/DkTpfVO3oV6Jr1hkX
PGxluysG6trjaCMnM/y3tLsBSZ5WTCJPbi/KpNsNRDzkP6QwW0+yK6UenY9gHjIUbtQgkBz/qSNa
cyxQ1oMxe2Vz39rY9N2wS3mEmuDawjlTYs/7AUHieFsVuGNCkqorFjPEXRjjHuX/epOeYhep03fq
LfFO/ADAK8Ufq6LHfo7V8jRwuO4LxxNwIPxym1VM7IbqYwEqIQTvWKHl9j6Ttcea8fqUEKWN/zSt
GZBFnnKoeb+7dTx3xbNN1fZCjs82/OSuekyZWJZ8n3s9NsKqfio4VyG9SbLLQtY1/Qre50o/+7q/
tA+5uuAUqKVwPFytwm7NjHUu9B06NxPdUzTRzSeKWwhYgYJ0R93iaRB9eXkYKpipSvj4BXdiqWkV
Yx/oFhdlcxozq73NBrGHpGZm5k9+8nUp3s7RKlOQCfIW49nQh5LHjAlrNvrZC806t8Qor7CEMjof
Z/Fg6jsoqtoUWf1OAe4wVow8etHzshi8zhACLz3dxrCx9RdXRFODyappHlISFeikaKZXU9ntHX+q
X6uTC0zhlUbv8lokLhogr4mmXZeHWx27QLxAe1xK0DdW49338Eh+WOy+A2ScBZa+6yrbTYEjo9uR
mFR9WD27EDsqkKlx1LbOxJc0OadA8p6uQ8kE61/bp+d0jbxXIzU1YYErsE9WUGwjjVgHU/Odg/UF
/PmlOGkcjHnAcEXXNMC3900IyxaSrpUgyGjPpcy+WokGv2nFxgjHuDDRwPQ3l+77XC5om72kSxLS
eguFGrgUyEZiUl7LfrJqMvolr4ODGADUyECnqT2JdVWwxFPDIgFQiUCSjJ8cwK34I4R2dozOnlNf
YchG7FFF3+wh48I9fQTqtHGjb9FzRwqp0LuQbsj3KrA5/cwIe9DV94v0qz96WiNwF9OHQGjPRALV
E1C+cZfin/MrlargMT4bOmqSc9IOHOVxrq0kFzg5GMx3bfehSH2wcM3SrbPtK6vcIgEkhhjJ/6IC
AvFdD2VP0dNhbiJchPZIuOpBgqV8JQRy0hD793D9DJKpJI+DngY2lTLR3AEhjFn8TektKs29tv8d
v3gvuq8Shj+/i5ka2iX5wDhudbBIrFyhaGZ5d6nRhXB3F2+b52CUqlgBBmedzTWeCWH973uK7JIW
9A8d5yk8YjgDLhe6xzIB/cYKBaYrzf+EppIbC4kFRA/q67rLRZSbqy4FeMEk2QFILsOAk3ATe2eF
PGnlHhvg6RUBARMaAz8eCO6IABgpQpFy0VAAwxwJ9+HQWpprA3yYUWB63oJL0hIgWQgLHlz3UBTm
A1gKFuZm4Q8J6B9uG5ohJ62OGePClfYyYOJ8zAwFyQq9orXyVmWaH6BaZSJ+/SGJPEEYFZN1Y7Bt
FYz8kzvT0HWBtCHjZ+hxcP8NveuK6Bm/YDy4YRo6sjMLGIwJ+ed5vmEIxMpVUpfZKearDUQVhOWX
yaPo4qXthJPKhhsVuZMkD+ExpUvZ8oovrKnvTuErtLjxyMNQzxFwXep4c9Wdwp+7G8BmPPN8Dm6J
iWb8LYdETNHC8tzxptS5K0O1gom1yQOBbs0x99aYoa9sPwOVPZNzxp8XwMNKNz5P0Vi4JMac9hVp
8qqF2pALzUlaATAuyyuaZh97FmUYhtu6JL/ksib/6/HaqHdU4b/BXBHwIe95XOGVXw3CbRcnIKJv
+dZhLzqheAaNwQQTJEBBE1zCeulH4EQpqorVbDQOM1wkKaWieji663x+gSEK8ZaBCm9QI0TCMBXK
+MMVA2PVTovb73X835LUlkt5PXErl6BhGnPxP4zA4R6XAhnTFsDDMzMSHysNnDWuXO4xOr5opgBx
TlYHuV63IZ6kgp6ZMmUgKOVXGaswyMOy5VT2sQ+04PBk/Tnfi9zTuM8g/0l5OjHjV5qhaaMGA2pB
9io5yQgyvtriB5PbT4SToidqV4XZXkjB5Tfv5ZM1eS/lVv+d6tNo2Tg6+l2zYJO/eX3p5SVeJVU6
cUS3TP3f+09/vVxcN+l6FjaMJyl4u+fAslyCKCqh3g0zQhUyZII7upVRl/k3TBrNjWsrqoifSOhh
NFdDkM9o/8Q1MW6MDersMQzqqEVZxbmmbfBmMvpz0XQsVx0pCrhEGI2NT5WR4rvVEUARQIXch4qt
CZCMXriq08MoSFSdoWP4PKDr/M1olg1ibSUaMiMreOe3jvB+MACzh3DXJ4Jrun5SskzNnKobvTGY
LV6JcZtG3aym5SbJt/nYD9sLuG5PLSt8f4PtEMIpaUCU1ZY0NGVILw2p2YnZO+aPRFxfgz7Dk+rU
hWeZOjNkUFvysBt0ZAu6ww2p1tvP3kS4XSdQybuMVVdcBsh6Z3GRQeDl4g6UYc8W+MI9Ri1y/5KW
ZRL0qEvjb16E/pB1MB1IWBu70B6V7RvHAh/7EBK+glSYgawyIRvPH9p38XJRvMJ9PYV0KOArGrVv
0YvRpWBbqjen9DHHFkJfSjvg/3+Dh/rUUL+bVOHp3lcvRzk/TafFWXpe0Qf/fKQKU2FhGdFLGX42
zcMi+LdNBvGww2jR0WBKrw+qDPlS3qcqWtK+aHFnfAWO3+GbjPwls+8IutX3di2FrXsYCgfJ7Guy
YxsXwoWf3/csbfZmbSL4+ovGfnJEyoeOYH+DDRmiGIeiPwuZ+ZFPRFkOyl2YCE1MzMXWS0/gE+Ah
gDmoSgqZjWETxrrGMjZmu0rZ8CDK3uO37YA7tllLtmaRNbpEqhyOwa7T8dUlkAnSYFea18SuoB5K
Ee3lkSkrKBe/vd+gZ8S3liAuBxVWNoZS8aUBNtP0dHWDRnt+QhFZa0n5Cn99pJcnA3wNTLLpCUKB
s8lx0lR4/bHen+ch/vildRrJvCVgWzDEspEDt1q4eU5ruUuWU3HXVE283PH6PpdY9lBLlAYioP+h
HZIJ01bNWE2aEiEm2LZ2YiEL5wK4mcaq6AHDhrRGvIQgzHoxn2uhrML3D1XUQ9VNLAQSzyYLG03X
6tolMWZKVNqGfMiXt4yqWT642VWxot7sKf6gCDBgjemO88F01K2IWjdBBzIuoRy4Mr69kdYBioMZ
KR8dJIVNQR9Ri/9GHeI+Fd+8O/28O0CKnM/4TivXouJSNqwj/LiIuB5EHMtM+gpLIFssGlRBFD3D
XqmVfGIDt/mGd4w1Z/C8kNOkSWh1m1qYW5k4BOOomIj9p+59LVplhZsFPsR/B2uStT7zPdD2uhpC
kIw6wdM30DHiRxt9OrmaNWsK0L0xtXzs0g4R/AOn4g9BBRTyJfLY6+CT+2sPh6u46PfsTni4hG81
2xKF1xYNpMKvR+nEoNQ1R/MciGFvwb8vMwx9oVhSgevUxKVdiLZXZugc56U58/Jgc4+StnIFuag4
qyluSJaiddEUSrdCLBbgb82910eFs+jaapGW6NRb7VIQ5EFloAbSoIeUUUC/W9BBchdhW3QeBkVc
fZFACgfnG4uPUMWTJIbDOo+104o9vSextUXaxLfGjVAyEyvhLfuChL9J+d16Du4Yy3P7j30/NYqW
UtJqLMgqXLb8dTcwcwPvBlwTXslb+D/+BUUiqOlhTSFme2Lap6TSGfTp3TCOr5KezQrfo0zcD1Zj
jxUmuZFi4MROC0tvSPa3evVRyiwO80qLJ1KJsPkzJ58WhrTpoa1hLSU3J/M9F52PODmGJS68VKaw
BU5s7sLKp3zqvazI/SM+W48b77hP+TKZlkyDNV8kcmmnOnnQDMAMd6CCxtaKMhxb8/gXQSQBMM4Z
j2VzphKn1z3CIUlrbWKAFYYV9EQma4Iy/CPAbQ5lZcUJ0dHnY/dwDpNbW5g6FnPG2R92LtwO5bfq
pA9m7WHHELi5MOTrnZ6wnFqFkYpjfbWv4VGBTvQtqQBsgie193Ln0Xp7PRla0eaLAUSrQDq9b0Qa
UInHm1j7IQsh946Vqf9ruqkAEzWa0Ocpia45EcCh8hu6lrAW4K2znacMtb7GBfCm8J4/OgDbvp3A
TvpZF9xeDqnf71lkkdbCqfv3wGsanhaD01DGAyY8UuSXNUOA97p0SsOEHDgBbCneSsf6THWbqLvJ
shvm0wVnZjwIJftWy4GWNX6fejM43xZv8ddKSN6Mqgm0CZVUK2RXosVSKznEnqEM4oTJ23IdIWeO
EIkQJ/6Q3GFhtmW37JjS0u6YuGUtQ1rmmUheGVeS/nWWNyt1wO1K1IsSGi64mMqQdYbKKmFrUtKk
s/GyFbrWiTPbFvULntntcUZ6okfJ1jxFPqRax1WJTqFdygUehC+MlBH67n0gVWiLC+Mq8qJ/duzZ
QhYce3XMDYPo9hG07J0Wbbjh4cM8i3zi55NPmIifIXOSs+wBT+x0S4Ph3Wn99A/q+Ej57/nQ1xD0
UZ9TfGOGze6WXCJZFhl8hL5zGmRmvSpvsI82MX48vTf8PgtpFmc0tXuJKhQelbQykupEc36udU3y
+OclOvxxEaHsk35c6k9GwiSqGKSo5ob1k/26SfwwD4a0Njg0F+3S+V3gF8UUMyhpZOpzFtyQdQRL
BVCXFatI0Etme0lRZs32Z34cFVTPor6NUxiQk+no5Um1fdbH6R2YXUC2LQtGkpkc1ONSdkNbMUHf
BcZ4a57j0Pt+1/Mxj7qg8Oj2fh/NwWKcPcA5nZUuq8h2XLxYwMMide8PyvRhrcJiKL4hiuxvVcdX
m1zx3bmYZaXoRQmXcmHHZXXwtK6/mC6qA7NR5NJshtZ0om0DYst6kPrLCQsisnaGpVcx8dxYmF2P
5hAO6Uaz8U8VU/h385OWjjWFp2c18FkU3qadrCYSLXuco3RFHKjcXUpc7jNjdh2PNY7tKHLWFjO9
bRtj7BSmsJIcTDId+7G4I8GJeuXzUT/3SVQAdeaWoDWDbj2c+CnqVqPNe7rPQmkoTaJf2geTRyJW
2iM0j0xgeegXqUUT0g3fjN5GhMiLi++d2jLLiK/mgOj0M62cp5qopXvZaXVl9QQE+Z/AtjWukWxb
jJqdXIRkEjj2TMb3vmCcsOaUtLfNadot3cHOCPrDInGCsxmxEkd6cH/2+G0A/TonqnCg18/PAlId
4R6ugtLo10oVmalNqrxvKwV/Jk0Jp3JJ2hrahmO5aqc156WbOZ3ZXYY5IYPzUk1IKsk8NS6hyI71
nEgT9T55WwNvW/pHA+6nZht2ijSm9VhSVRNrzdZlyhfxgPUh15CEU97ZkbNAGfGGvuU7dbcfaFVC
tHyWBDzy3j0GRd3xlO7zljOPPV6EylBqG167MKWhohgQe79Q5GhXgKtU1grIKTW9C8zji4Gh1wvf
Ec/ROAA1sMMoJr9P8hKzSRvfHlFk31JgdAibHh3ra/wVvhXxu84D9h0Tl5WXO9Lxdieiug9M1KkN
Snzm+xfKh9XiGrsXXaFIa28sV0kOMkfRDZpKkpQnXTapQ37XEeSDFT+vpiYh5pusMXLTL57ZX5DZ
Y1bFg0ffwDKWEGlhm98MITJdsJ8GBU9kS6YcIDQJUj6iqFcBGZH9Nd9nYA9XnUpOeSJe2RhwZNOl
yauje11nLpVQt4dB2E51cIS0p/e9B3GyFMu/SSmNVKtQ97KQAGjNJtfS9MzQlOmWzmIm8PXmXaS0
gp/EYV1jULtuwSYq7G9P79i8VhRuYbtiNRRlZCovvquH/y/BDTZib/NpDpxaBeSDrxgtn6EM8W2A
ySD0jTVnsjvbG3NwZTZlrusIEtCWGkKABhgky1v/975kPGOiA8LrYOiZNNgM988twcb8crLj8Egy
7Z7CipKcOktHO+OgqyrxA9v96MYzAArwYPxKjZzRS3fRHuslkdXNezMVwrJKHrSMoX/FV62vd4Iv
BaJpnSdEtCki/PueDR10y6asQ7nSLr+1tjvZBsnIcVsqLIwBquTJ0LGB+5C/pZm2Lay16r3vtUYX
xa6/U/B8HEE5WP/xS8r6OWsoA06xZ2ukUreh2wz3MnUiSvTVKEF+Wmi9IqY95SdP/3OeJMnEFbGH
wWeEG7kl1nNP129AGTO5nmu99ecz0OUMtOvu0cy5ymsiS2M/1jqt7gm7Xxgok8hJoZ3J0Kj+syQi
Sycn8NZBSz9pnt6QH64Rep4hWENy7jsyorA+QuaFrKz+WnJ8mz9cLT7YVO5ek02v5ZmJYZYDG3uw
jWxdl755uhTUMqFgCTV+sF6JeXSu/zgDi88XtQiELZtqJ4KhvcLLLqnl+c0ycxD6XvsacZYJg0hx
BQvNrDhffLmgxJ9QbMs21Id1W7mEqdW5/N/N9BG0YMJMMgvet9QZH2RkMgFRPjDlGr6JJXX/rl1J
fO44A8CPM59kRb1eAlwH4cVbNkefXqjB/DZaUUzAe7rSrv9tPqPWyRGSsnhE9euAhoeUe029kjEr
GQgsj4eCqOC0eMlCLANvkxSzymJIHDcZeH0ut5b6w12PboQbOZJqoaltuXKg2mzsRJIhO7hjfn/D
uJOtKDS3hU8eKXCpCJEfHtoTV2AkxrIVdKDbPHSA1wasmlvphhZ+uQ6ayFcfj7vMYInDbxTYjc5U
WHPZYkWJR2WlMOUoRhF5d6PN/kKVguGv/ZUkYV9MUZvmdPeJFD1GQNZJxDCzdPIsxggoTH1/LGgZ
D00PRZAQbTe0u+768u/4mICAcYxbN2Kux3IWqEZJFKpnVUJOsnC+NoaSLrXJ6pKowl70vmd0EWGx
MNMELkoHQtAfr8NeCbwFXhF0u7OLCsbo/ckPRbtqK01iZEmFv11NLCdnUseLnkI/uPaS2B5kSch3
z2URo00ABeHZ/M5b+N2NHXn4Yl8nyaShXkET0tzNGyXtp/X3o+dEtIhtgBnOF4wFgKLGb2T8v21c
Yu2UNLmE7CcgIU7zNfEJ84+spO3SKXXOI6nS3qaXmLhw8yMWuAFgf6U1jFd1mXPqqVpehKJLYihp
HYQfT/9LV8INiUXzF3bJABEZd1m+IasjaEZ+XI1aLizGd/6olNRjqyAftke9lbbokFPL3KfHR1Sc
EELNyip82Gc1NPkr1pePxdZmagPKj50xkqdkatE7HoP4VuHf/Wh7mURySbz++3ipBWpjZpjGOZqj
z+37JjU2t5Mf0kdUcQTEJPXFccouKsJyq2m5y224nU/Eos60GXwvum6Z4M4eHX/5AyHIkIDl2Ibx
+u1gCdc6R4WgvI4qLwnEKIyXv1AjbcAjJbpC4rDMwsiH6QZJLIR7kpAruyFdi37z3P2nHsgnvSpA
jLtz5rjoRdoyM+SGkJeD7WOvfDOwehp0WB3P1MkECkhIaCN9xaVMjZsvgvA2ZFko0zPXvjEEXcZy
A9UgbaenUALi7oyGY/3X0QDkoMXJW9L9bW3aHJu12EB8GihgTRkaWyx1Vsqpd3H+M6IJueM+N4Gq
ln1f50WL70NZzuw1/5gTbRGQr6YxfObn3jUpuA2Xp25S13v94r6u4xivKGh1YEKYVx/3nqQiKiT1
27uud3c47dUGLwyKe5N6BrR6yqsvc2jnCzyH7NoL4MVjZ8BadgUObKdTHtEViSp7M9BYsskCFIQp
WBdPjnZOOhAJfGjRcIojRYn7s2iYJXoWRqKTMMVvFDjZmRZURTIOEIS+4w/lJPQdYiRb3r2QLRwJ
2/1h0wboPtBRCQf10dkk6MekRWlzCdza0EcDVhDg2JRJsVS5STC92Zx00a9ARu69VcXXlzpYxsXE
rlzuuL2YeXkKjtGZIrnr2Xk9vj/tBpGW8y8jxiH3vvx5pa9r25tJvD8XZ9744HxBzvkWp+RaGtXN
e51vFQr2ztJC0IlnFrMNbjxIgv0yjTFQp29WmoSSR8uZRh4GFNr+q5iMb3T9+IqpMOSkJSyAUUKP
dzmG/bLiLd5OMGHg4wPUFbseUsinAhc4K/qfPmXRq5jSzpob6OhJa9SeHg/2kKMRwuXFOQlzLSOH
1zCtIE3+RMP79cNn4qBuyKUwvuKaAQEHoUXf4Y8i+dJBxF3/Z8JQzdm345QC4UZKeE4c7N6s+z0u
ZuF5Q5XBAzM/jo6+Yo+1w8COKuBfQhV4CKz9w05jAtxZzOf64SYL8qOZdYQ001Pdexb9D6nOiXSm
SHhGelQPqwLUZMEA/MbeLCEk1uZLuCWq6Zn1U48/7So41I06GRtu7mpGwbZjjjgf6zg7Dxg6vo/k
s8MmGhDzPGvd5r8fWvIozsz75VCRKT6LwfbUQLyvaYorICd/OKyhlxhcloMZTbKRGdL4SkFp2cjZ
OrLwkQC9K47Sk3htrdh3B2+OkuhGsRPn/7QkLEtcXp+rTLKqJeU93hGnLipn9UpJrI5IwSyAMvC4
+ZCEcN9Pb6StSpkvoOLNgk7+ZTtLhGi8DWc5ttAOaopvTg422Zo5JsXTMS/AgpOnmpRaIlzYtTAW
3WYFTKqnGUcSWxLvjwUcdtW4VlIOrTxbnlQHyRsOHqt73fbZPMXWOqeXW3QcZ0MemRPbfby0Ymba
PmPLqHqrE5b4Hwzn2GgsNrwPodA0b+O10TDaKELBhmTqrztiuRdqIO0aj7qFZb1wbi5dNyDhwOAw
7wMkj7D3EeHGhjlPG9f88vQWhs99KEDTby5GTsUiOOgcY1jrmZNynUfdgQlRPhjLtjHb7PTZGiMH
Aone4OaVO9/7qtwVUhiJDD/+J3L7xDH8C5xKHBc3mgjmmWE31yQJrNbTYsRk8inQFbxvqpCKvHVZ
yKDj5QgpXRu4xHQ5I6cdxA67FGjeagK8r12dLQYr6NUycrvp/nLzruOEM+KNNjPoX8OZmy/BXRCE
3Tc1wDlAgorW8Ze+t/ZEGABbA0rzfnCldRcr7e+CqM+OSta93wLvgXBg0xfEagFVpeehT7Tw6Geo
j/IFhhJuUi1h5NG/j3Dqg51Fr+xYlrCfCk8Zk2exZNaQGjUTJll77Ub6gmvWsTC+452C2DiZMRcQ
U8yntxEYXhwr9OLHDwblWK5gO6O+QvnZ/EU3SL+4+itGSz2aJUftNX/lHCiDapg+GGZaTO1NQx4e
dyDzN5WyZfI9Pwtagjm8F3Mq0afwKXLyKecgiX0F1bdiP1iT3HQc9cKB/QIstt4jXkoNnERyRIi6
JmY2fQzZhoboSD4Ya07mKMF3+En6NBLG7HOeC7rSt3n5ZJWH5CpHBWrr4mlig7T4/QO/ybM6OS/l
TWqYMsWcyNQTOv8hstUqREAg/tWhKXhLyTcRquLY/X2Q5/27FvYDgXOxkB2+zRq41ebasZQuyDjG
dG4tKUHz/a4fMxAU82JxpzxBs7oId7GVcZrp4UBqEo5bAt6TnjosXatZU4WuVQxS+8KVCfGZapaK
6e6XMRvRyjU92vmrInSsPxjC2OzoNA+YJawcDgrgvNnHR2IpCf05StQsm4QHYRlrIlVGUOJ8knID
KmgUgUGY+5kSw/ISwmP29fiDwAqA+ROLnVrw16/mDIFN3wqqZ8D8cD+/zMNskMZ5zmjSCMvOhSxu
NARr7eqEnJKQAnYCRpHMmC1w9OY51lpTf2YCVJrx+t5ewEbIcHqKBfXGvSbX8wbbqDg7dtV3/H+E
kjkiTr0cAaaZ7SXt0xArnRebpFaCBcB83LvKj2fJJZWoRIkzcCZKUSgeXEax74A9V6kFzO71N1Gm
BYrbroboyjGh2kXygDnMNPBTg64oiXVjohn3amYiDzKRTGykshRy9UGsbLCutdCS85AEHXxsUJdB
m8lAehoedNiVBpmbFd26c77heOKWFCjBJVuEpjhh6dQof1ZPqtK9tI+0xM4HZ7BkM7X6bw1eESkM
uO0KSlbCQJ+zSFai/ywxDYHFLleGhvPcinB8aRzrTtOYcshVl9g3p/QjoHqzKTi40gr65fG5xrfR
iqmmdZ0XTSHH/Sg0USWPyZJovwYxkaac4/AzekTK6Kp0DmXBon0BejIo4R4U8ICjtrdPKm1tHEeP
6EIEHjmTaScW2vV7aAvPyR8y/eGK4Pjm2AHXoWu4WRApBfi2BIt2n5csRJ6zuFXwb+vEeAgiLBqn
1XdSXifTdLxOLPBqqsFhsI2I7INEJR1tNBS5uPsx3zZtssz8L95VXxLUmmt5pIsCKZwr2e4KuOMX
5d8E5KrFW9W9eYpkMkG0hTcz9CeGwRaC2zpwuS5p6Z3459t3UPfczvHX0+nDLivk3k3p2VCsICUq
H/zyl4GoJ+w6VRlzPPpnq5EReXWtySTNvPB3PdFqVljqeUN88HL+ALdQVkxQGm/x0PuGgU/x7JGB
aqhICBlALJ2pJIUnLrEWPFzFfAdU0tBkqYjZNsFmoepcEikz8DFPFcQOFx4JPp+DAEB9+CvtCOnj
2kM0E5l5SblSN+WxY9qYDJoI/j1mQ6kP0HhK9ZrYqGhU4/QxdYRZKOQw+R35/wLz0U1tMZlJv9Af
p3wPA8JjpY1wBsj4KeDmhHX3iWQ0HqUjSHwq/bUu8uuHeH+Eo8PAcNN6ApbeaDPJg8AHDqtknncL
Ci4D4J30YH4cO0eSzJj+GO8bRm0sYM8uhbnQpni74tdSBbCbfQcwTlXtRTOw3kSu4i3e0jSehJKY
3aOqyqNRnvrfshzlIEw59XWLvjSRfsePEVz41jWSpH4Mtfj7qy6a+vMVcqFO2ZbKIC6NqSMVyjK4
N5iUgKGWXTUqIitsEv335R8Csoo8TDMJme3lvQuTaaSAM7E+RlCMdB0piQlNTY5J55U3b83icMl0
p3QHpA+/GBd4FXsraulGqOxW1NPdo5K/OCfP/RlLcgt+SYXzJtw9AAyqGh4PgoVn2ldw1mvjGh9n
yUb6lF5HaakzuCw9zgljjlL9IZq7nsbjyXT9CVBf/zaGGXNnd/JtFSNlyhho/4DwrZyPSwdaHhzm
Awh3rAztdJnHqVCcGMY069IJrlrXiaIe91bTjEKznvQo75Iodx+GWa+R7PxonhFzn8MJEbs1tbY9
F2WZHLAhMObyYR+0FehNRS+P2CI7dDp5ATedXQf3vTA9K82y5cYNQKefaMefsU3YqA2qulsoPw2r
lzNNJ7qnDyKHC8aCWpkaSRqnKvTccnJQSLJRpHnZdP3Kvxf6HQEx3furGMS/X0qmSI229YuuaZU2
WuAXS+uGLurHujclR7XXd5JrGZ4YGaPXrs6OGlopniooohOfK+kHdgAukJQdf8aIRbdPA/dVjg3d
KeLYKTIMrXgNGPT9zN/JfptdFkjDOZuff+wizbL1XhTSGlAZNxRVSiv2laK2/jsTzHrW9Ow8RJYf
qoR5SRXmIOfGSxVE8jJiS/QmURmoptclJjfr8U8WVGjoYcWRyeAUFUCk+VQwTmioJUiykjM5xn0x
4zB955N6WPgIqceP4SxDu/nRjMaPmi1lC41yVwM41NDhF9pkjW48iEGhBitYLc3tmTmew/8y2PTr
jZ90vmR2jl6Yxr0BEZSnCrLwgZ51q/fywb6nGNd3EVfkY8lytTShbIl5DzcvLtErBUJkso4yiFyr
Hxv3VrU5mGyXBId7wIsAlpyVKGGGEyYtX6lSqkUlrO4lRo8mAlsvn84tPwx8JgUTmOwCD8QdXDKC
at9NtE3WdpVSKsGD7x73JY7z68DIHpg7ypnWtzf9Nm1GBKo2AQHu1i1LthUAxy2fhLEIm9CBGdU8
fFREy+Q/hGLjglmRqldQ/S918UlEm4QJYL1pTuRNWIOtr3XeMfA6KOF43UuT/rG4xz9ymHBcKIm6
4afiPGz5vB5bI8e8226itTINY8tViNNj7g24nsskeBbgFbWhYwkHFi87r59lGJPbDRNrPOis+56T
zoPzmGdoxF32b01z6OIQPeGlQ2X4bQAE3dmSbnXksbhG+uF6a3ueIDZYdNILTLbzWt/bSOidGpgl
1a6joTmNRgWzA0ve3scL+C29hGjT/uPT1+NF7GWk7aD3ua2sUyVaLfX6Lp1eg01+gnNkv1ndRn29
rmnGnQRJvyXWUTuL0fWYks3u9PC9wLfdHMzEClCstYt959hdTJ/PRpfzza+SAIohdgn6fORHZCtq
OJIjFRHujVCFu6/ssvbK3Dott8PUPMaYpqRWiY8/vQIpRpwlDTwuupYP2zONITBAVbhC88/pq+3w
O7wn1X58cmEWxk5RDkojEAB4vAqc5W4NgiDyoHX+EUh5KZGHMH6pieTlFHzbT6oC/w9I2CYYEpPg
SV5uT0X9jPfhZEPmknd6L6zMTUDhk5qaV5971TtNzkq4JIy2ON1mNmB4yHO9X4BujCLiju0MAPRe
p/6trDZKq1cm/H/jHGo1D42e+vkvK/gbrs9APfVJ0LqB7NEuJf3jMaLUKZ3FS4mwhzZ18PCQ+VPR
gNX3IWcAov7dZDEFv5kkI8f00wUahl17t3EWJlt/6vafryWgYFb8yL1N7THZ15EO73FbRWbG1aSl
I2xfru2aP9jYzaHHp9dKC53hGm7ZvEMLy8+LMo8+LSGZuOBEAtUBqQoNqvEtyHgnbCCq5i9aST8G
HSzQcZNKOcVEQTg+eJjoQdqjVKPDnpdfQ98aC2CglpiIKD2gpgfGBzNAFf01vq3/h9vu1Ya1x579
gLqKzP1OTfomFMKJmKFZ0k4glVLaNfvqyt+4J3AKYl5+UDFVAR+8dEBUqXqjmjvdtuj0CRXD84UZ
18nIsyCVBkTO8ptAKGAXiY2OtlhrMKH0QctmePy6WAcr/AlxVOrQf6fPFsnaUQ/ESugoKKDCSbHV
9g/87SmN8Z9/kMAFNUhzxaQpYPg1rrvXm2pjw/l8T5oPONV+iO9SzFfRORrXfIYSztN61H2w22k8
AaXKC9LTbd0Pgz5X2wICbCyKmX3vWd2MBhL6Ahf+VOdPwOWhAxdNDoR0qCOZzC6xbYj2GcKhJtno
XsIhzj7MyeCiazcfY+GtWLJ5U7iNXhz7dVjz0JH8TrxM5vZam5I71xEZ2u16RxQPr1RI2BN+6lJO
T3UvNUVw/fqIBl0X0z8A69wrojEI35mnwesNSbpbPdXvdlefeNR+vxfLHI2P9B/d8ukV0eyTJ7f9
DNcs3f1IeBkIYTmD7028Jbuwf2JqbsG23Ja92kJ6iro0clfObALtzpJSF1O+pqGIq6GWrW/35YTW
5FU3dt/mupg3OgVKxYcPq0+5y8wxyde2qs+xLOsSxUCc/SLTGKksqIWAXlkKeqJFzSWjuDn2JmF3
Q1sSKIzNauCTLYMFfp7z3c2N6CmcxTWeWl+H9fvHxDucubgNP89ces4AOAnmBTMavClXcLDPMTV/
MEVD13mO1YxpUPTQ0+urLJ7JlEfSVLyg66Sc/zSuRpxuJY1IlWXB9MLC8HbInP7WuURJ7f45XNrA
L9N9rZxKg+k8oqmu0IOC8X8Fg+YJ0WOO7+6GpszwbM9+P2UnaC9VBMr2EcWFNlMDe/54ZKFHxxu2
9D7Tj44c1fqTPxAJVw9htD39k6TBJWjBTixhM+60EvRi4bMmdQepWbGxj/KI7+H4DJ2VEj1Z9zm2
bhVRrzVBVwh1hZjPuYWrAsDaCke9sSAoUq6wC5sFYp8PLbyNN2JPDMinViICeZ04MzX+jdFq/dVk
sMdG6F71f56HSjH1RBvzn6naqMbByDfTF55oOuYJh89AQrnidev+aH20VYsw30P3AcDNHANaR97R
H6K6xSTEJuJths4jTJLTE0rd1xitbiQhalpzvJH5Ebs1/ctW/ekGOAK6cwyMOzAmnjLE5EHgqMT2
cvmLB1Q3kAKbw0T9Rk8x6Mqgg8s13Ez4dyetNKtht480oJtI4DH4hEHWgqDxK9Au7QVN2UnjfDuH
iZJpqguz2F4SMPzlC+vX+PuXyW/4FcCuRBl/q2L5Vp5+H/VKS/YZ9hxoEITgimfBv0rNgDYxqaUJ
ba2mHx4f1+Hw+hIU74OcFicc1LABagw0TURbaE8fVXvtDEQY9Cxs4XqqAx3FXmcspIqWNKATKhEj
HV/oAJWYBUvUJZWodYs2qacUiJN6cJ2dGGHTHDm98lBGDYaoMgckbIirR5Mg7rM09A/QY0zUndhO
yOpBwvDEEwiW1Kt3OBWbMRXkiMprajnhz1R0gNLzpeB3sIEmEtI9rBUivzB/7KJ1Q8hwAc25xLWa
W3PupiEbNXReWRLB6xhRn9RvhlsIswFAzY+zLlMNcSL0z71FObKfjjgxol7CoyORJHU6XnrDLj2k
xKFFK1BWfoHnM76A9zQ+HrxLNoxF4MZg0VCwOxCmDMULS2UofXnC539VTPukf9GynNXmwm+xzyRo
USPBnKTkhvwodGHeJdevmrRuW0AngOSnK079bNLaS3nEavCwImEnZ1kR8sJ7DvxePIqPnqwAjH0J
CwOpx4BEVjhUS+b1n4BIBjCx1KPE/uGjYViA7oHHeOWGrRmr+1UleK9PFzIVK7m4ED8ELjgowEAh
9595BEbeCc/j662CeIkkT6b69Z1p4awC6ypS7QnFo9q9ffHFlAYogaFdNcvhgHdschFe78qzuj3D
iEDzlztzO8yzGz5hDG0Uu8k05VYXawyimQTjv42eMkh5gcKtFLHX1UPJSGj++d5BhdCWIiEzRpY+
HLj0Qa3MEjafbXA0zKE3lICrtGj5G5mQDLHOOI5N+AH3c1ugbEmy2aaimzpiwNGSBzRrU/CmJTvp
c///oj2QizgCjQcEVvceXYU5mNHRhKFnt9j0Ck3yqHVSu/9Kj07Nx8tauuhT8TBCCMNZZzwn0MuI
Ni6ybmuIclWqDSCX39ghKO5pZ+MKPzyzdn/f/PfZCC9ILKVfJF6LNHwiZwX2zlb1QilMHFo8SJgW
CRc6MkoPA/y9SzNrrG+QN53GhqxypoUPMoNwuS6Uqm5iYekIPw34xK52tT3DPGc9hwfD+uft7aaF
J7QIBm+JA8OoYN2FodWLxLVQbJ3U0Do2FoG+xgENqLvgZR/a31Zs2KA6nWAAGTYcsucQhScknPhj
QrMhs9vYUB/Qjy2i7/UxTHQ3Nl2xFifjpWNIdXyTB7bPVwHzu3/0WtyMoQ8B1S+Tb0vIpGpkMrFk
/lwxnJQy9j7FpNZaRz1aA/o/Zmw7vOJc+xoDZxn40XBYPUfQzwJNZACppsmLfrL8SfA4/vL8TVPK
Jkx9tlI6K7y28/GB5vFBw82dwTdfi7eA6lxoTYCjZKwDyUp1oDt7D1/N87E1hB0gacdW9jTfcoVG
j3sDo7Ag7Amp9SZmdciBLKVWkNj7y77f/Kc+M5eZ1JqX7q7YBts6Xoh2C8SDQVLDeG8lOyOrVg5o
cf7YyXvUILz7sgvqZ/wPInkOqaTXkXfzDVvD4gihoSNMDxlfsyAl1Vpe2vSPzq3uLD+ylNOg0pVt
QGpVAvdgTu1Da4vHuXvyFae+EcDdwk41uZXJTQMXffhuA7UqAbhs7L1XW0AyWYIKcCMLKhM5Khjm
NeUAQGyriQlaO5ab5QdH6QroEB+LNoMaN4EvMs5dujGK/0mZCfNcNBrE2Zw8TK5XgMdxckufnPD9
nS62ajc+Se6UYQD6XMAUWaFqE7aSHJ/RpVFWOexdbrgL760Ty6so97Uncvy3WXBJ4Lc5NOWzMMC3
0/jA0ZzHgjkbb7voaKQAnpL8u/UJ3npxug+g16Lm7kzxwXbbUVJ1OxNisRqZZAUp4TIv1u2rBPFo
p3f1KtUCcD8bWE4evrPdKNBOT2CNGKQzm5YgAvoOFUG0plwZz0ADXKgYe4CY33RudTGxZbZvPhDY
y70Vxn4YaaUft4tGO7qBq4ptciw6Me0LNCpH6/M1TNXZWGbEEEpeSa47wepQUCRxUFYqxPqLcMdh
0R1TbP43IjC5wtLk59heY0IlpWOx48zjMtjOB113ISe+Oz+Pb0C8C8qXGuh0Dywbiqm8ngkcWvtx
WrMZ1m4mCr09nDxfYdUThwanPhlx9MirUevtMWotVNG+d4a6/sGTINSWN6ttj2kvrLQiuv/Td1Gt
Q4A91zPquni3cNj+IzmLKGONgQD+XsKbnhoRmfaxu1V9nAuC8rPwPcgz6EA8z85/l6Y6VWdyw0yQ
VdXUS41cXUnthh1NGIeJlSMljSc+uMT9HgUCl3Zam/sljSbk+5nvDboidbq1IBSGWzhSGvPacC9z
3mnXXGrTU17dGpGj+PH3GO3Ng32/8cg0C3SGguS94+t4IbKG1RFfREHjWEKtW8TVhH2f6UTs8hAM
/Cw+vxEV565YJqtsl0HP7yVsQCQl5moTm5nUvBhHLXmAgj46Q+z9nYDXwAmTdO896CtzzGAagpyC
lAyRXa+DGUe1TJWuov5N+e/X/fpILE5wAxbB/rsHXQilXxTg8rtNxcmt74WvST0LHFVbTMoARaEn
nl5iIUKODbuNNdx4qnIRjxrJnx5nRT5qysVO/SDRvITGh9372Sk/Mhh59CWY+GwPR1qE2/cBtAzL
KqUpp27aobZRf4r6qn/tmOVCJrUAWcQkZkeV+7QhODxobtlqIxrbdJX8J+Z3xg8gpCLyoYfRIvLU
aA4QZF2d6tcuGilwLByAjziSYFZivTiIynLDgLbuG8p+jmW2/kWJzwRzDHhnnxVhJguB0/qUpHjp
XUzqaiCiLqb7TZMGNodfZa+L6dJrwVuha74/l5J9vzp91GNK3Uxut4ugxWHIVhKT15yn3X4ZvrF3
05q2icUshc2NUO5A8a7iJ8ZQ1UnwiFO935o9G9KJmzKODRSK2+zChA+HEzpa00k2Y8z4y/SMa0ZC
ozKoJo9c37UlKlFrtRwV8eeyOTO9l7sXuI5Q/2mhoPebp6J0xil0gN928cuMLFuqBbbPQYX3FZmP
y2u+lOoZaKahTKIhnvWtNo8XU6VOH1li2HvKk9gCd3mX1E+MKlXtnD2BdOiDXo2TtHMuhjdK/V41
DFrIfjokmN2XzlCzgvXvUOiDmhMyJcG6OWgLXo1TiZDSCfdWLMIvKvmmvLUFgrnomzIpI33tDYse
7ec/H5EBz3Jeh4MG3LzpiWGX4FXzwbIW7khG6urm5apj5yOm5QRDqx6lxeTyiyiMF+jGCMjASFf9
auyST9q/4j4qXQ5NRFEW0uSZRwIvPh1RchgRvNxfxKlXxfFIaC7d/8RDim//bfbTCEYzTJYdGyR8
/toQpbfC45i8Nb6cPV2eu7FFraPS36snNk4kQh3bQAoU8ht+cN/QmnvX6IQMPen8tUX9KyDo1O1M
Q1Aim7qJ83txDP5AbUkEvd9ctSdoY8Bm9TenQtIOaIGqZYKWA7S5K4IOClBzUlqu/GgomiirWyLS
bdEnP/dNEDVGIII4X4EP3KlGXMg9Qv/NmsKOPhHCdhId1mjW3ZLqFJHCrPKZScIrOo83NIHouNPP
UYxASyuHX/mrsfiJC9FBO30qJ6cBLUOZcOhbgCxUFjsB+43quVwWq4n7X4e6HE810+rnB65d4BvL
rO/VUBZXIMhm/t1SE3ms9purP4PCDHECWM3ZPXjwkGKXJPkySdLwTJeUtqp8PkcqqsDi6RmoVGnr
fMTbmVc8j51mfy3ZGCjh1WebrdPQsaQTkT0oZhFLKZjIwGMLyA37UvoiCOF34N/Rs3xg3NU9Q05L
AN0fE9MfMuzTwdjRxN1WnVz59XHwf7e6jyuxwkT17XjAL9c8qAKYiu8Y56QWDko0VGUCsMheUxPV
k2PxIRFHvNHniB1CVBazXOtfi6lp8jbrgD4TTCUVOR2HsvSUczqjKXqbPpl/hXaZzbKgqLDl/uOx
o54C2WMfvAftiSRfp41WBLnIQkSNSiR0vR20l+/KayRiMR4FqmO3VpZNX1vB6MOpr2gB2gZCTniL
nbqJRWsICMycZRBAvP8fBdBVpzFIZVuK+XXuO7JCtPN93AfyI38w2jD8YP+aOFWzT999IHgkDypg
v/7DqjVx2XTnKuuBtSWjpvlH7riO6NEJgFHeYhXwW1syuuTyIzB3/5tBMKZWNBdDOwaGfA2LPUvS
UAKG5PVmBx5zQfp0Dv3O2tJTMcJfVpP4pUHu/2kcXb8pD6lxjYf609LZgETAjAY1ZuUb5nJnlOkW
gvjpw4jW5ih2yHWzyHaca2DpJbpnjIWTsKHKbsTd64zjInmX/y2dlPtlOHVWvr0IeZq76Lu9vuQ8
f4bnvNTxGpb+LU7jx6ET9CYGp0v1Q4kCU2wakqi3nRCxPE0+Xsjbh7lEnydqwLvM6DxCqTW+oMFP
q856AdW1zo1GT6FRi/KCAAI55Muy60iYWqtwb/pIqvV79PRvs6p7DKJf10ANVc8NLt2AxSiX9GXy
qgodkAV2qzqgNtNU6Sdoyv8NHy572iuwvPhChg0Y3/c4gkPZO0xQJXj+4Zu/kmV+0KRtk1iGr+Xy
4w8EqMlwVcPgXgocAdeEs038PD8IDOkuk/GrPQXsNp7IkkiTlBqUJ4H+1BnBu4vS3YvvKausOxz/
2qK8eOfifGSdNT6PnLS8UGEkG9hwf6yUMgkOL6r/mVd9y5OYFX1J4/qsjwdGmi3g9JxvSQvYnC6x
vv9Rc/efv91e25qjVDQbk4TkVB5V4uPpelz8x3C7KWZQDgGNulXcjb/xhI4DV6iL/nS+z6lAVmX7
BVRSorkYLonunvTDmdA1HNgkUTXTjhy3OpooL/rlavHFg7N7K2CKHQVD/DcjiBIJrzVrKWXhSmk2
eY9hKXcj7tkLZfh40f42hZ8+mgfZpKti6pbe/UKdmLX6umf/ZqbB0P6GUU6u1smdfNiNshZcRaGX
7XtELuVD2TWShIa7kmmqZp1II4EouW/byvKcfJznoifBQ5rXHwA0i1eF/iDsf2RexxHVADPUIpiG
ZpEbekUarqQcxOGifd9EunEt3KsGEYDyqi32Kj+TwqCg6/GeX3IT3SnVUby31Q9w3Oj0GzEcT4a2
MZBetDkPshPZWX/fCeBfpc3LP9jPD0yd5Uetd+IV8lm/qe4APyBOPtEbthvgaECKMq9CpsSps/IC
Ra+x2Ehsn2bdJNZBFGgprfgeOofqR/iRkemf4fp6DTuQWyDdiHnumwpmDSMCIOl+SRkuQZDLNR5K
5vGljwxITcQFv8qoVEw/18aibFmLMtT8PIr2XvygpWCVyG4X2OwB5424dGbcsZOFOr/nYhe+FUL/
YQBPHP9QP1mS4v0mMfXbxKXW+H/6qgtbFUEXQwlSw5rSd2DStolVtLdyC3ck6KofUWJ1Er+hrmu6
cNBrQweCovaRbLZTaJu74imLASiAqSKOWck0qjIDMF2ujhMfZLDTmv8GMdCrLqzfvHXbmN2OJubG
jjj/0vMhRgif10mMJek+Q3d+qDoPw5vOCdfWhzmZQoc0yrBvvRn8aQasrPxsHWrCG76dCux1xE4a
CUydjxlV20KIK7HkyPKFvmVWW3WtR/MTpV7VbXKe3cUWbG48089GDIEw2ZHG510KKXEMPVZ8HqIf
N5QA5JlmKdxzKyUhV9cvJbgknpnXSc+qzzH9ix3IDrUweHh2KjV5HT+JCqFED3yJJxsWxVR+8Lhm
y5R5EQ2naPfay+eJslIru1/qjifOEIfXWxIiqt48tLLG7C4s2ITcvjq/QP6n/7V+TulhzemGwyqt
AMVBY9mpagrso9Jol3K8GNPQuD654f9/naphnds4cybFaVI02bepVq1vZ/ktFoP77syrfq5EhXL/
ATMcYO0cUHy4FmADn1xqWoL3AMhgLyF0OcrzNP5RG7DLDRD70YJqA9Jzm07L0QW7YNL46ce5VkSy
9jiqh5gJSj843+/bfkKy39gU19tueX/Y5eO9UX4w1FJyKTr8keFjRagmqN3U2zq+VHz0zZ4IvRX+
S2+2Nx9H4Ee69V86CV4RUVqIDjVBgkoNsMBuR9nuSZmhri02TzYC/cI5K5fl4R0h0AyK5Slsd+1B
7/18apuRFG9VHxlYxk/vKgy62s1u+FtxtjLq+e5JLOKTTpRdBYyds3dKewVX9Tunbq1yOZfZIfui
gcngNWvQ8NsARUIiFzj+ZuPBO+oZEN/kBjMkxbKaM26BhSbBpfS1ZdQSUZrRPW7EHwvXN5HtKgKU
3eBqhsoR8zpWSFTW2gbQrTXx0bjO/eFoPOmnkXtN4ngSy+ZE+hzOuooUDMjzMpNxLLDtpoFHv6sd
3dOhTBWM2DrSainsTMgc6gmS3kN8Pml/8FVzOLV6mLj/fIIZWaxRy8e7HKrUsL4NA2P1YT9yOOwv
I1EhP+fOjYpZLAyl8tz34I4AdECW/orT0bgbWcS9RBBVBh39ly/3/PIWUFfkCjC0gs9HtSKbQ+4e
X2wunc+Z1WtuLVKn8W74qAXgg4ffY0frDCw7Ty9A7t3hlM2lj/8lUxddr166LGvhkMapaEz6sU5t
I+D1WLLjHIJvrGY+canFzVd6IZSpaN69tCf58duHqZAnAfvV/vkA0Bn9soQUB0gW1ykDbrGqig2H
R/79c2z3kx5fcUJ1dSsKXtad/47HBA6BXZ+o8tZC9nXF3GJ8ubgHAaAWcLHaSr2eEU+VzyFGnHIn
FtbuvX/w2ibGo6oaOqtx5AL+BXEpVc3BhdDLLT0rP3hFeefCWj78gqTucynkjpi+T6sVkKY23Bty
68hF7toMZE/eB8At462Tdi7CqozzcmXzvt6CT+gdJ5i/+erjDuqFQF/z1kKHKW8KJZE3x//5VGnN
A7B5m4BSC3z96UVE2mSAx6/G5Bt+HVMdr5DsyCJ+BZZvS05rwUYnvWicFeUihwlq8uBl5094mIhv
0DtpD/xkhs+ZAny6h/nJbb4bZ9rJGLNzRNp+B9GWS25lO08nEwwimXyCduWe/gcLsuO20xR0yhhi
5H6IwDSBKUQJ7X3W6q5/DmeXVfXwsSF2kdjY5q0SKYlJyCUQtOGximAQasyxoRGWo2yiVPsRU3o/
UOKnXribhjCjKE/DkbYT0EEwLypjJg0W/AlNL4AjPpR8VlvQrQqSIRC6B+V4mYqLooi2UBg7gyAu
cGAult1J6yZWVH04Z5bcg3VvVbwfqTijsu32cg/AKT5H6ZxFe8dzH25edhSUp4wItYdC7mGnOhBx
s7LiP55ekSS6t8PPtdkoO5QiG42gXd2yisFdbEg8ZA+O2VMBZ//fpqb7aXZGBOyj5hoF28pY2cbK
KrCw8rf0e65FsNbuPiOrIHfu7DMfzxp7H9wzptqp1Z7HSvhPc0YIkDWSPogY7Foo82GLHmZWBUnA
ItnFzhrAnDwpblFxvmNpTieTxa1KFPPFuXUEuW5/wXmWZOeGNPvqzEnAT3scMgmx4IqbL7a8tOEa
DWOlCOuq1MCN/J8U7754KN///fGGmgJsg673Ic0VMfMgVLSZdLVSOmeos+c7csgwA8sBm2Ax+J5X
MDQqNUBB5nvDz2JYIKPht5jZstqHWSq3RwNSP9pD0Aiz23ErdGiUA75xde9WbdQcGcXFM1xnEWta
xQ+9uc9bWhphG9mtF3GKSGM6lgAiC/rjAVp89ianzO8uLeZaBT8oUBvdsnG5VBiGiVAf7Lkvrivv
vl054TmhOEOeMct+htMEESzLpT1OF8mVFPFvIa0tPr7GHCljonkOenAVtyNNWqBwP6ZabrrrH7Tn
0uQa14/nY+bMywfn4PRjan4AMCpugdVXb8Ou/SONC9c8gXCjUyRe/J3dmJyweaTxRoOSWlLt3zDG
i4WkLopt9g1XsP+AJxTVGHjg21hwY37TJiqohZx//4meRhWbZqq6Yjk4jGhpSAh2j0aVnVxa//0I
qRGbMxwY3LlR/kXibJrxidSDx/gVr3HhuzH8XHM8h6x1YetpN9n4+BeUAswnNQOHyI5HhF/5ukCe
ljYmSYuH4UkWEeRgpNpPYK78UMR23DvXGtfwtK2z/3KyGcdMsEM69Zq0NjZ/wJUcHTLmncnQMqSJ
x3rhqnLQ20vUBwd7exM5MSlNoHjp9XXEnWf0tbs80CjW1jPy55FmfxhkUgrUre0MBxC2GctbhAkr
wj1YStMxLQLrxsoAjVGM9xs6CFDPjAeXYeG1q3uqAQdmI2u4FrL15ZnF+rk3NHUVspFPYNj9oQx9
7vOrV+TBXLnClAh5oLdJjeEh8vTGttL1d1rQoInOShqOe0aKjXfAb5lpA75WtdmSlSJ5vJh1I+1u
mTVSkqOI7BoIiOu7/Ofoypf3TFg3M3KCC56K/ynlkxF/173CxNuTKYelqfondcP8ishFs2uYs4I+
P6D9lovkjigQq9BhUcgYRJx+u2FvITJfQ6JE9XxeevEfaSyTFmvEaF43gubdzoPNVkQwD2ZapZZ/
J4amrm6qkxzUkDcFrGrHWBCMb8a34LF90KuZ7LtD/b48tIKuIsA8lhW8v8H/CA0Wau9FoSirfasX
W8rYCZELB8E4Sl5gpnaISxm41iu3clX6YS20VeGntcjBPW4ToWx31q9QPcDb4Jbgp1AR2/y5OsPc
HH/ByCPtpKWk2e+Va1ZKGvD6MZ9229moEgWfPa6dU+Ffu26DrpqtpCWg/MYgnqE5ZuZa950jQlUL
GXMmfjh8QGEAGLaZu3OEyBotsmcUdrqf3VepHnBoJ1KM9SFU1bcKLC4cX3c6wrOpwcz6mAfbt+1x
SW7jIc8AZUr56afblQY+6HmP3OFq2J0ffscMcBae/Ig74xr8XWPj9lNjto9RmHgPLj2PEzjjGMwJ
3BOYURs8brrK88VedEvvDqy7cULVkWS7eB6ViobIVnPLyC+xvxNMgScFm3GgZucRB8qkMK1hzPbI
+zu1RGkZNZh6XDJKFb0c6deSjowyAG2YFC3pbOjYb7S0AWLW/wpjuQ8vKGWf2der9ohBvQA5bCrj
1jSGjvhoAtIryD4KMh2vhdTRN0Zl5YuqGWV64SD7pcKjQ321w4NXmrdeWKeOI3CUW8pYW3CkG6RS
MS8+KKMa3IcdXtmhXqdLAZNpvLMZIAgMRYbvHXXo+qW5fbs5MkwzzY+RNwZMO/wHHa7jY1KwpXAQ
Hl3u9rDB1p6tI1nbuDxZ+eszLR9o9aRDtqFs5Z4DoSZbE78UM+8ncXFusz+GOCCI8ltu4tZlt+oE
LFrOclwXH6VktBmQJLxqYvXgqNW8B0yPQ021Mc8So/yoJcu3U+fkl6nLdI10PVKfBH3itedcf0dY
XL3FJD6Yc7NPqemf2+DTw2s6INW2pTd4QtTchNzBFsUX2TEOhUyuDJfDMpZBXcrLZ2NvUN93bKxb
bfowitYt1Jb9fg3bM6LN5QGWmR0JPxffVBrgGFoGc16R31wWhISifXPzreHxtSQpFb7vW948v1pO
MQx0NXa0Ad9fClt3oXUBCkAy34ykutN2UT5BpNexeQ/HmWiVnjRzuEjI06mmoNuoGvJ3yM77xxxR
wK7H0TFGEKrAjRddxF5wLxrGDByD2uDLdQNLd2SgIu0VU1CZ7yixn21Fx4bs4GLGKCcvN4WLChw6
FgrGgmI7ktS0eiTjH6bNiVBRvuzVnRKhBJA8lEsV2vJoDf3ArNa1sV6hJ+vua6z1493ALXqJWTzQ
1e+sjjl7645Qg5De0f9654UDhA3YoPQJLSa5LV/2/54YQJ8Hss8CZaqNJZaRfXOiNeiAJ7WLFzmf
5VEkgKCx+yduWa031pBXT3jbZd1V0mc4Y09016jn+y+WdVFHPf80nSeB9qfIVnaDPYUpYN+GdV3/
hdNzENp53I3kGDfbTjaFMmBOsi7mjB1ix6EHW9/KgqHmeEMfrHs8eDjAZPLChEA/48RlRZl1H73u
5dmeuiZbYZnz7RRXATnFtzybaM8RSkL+unOb9l1z41uIr1bD3rK7/ygIZyIhNZSU0YfEsT0Bssse
jZmLcll89vh7l4dU8JboWMBGFebmog5Ekj/bPSk18fPY9c60ahAEWMWpt+xhRRR4zydP4AeNtnNg
eXJOKWnj5PS9JR7UW0Aqihog090ctOIENr78+KYr2gLzVU6+h3dyGZ/k1B4QM5eWJRFIFA8E9RRn
3+G/gRQKBQ6aY7zBL2pZnmFFCFQvbqSkc+3NYwg9FghhYb2N7hgz/ApdIIbwz5y2T25WLLaM2qPP
9SJEDNzqUX4IcE6E/V6hnia2ZZLIoyhZ5mjjZwUys9KlY3K1hsRl+4pV3ztyZgJuA/WZyFgS6x3/
SSOfQz/41A8bDIGYLW8Xc9DZ8OcK16uF8OxgfVTn5tjY7eajkSo8gtoZ53pELarDw04GwQ57WWdD
sVwMGwC5vU5rLL9XRf8VDJUE0/Sd4i7XHnWMj7EnsLEeBNSIX/PL3yWSzvvzC9G7fN3YIpY0p+tL
78RYlEuVqsUsH/6WBFO+GD0fDmVNVIA1UFdtKn9FFrtNJ7VYaEFB+OJq5zzkznQJFx2oGUTQNQaP
JnI/rq3Pu3Y0soUsVw6X6qb9YCyDl5LX13roFjXxMW2AO+icwgSG3VuQTCAbGb5ZvRvJ5bHqK44i
ZWYKrr8kPprP6qGtdN7e0fS9RtqVrzRw9W6swGJeImNOGdWi7Yajge9LyU9sKScBWlNS8pC4I/iS
Tg26RXrO/10TB098GVKibrY6OFEXnYnY01ruwffz9JMs+1aeLPU+uiZnz+jEvLkkJia1Jzb+IpRR
FxR7p4CKaq8HM3heMsuUC+gMvnrUwJDRTEMDc/QR+17IzXn7VrU3UGlZiYDPAjlj9xJERexi9SH6
kjV9mAG9wWpH0k4pdg7YponarYhV3f9npYnyI+CcUBM/iu4I+UGyqk5GS6bD+PpKzb/OImZJNinS
kvlbPIPbKTKKxuRmJCH01h+JqcN6i/uh1TJb0vT2LEMFmU+k0e56WiukwBFJsX8cwUYvwMON4B2r
4FVlNfRZfqSqmaynPnv/d4UTffi3ZSbYmtka5GYaYl8tpe6poAaqpBqlPtR2Do2+MePwHotByY16
TjWUbNXOEOXUjlIQCGAEHlLfQv+DIHKZ7LXV8TLe2g7kDQEeNEZiN+CP+cjud86ZzLXJMufLg+ek
vIP14BeuZLeUuskryc2KaeEYQoQrIynTApGIzRtaGXQUGA+UmXD4ZQW3g/DEjAdBezkHgU5CCiNo
m1AaHAwFbQsWVTgQUZHSRfsbP2uZj8/Hh9KfiYD9HcppUdPpjV7gSuPpyK4pyN+govk3a+azpplY
yXmtvT/VtCNE2Y7Wsw9y4SY6ZE05rGOwOBczP3S2u5POzVdbSXx/ZUGiwkNpgRhxl5IHpk3sAEQj
kc10Auw30pQBsK9+DuDYo7njuPVdHW5dSZfPs2jV+dFtqPcWQ23ixidUgus93IyoFagjfquZClPU
cT5mPsDgMNlmo45JDecQs0sh8bsNUGq0Mgz9rJQQG8khGhoLdUmw/PS106oXekge9QHgLP/snbQw
n9k23LPEMmXGdJ0hdDcPbHo6+zJ4vaj3Rn4E4+s4us9ksjiVizMmTR/VZ/Ll3vbnOnSFBk/EPwIy
36ZNZXaa0dSjfrSob2TVuJW40n57fTTQ2t4e5ZW3454s8QjAtrHGZa0D2TOVOpHhIgCvRC75i/a8
eC9DgNivaRTZEUhQLvydLagvipo7C5XUk/HpSiFpjN7SHuHKNO//yEwOxXcrhd0B2GdSQ91UwAgL
FQEkrZdFgY9UXteBI5TmQ8n5U/IVoW+OkOA08m0IPUaqKtRndLlJZ0zeZBFU+TaGRJxhKzWcoZen
IYgA7CEAUZMkEaN0SKdnEQaem27gYtcav21s5jPI/yPf4XS1kzhYvNRGIqCSpWoCOAf0+lVnVOor
FNGuSGRxN9PIbqIV0hNkB/WVCpFJ7cMXG4Zs8xvf2W5alWwSH77ws865C7zE51RoChl2CKMsd41x
mHsmtgvOB8mCfRYMoJHbcbMWOfu4NbLnYBatIYxHM7DniuJPpxCrfjbMhdVOnPIZwYUCkD9bOQic
B4qkH4To+n8+Bw40OhNsym/lR7omhWfpHjlq8EhYYpPn9/QUaQcwAUZyhEKTHVQL2HSXsee5dd1i
yvwWEmZP/lNQF7wH4+ROYctgKsMNQ7GFwZ6fh9v1B/Zpawhq6qbl50ss6/WTJtvoX94CH3pAQF4r
EuW6xGCDkU1CjgsYoOaEcYxVQlqpb+heXWAjgMP7KClscLeYPsPDXdYc+B2Bo2WsmXH6kpQKQp/y
15wQDeKuhs5BWOSH0QZPt6DBH7z2atPyCz7IVf82dfsmQP0oIofgxupi5VDQkC9XksSEnzJL0Rud
E64Hz8ovLIFA7k4JNl8AlZypVlvXGbjcTFV5Q0QiYhTGR/BRdAVMjDxBfgHl8Ht7dtDkzJ3VO578
O7szNOr8rqu4LDzmP8EwajmBU7nbfRX6pjI14hUGDZLYNUPhfRXT+YXq+HXvotpT1bBTJ0o8E+jI
edxMBT/IHHk6+tMJFxYcfWW1U5P0fU1jEuRYChEVV/QEx7a0QNMSFKvfkqmBf0LIylDwzhBigXez
JRmsawhLy5Q/wVygqXfr5ZeA0EtPOAemPcbgeuCbEbcAheYek4wI/WHZmP5Z4amc7WutmLy7s5KV
6RJhHFx7Jy0EsAxey1W361e6CIONnk8dfD+ObKYHEJ8GdQzooSAmNHhsLCMnrckGRNeQVzdEMf6n
t/KmwbPYXCJyw3N27UyGy2gOCcnZ3J5ZETNaVfhpvNkwYMtmFbre/yoy5IWPOMeFT66wW6rE0Al2
KB079CoxxKJ2RwvGblqJBvrBtKtm/6F7Xgmd3UM2XmxWAndEO+SwsooHJwkBXRRxdB94O9JBi6U9
hLe6urhX6vGhPev4PAA55n/AKP+04/uwViIfjFImBZ3v7+5d/3CIg/+ziEebEf/mkazjZAmxU5aP
zEE4xpeyYxRSeHxs7L4oCCF9VVa39lOmxwbRkgk8cpnJzi43UuzvaowqqABYjuWH5y5+PPhh9z1C
VTq/Q1uLhuL4PisB3R7TaQQFVf06g2gHbk4N11a9UXBPp4eT/frrH9yPqb2VVXLiADGvJJmbXWdl
JgGyJP8znprQitrtyJtA67C5N6E/SHHbfWwdyXH6p8Z5bKeeFxWHreyvRYnpjuk6zLVJeDH9HZT0
RDaV6CajYhQtchha3NTDAsX9SAPEJ88cHIp0Yx5a4at51jLaQMaXfUUO85zswZFkG2urJK48A0Dh
Weo+0qOJtyBehMxBx3IgGZGUOGWh1Lkq/42k5YNLFzTgi3MdTcJ1TMaXcfM79PAVM3a1ySnjsH2Y
GpMwS9BdUF83sfBFmj7W4G5uqL2aDf5D6Ib36C4XDCzBiiqXEzux9T1vEM2CGzd2AmHircgQUdKl
DjzN50JFQpq0aeLb/pJGIEcfbAl1twgg5meqrBUYoh/lLm0WniTYFuDK9hGtsGLB0s9IxiVRW0X+
GPoj19BgQF8FJV+SoWbVL2trjj1wsoI+/ubM/JTxokZHsYgklt0lU3MzBO1UhwN/myfoSBUHX02D
gIEPQH8fnpmJRQ4hVDPRJKjOTrZa0K5kxY/Jof1sa4DYczywCiH7r38OQDfWKk/5f+4dYSoREOt5
TIa+SB8y2dooj83QqQEYt6SItPmnCufxmxwt+pgpikH6d5vZrefiM+Riaf0ekE5E0DLaUfYqvlVP
BgqCGu5clgQ3+YtpEuhB4tGqQKXREGL5TeHBwojFgA19v07OUsE6JoP5QWzcdCf609NhKNXiJjgk
wBY8nW4TLQczLjtCw4yF78MTuwKRnma4go9Jo8hq1pQF+fO5tMmY3Pb59Y/wnkEe7EZ45f6xwlzl
JdIJHp1Eigvl/gYX6eLK5wH1ckIYbwZhYSwbdeUvthd8vRYF3Pxayv/rFWA7kcxkZ5+FJAY4j+Kb
qRyQcRbOo+/J3cT0W4ODkcYXY9BcdbzPVHBCSHbGF9A4cAiUxhQX/M58swc3f/50/UvSO9myl3kx
1GzBfVNHMMPdB9Y7hs+FWw0VMt7x1Mg/GPv4WCXjBj4s6Ua+pr2SxKSwyqaasjkYbVivfJCV61PR
encqi3XgVO7Ugzx5kE4jojgN2zvAYnvq+798tnhduOKk0012qf1g9Ifz20ezKLsKPR3eL40kkLBk
FiagGf1NGeSCbHIWem22nW6tYcdGgZUgGrZxk567geW87FPqXI1wfzAMXUZN+aDcSeNYjKxyeKPV
LyVlnc3zxSDwobzyl6m1GYUVMF5ZipLaIVyZSLLPZ/rLZ8O+DMRsP4ZrjFC0wVpPDggVttLs5lcV
2GFxG9R5NxmU54CfU0fvGXngUpY2GDXW5aVnec3LvFVD5jXE2lH1jJGxLM1eGCcbZj+sVpokQR/U
oY4kK9slfkhBHq+Ni++bU+DJ42pUq79nkA+mldQMKFqBFYjPL2s5H77XEdUu3HO5HZOi0A3bci94
lJnfnEpNRsLcPgUPWgMAAwEG5iIBfXuXo4Gr/WONvzuIR/+T7QcPnZ+MVLChUOLPn1IPoppplN2F
HlGrDk34loPzmV3GBReB5xO9HBiWU4rf9ooXhawgvDTSeUdln8hDgY3I3KC88jCYbFoTU8O2wtMf
FliI5xwm4NGKbcctew2QltZAqiMHbzlWVabAslbCTSEYfX0cmCHZsUs6vWv5XdReqWUk6LdyIpLj
+Rf1jKIrjGB7DEZntV2MfIickMRkgLb+sXJmSVBY+MWnnIjcLsil/NgMmF4WJzU4P5TH2LyFpTbB
lpQx6Zyl2EKXVF5tG5gfir39o7SlMZt0CG9qtk/WMMWObOKCTcyEaj51sBKSNpjtjFK6sLW87SdH
7G3NoDJfVERs03ooXZ9alVFmODNzPDZtpQ3+P1QY+aGKwfNE2zfW236VtGkQoSBvdFpLcE3Fsxrj
CHs3+JspM40dKFje8z0l/IaQLbEYv4eHsmqLQh/HZAWyr9/iM3E8k5ywdLfIK3Sk5suVRlr7av9h
zn4ZzNlymf3FhA3Lq5PoIncrX41jLSpQkAr6K2tNfvBQb3PgHdwgGX2qanojrVxgf70+41s0w68c
GwR2OxVwY/Goq8ouocYGShO30mOHCKnvgihtf6r1cO7EnBJraD3AxOV+QwD45M7OTGKJxnujkV3C
q3y1+EIAFmMPFXplD/bo9qEBLfA7ShWv8vFt5xGbvQqT7shryzXz90sa56UcrAw2TTurl2Q+TQL8
Rz8bAdLaO9FxMzO8BXv3eZ9vGmosnslIPPCJ/tSUJV2Ran0W55lsbAzj+O2GZdBojiQPYQ5FWIBB
F3dhCB0u0OLzPbgnxK1fB14mVz6KsVLoZArwEURK7Dbi3S9J+HgGpZq+g9IXuk3JuUgoXeybeqzQ
rj+6GJD7z/tFhCCbdZgXE4O/JuUVZI6Znu3VyH+9HbkrZxBzD2dqKLbEBK61f5alPadQR1mXmDZc
czLG5g4lRXyyPi1bHytuXtAspsCSJqblyJPqTMVnu1WOhtwup9DAoExcXXgwNskcCkLbqW7FrH7Q
1vB2lN4sLtqaU46GX9PjzH5NYQUOas7jhpui+fLabMb6xNrKBQ0k+y8/4g7gBzGuJuK4Ahvuq9UJ
aQ7fJxJCCgINXLoLhon3ATHcq8HKcAvUk0U4IY5f9T2qNDk/sPKe3ZRLf5N4Pvt/ziw0b4IInTSX
2Nw7R1C2rBkqebzJ6jr0o3bbNeXCcaILz8XWz5KgkiahMHJkgxvDGfIbFzain2fFIOLNYt5QcPMB
HNkS7u3XsoO6fL8TA8x9tObtwjQBjuB8Mu8IqU6MzeWRMr5MNxzk9r/48WLOV58fkKoOkXx60rmO
QIyEPsoiGgYnsi0O+22k3Q2EkjtRgl0SoycR5/NMMOTY3Lc5MqMwEUXjVqpb9dqTPZRlnu00SDPw
iNs6zE/9Uxm1FPMU1Iwolvq/ZHn01ywS7NUS0MP1ro1nJWsrhoWkPo4WOpp3H5T6vtBPEtHMmAPE
c1JTRjTKRM21W2vUh5iFBx3Gg53E/GlR52rumEOrvbutxouevWHjCwqNYhitX5ShH4pdvXgznFJA
xA6qbVFXUlLjz/6bZw+Np2DRup4dcd/4Xgu21rDTd6VCtVt5b+BNhAWrPIaW/UdA7aKMzPTbbQpD
thIMTDfFkkMuRkVZGntrQTKoGzAcWSMlvTs9BnSSM+saV++PWIdu2aHENh5rHY64AOvQQU4MPxmZ
BNdRNnJtmxSgi71rpp/NAiZBCrdYp/ihhQoVzEMeDsp/U/LBj+iyypEgEUqdnxKvp+ErD+14YkJS
eQlUUjQcWK4jBe4mWBeZVP4gXzrQOdrvaaOjheL/5XgpBj2/7+jsZP7eP0Wa9BN98gBg+rxmZVk+
5/5pIpHGCo4XN6wkImcNdO47s/sg9n9uMFRxVkamcWfMrq5pkBmnrGgJu/26Dum4mhuUodKwMvWM
gz7o5MmP7q2bewGE+lM7ASuER5IVaFltkiy4/36iGtOEJtkb7VkQgIk7QtXeC10BGCjx4wqMyct4
yw2ce0o4c0y+rD11FO6voj0i7rkmO45XseTRUhCJSV5iuIn73o51Edkt6ZzXbkUUW0HXglbx7kOT
jIC9dapiahJ3qhJYSFHGP998MdukJZI/PAe6dFm7opLV/ujwIVSKsRpH/pyFuJuZ1ds2IdDELGoH
gpT36JZgSflLvGVkazDFL9jwjvfo12J5A8qsX3lNCC0ke9518wJSAD2DgUG9aM8+01Rsmh048f+b
syUL6BLoNiFjT6t7mio1JYAFSyfKY7p2qXs85+N4PxnRUaP7wKnaPFAD/10J4YEIHPJXgzwFZAiR
dfgQIscRyxjoa1cQTMHvr59cS/DUzsrf03o9r1GqGuS4k9Iwb9OgyUGSm+a29fhIqgwWCAVuBO55
14dDnLv9rh9aeznZPWdpyFDxvLqTx63T0I6MUWtDnrr0pxnWOcJaHEg5qR1xFJp7VC5/9kHy4uoy
CI/5MlrljZ8xSj0zbbVycchA0xw9nU+yZ/aqsNGzMTekHxBgi64hCcQwxrIQtBFLk8D/hkcSJ5yR
IbHQ9ZlQ8ZCrzWNXla4xD/6ILy8EBnUHgKqHUMk5+rjBBYvmlgkhC5uA2N2tTDUkY+lSOa84q7JP
3mYG6HmzjeYAH+mxYUv+HqvkcK04j10RcDNcSaaoYBxyKx63C3VJx90lSVV8yMCkETEX7XO76laH
iq9UDhlGJz6Q2pkUFSyvMCT8XtLKedbhemnMBUGDI//1m2SqSocRXJE3WeGnMHTEEwa+DGJqiDMg
ATTLp37nHg12lu2IVazh3A1bwsocc+NhJ2/I/0M57epurCo3G2vB9Zdh6jPFuKbX3vTCUBy2PI4h
BvMk1sm0eRpu324tVROOEM1NRb3gUylwykGc9Zq5MeF1m7B68hrAnWNG4SIl4FBIbxLTuEgt1HLI
vHg4IJLP3Ug1ZUQhOWtIfuqceKqt5Tq+wyg/W3WsbdfAe/GNnDnPNa1SBtfPd17cyLz4cLEpgAPa
TGuyv8aTvWTwkxsZBviw4UwBGAoVWyVaIxOidNjRwYFxCH1Tqt31NdspCdy0ZS+Q4VZwVuHL8Qqt
JRgzveOyxxpztHMUA3JYlSjjKjH1tITn6rRbSwYUiImW1p93GfhU1UkpGXMSqyfcDGEPDPWtWrWi
s8EQ/L7CGfBflxDc7wf1PnBuCBn0I0SSQi2rOgSCE6urk45A/8Vb03CGLlNtuacvmxUIeSFb73sI
mOG4CspJ6MVxU26fhkTTurraBVEKJdnIHQPinTRZANlxweG/6LKDrKfJDOFj8Qxol/W7yLynamNg
4qvTVu4Ni13kRUfuih8CJ5DOBtMBCwe1Je7/wrEIX2J2S7VTypr10KnjSQ8BBkss9sHtpdFOIW0a
i2oQXLGBnDGLH4mqxiZQxIezq+9clwCebqxc+6fYjyGr6j3RnlMohyiNYRdAPt5tg0TnJ9m+aGXw
Q69zX9c+wd4y0HOJSnqpGpT8r2GqIy3p4Qnz5WOS/UU0rjrutOBiVeQKlmCEiYMAvzZNyHKHBf/Q
KmhvvSRBRIyYMBAwqqOCp2rXoXt8wW2+UsXvYkGwrR4z861U+PjZu7+Ye6MNGpUawBArwTjVPa5V
6pKIuTuVRH6DT1mymSxMpG9HMxbZNVCrQ51BVWBBtRIuFtv1kuEwrWwxUa2J/EjI/cndMMdRQc7O
4s8Zl/df9tsj3yNF4JSr7uhM6Qpdj+kgCZul4j96Kv+B/adtnYRE8fWfSmSix61jEKPwrsp2z/Or
kfgCY+wsgSJaNe0mvWSVY95b22WL2OKCObNvl5iiB4k2ptMwejm1M5k4yPaC3LFurYRsZzNZY3j4
sCCTMjrPe9QsZrMw6MD5CgjaUJ1uRODS0+i8KxEoAbeWF5cCP01/xYAWBGT8hSa11TleS3S4arDc
ZnEzJMu7l7HRry1573fC4iOskev3zuGbZ3lZ5mJ1aEKzqZ/doURxErY/CXzEyPPBpMxjvU+3MT7g
EaJtGQVHQmCvdODLNoyqKNr2eA2xvBjCNVfGIY+IDbDbU2GHM97cogqc+81Dc7UTjuBuS0knwgiW
jgApl7nu9MSFoFUjHUO79H8Kh+DS0IS2Ddb7XszU/7Po1MdLTbW+jNlj0GPiz4VJ2l6BTHzFckGZ
sw4W8jUZdFhaeEOykJgcY9c6mdvU0uUvZKCt9g2gzMEheNgL1H8HbaSRWEO1VqBwwJRsxYkTrQY0
A/NauurM/G0WzNZErTM+U5y+RHnceOQLS9evsDSJX2uMCon48BOliB5UjVmwYAw/wJK9bjKNHteK
Lke0TedQa4TZ28UsLFUwO0TKtJWHhf7yB1ZTvSEa79+wYKnqcRXLaNj8qDSPOIoPI3hYc4VJlyQm
I67dYh0NbMfydImsSi7rseUgOBE28T/DpcvGyl1EyQKAv7uipgUfb8nKffhtB1uc55bXTVdfmCtq
cFNfP1AoXvDBvCEkAGt1418wkhCLCMoAJzCUSk67Jq2c7vaLfyKFoi7+/KHcm99rRn00gpYDqz2l
qYElZjqipkltQnpq9XLApSUmLHtqo+5f5v1f3g6T1bWB1RBDu7pg8muoJjC9egxE8jvRxaX+RI1r
J/Z61CrDLIFnqQIHByJdjMIpwtRlSOngk6W4exrmd+s4o22CgjAASESY/b+g/lqhDBwWoZvk9agJ
yjCv4FzFYxmK5xVO9zk8IzEFtmngbWCPknU2NPSLwJBFiHc8l/MSoqlVJ2gUXlY8iGXaxW1f781Y
R5UWM7HMeIthRGQ1oU+DQQqP+v3XZU27jAsB+Nnvw3Ea166p6wJb2qMdkte1s9j9OGXWfOALgWaA
NaJGa6w/6GyKHZIWGoMoTOJfm9EAWnBpXrZ0SFkiIHzogcf4LiHzbAgLvwwzb8R10xr2KRhrCHef
WKRyA4GxDoqgzTqoawunq75rEIp0PNv8+AmyNRyD4Eimsgyor7gj8T5gNs0ObZS6GtV4Sjuhl6mR
XMOzNuVgU6rodYhKN9ogf0veSBzbBIyuINTPrj6UxoraqmJDIlnv3yYxuuU5bXvU0IWc0Le+MHth
nAMu5/TXSVIiBRLKhZ7WZVsOX41Gjj0X86WUFk+80qJmDXCSbIeQ9XqGJGPSY2aTUZewa2nnNmzU
xDdM1tkoLzm9G04W/BGBaxZTtTqQrPAv+Ghp/Cdx1ZODagEEBjPFI6vx3zid0vIeZ0OeUQvmrCbM
Oz5z3H4HYZurtro3nLprQkWCng7+0ZQLC+8TyvSgbnV9bf0RH/s1VFrUyIHsDl+arh/0vXQqgK9R
uhc5Y4AAfB6VrZvYgxSp7L0zi3zQTu8PT0mx6pCP4DTx+sXiaEPxoyuOA923X4yPSZvwUPoIPIQH
2/XdKqn59rqqVbeDsWowtIbm1BaU9tg1Nha4as6ZbeNJz0VtplN/qrTVrSfQLR71i73iF4EHHW+m
1i0mh+e++/cs42aKI2RjGvufRt1PkQwLm7AGhtZ4OVuzqGVzR4pu2vCfZ1bmC6HaPmZQUEzt7kqT
rtu29+roNe/o4v3VHGqkTbRk9ZOTzm/VTadTqPVTQLKJmqJQ786s/LPY5MdW75ujvhYSvx66cYQK
8zaIObFKxnGyifuuBZPaWEGi+l+7tMBPWWSxFWI53B7gP5s0+XZNhonxtM21nR28CegTD0ZWWmpZ
NEiok3jBC3ypzAcUDCZ7L1oHFVlTrcKb1az0UURrEabiS5hFYI0OKaFbBWzi+sJ3bTXDrcEhaK+K
78PEuUWC9n2dXUqSplbt6srPpQ4xyQj0Dlj0bs/CF3B9PecYqZs1wipU+JMyVjoBEh3caSKnYQvS
KIbOByIwDfmsZMAUKLlJk31fXiY9f0l9GKOAUT94qy114ym3rzKpRNW3vxGgDE/4P+gE9rDjXk3Z
OlI/3KgVMhsLGxdoRToWJqrLUKBJ4XQ9PREe829wnSA+r//+wxU0HHa6np2IeG32qxJTLbmi00Th
QsJTYYR2G7nOW0y2g4KCsPGofqcN4vyNOjvvNRapT8+B20g09mSVREq4uvgCR5dqtu/Qe7IepR9K
eFmx3f0vy40XIwnhTqa0LsgJcp17VJ1vrlnalIzcLWixsnyW0B0ryHN4GxkBK0alu/XNrT8xKZV+
jxmlfkdW8rFY8ZXtpgqb/j2vCwIvaBHs8K0uKAvP41lOouIH+wf2P+ovZG6QnZCMdGtYf6i2YEdv
TjFQDsYKJ60tS2ev6s3HHtAst39igoBGQx+HDLpnEf8aWYwi4dYpwHjSpdJwT+nQCMEquQnTnf1G
gWnm6NOB2FDd8HYntApKXFJh3J49S1w6k3b6fKNhgBu2OQd06ywmY00GtVZx80vnMKgN9B8Yj5ok
Lk70+gSyqne+HobL9SopzS2YmZk8WM4+aG4mHdl5T3/JpfO5IX6K+oWDWCYFkjPKRgaJuyqrJaL9
Ac/7oDQuRZRE3kVfJgEj+//dmx0bqycL/XDqwdT4VFv32XbQfl9c11Bkgr167K8bkzZPFeV7WO2U
erPQGBF1fOfhsl54/LJPvSXZaqlMoUFJXfta1VE0R/Sub3oA02itV8sQYztUPMTBzmvcRb/0UaHX
v9+UwmWnidiGaKz/+tSlSpzVxUC6fjGx+kOYIn7C59lcHjPtS5nuoRiqijnKlIPQzkB8ILn2fIYB
to0BYWzv+xOYQ6ZF5BdwcEZM3cOMw06aTI8ahEfP1h1v1LlFTscchQ5ZBCfbnBYsno39ImH0GVuA
flR8cpd5xZD9UHE8vCsSB489kYTmI2ndYIwwdsSAuLlj7I+sY8WBmfBfJKj5ao2FHWzYzBV/5xb7
NOz99j2zZbV6Md6w1z6eXp1NuR6hswU0716yxGQO/LcrYnmVscYC8hTES1wiCRn2Alv0DRvaJmrn
0ES8M5XabJR63nn/DObl66dNZ5bkdGpZHGZjEiwuu9gunlmVK0zXJ2YsGbMH+BMTElUyBdWTvEly
0lo6cSmhnfMFqBMO82L6aOvfSBVEFBzmxbo1s1z75PHYbZowOp473hR8g6PZNj5ETuttsrsJV0bl
MZ2gGM1kgwxOK65W4HdahnMa8ZrOrmVJj+ALf+IyM2emrM/kf3vC6EikDL0UoxYJDnugeYG6Lz+K
bGL7IMi4VIypeqnGyIV30ScIP/pwQu+GUwhj48nz/ELKQxZh+xj2pEq//BjMKt7t7Hbrk1+8ppvz
MW4GkxO+QXwkD6aaJ9TdSlHrHV0XbJN0atvs+w1eVWjMa34OUeQKPFSxAwpEWmN8B2oCLhoFaz5Z
zGFV3bW+ozDx0023rpuFMD17JQBdds57JhVF/F3dl8A3elLz49rWtzBRem8jHpTtUOMkIow+AZ4G
DTFxf1vjPB0Pk7A01zQQBhrSzMqAVmin/DKW2kwn8yYr59CjiPcoHNdS7DH2aX3nAJfN0ZTY4D5O
lpPm/uzjgRb+GCnI6QWXtndCGxbwT5mMxIMqRAEBhsg3x0+zN1faR/tMgbWnmcpa5Dpj8oMpvm/I
Q76uNaUcrijEU8tuwfzF/4tzCmHqRQ9wG+RofYgdhDghKs3rZoiozuFwTzIbB5NhdI3XxA6HQy3W
u/wzlPppn8XwTZcB26RGAv2gZb9ZOHxivVVmMJNifQyNpl0RjDN1Ea6gUm5SmhngE4qukLGPzI7V
bt7MN5E1AF2M6f4z3HyWhUv+sc/fQ31RIbcpsjNdmsWsi8v1UwqoP7rGcVCZRUll0OPh9DbExlje
rK1PNhAbnzJEMh7fAXD7/n8KlngHb/6EVaY9ldtJDrav/8z0KLMDrZGF0MbL1aI1OYthnL0o+xtS
tSXYUR6CR4lfRE4bDBrO0w7vOLFSZG3cr1y9W/icBL/8vCs2Q8/iB89YwJCIDU3K/LLeo8zrwg+j
VUqdOOefAJxPWcLC8bb2HCQ2mDfZmG82V90eg8GbLVbOqpuJiWIQVmp1M+ukACkAYS/MroSRKMuq
3Ycw9JnVAb8Z9fP76UWH4tKl2206U7VzKvG7aKn0LVmQ1mL5s/JguQVZDztiiryN8NarzQiyR0oJ
+ZwsMUHFw/EWpUvvn9StjMJHoNmIFMded/fHb/tSA83pmI2U430VQPArtz6Gj1vJbz9xE5URLMG1
B63fJtKMb+FGDw0l4wqwN2OrKmY8mjgl1tDANTnKRFnD9K2dnKPNUi3w/7H5emZ4Ego7ghsPCBho
2ykfv1MNqLwnGyTxgoru1V4kjYgnmqxEaI3XpkoV/U/xIhbx8XZIYIzBw+Z51g6i/Y6Lw259HHwx
GXYYP1Mpq9LPjjp6C94eAU6dkPH1OkCAfockT4rRqKJTUrcjSXyE0Wu4ZhCa5in7Z9HbEsrjPESf
vxJmJTIeqYWKNxgdkYohjwto0mpsz28tDJGH0XyMa0249NovqkiVz3KI4HiNOz83zMUbYH8HnsNB
ZQRtYrGjoYLflXw+ZpGn5imxmET7MbLSjGc8yrxQAW5xvxE5qu5Z0a5GTEFLeFSK7u/D72qKPpOf
0pDSSCbzmo7+26uo/aMT9TrNS6GhBQBltCTm6F/hnbf0rZexlwECbakdRyszlm1CDKvdmDmtnaQd
oz7P5F5SrgVFCjMpzGaYPTidx5rLsRMj27g/QaRc5EHxoNUMNWrwyv2vFwI3XtKtIt3I2UZ0fLPk
+Ch0X2yxWgXU7UZ9ImLDsRYBvjnx9daFsLPYJ4KPf5JrTqH8bGDMK5OvaDNmnN5UZUhCUn7Xq2QL
h5T4eRFKUV/NEm1MO2TMhWl5ya2N9Y798HokbYdu9Q93XBr28UMNtjw+btvB76N7Vku+dtGVJEEq
rwlinuFR08TrJ4N1T9pWvPXuEkx6Vw9dl81sf8fAiziT+w0pbFwbVWz0Yag1x9gZW0MIoqebjkt6
3iuV+c12E+E31D+Z2kqavckLj86zzmwP+IRuecFJ9ZTx05YS/iHRVPZ9wCYMIHVnxgsdJB47gahx
oE+ruHGs9Owvrpcb+XK1Ye27MQKrWHvFnlWKdRuLYwWJLIeCazbFY7AGPsbCxhvWfj+V/uq5hhnr
BSLcW73SxyoxQcILy7nppO8DLAOCjrMmJOJ6HWUj7AJpYrA58bcMTxeqwuPC/p5+UjX0bmXgXZBw
gRpTYgKstQw2fTHbgqTPaoT2X6dAA6Zykm0wTPZIxDyaF6hMwQwDTpYuZqcFYHiwswPuscRcueS4
SHlrukggCjA7WKBuUqglX6a8MAkBvIbxeWwtNt+K/QQ9+FJLzS52E5fsGGg9F0e27s5jgAK74i1h
8q9cAO1BUTVhhc+KrXL6Tv03GIxSnrztPkL4eVaoIrwcaTVrvlal0mOGXDlnmQo/yE1eEZUQay7/
63zrkTzA7/SJ99wVUjCWD6fejWTuu+4gg1RUfvlYUGzWbPOI0RyZTC1eQaSuLgBLBAQ4ysEoZgkj
yxQP6TxbhYKUv6mm4+jNRpgKjIgecoNOKKtbWWa2chFtw7z9uYh+pppWXm7pTQ2ohHrCfg1lRnoJ
ba2gk/JaGX7ak/WerIohybPzu2QuBPzd3pRQC+G8/dRSEMGg548lQ/Qaiuy+1U6W5pUC6QDwgWe6
1udjSLcuU0v9zcAMLT5GQdPamEp2spvWlV/pBjQ2vuM4WZ8A0n6nMj8XVFJLPqzM2AQiZPTsavvA
qd+MtiIwBU2vNEHg7Omm6LA+MhbS+Ni4Kw84gsy0wcl57z0gvLbgS1UO4DFSqiQ1SWuwaXXwSQUo
X/HAWpYlyRLnn+SusvTHlmHzzqjYjMQUVtTygAe60Z3oOnXVXuCdUIZNHgncn/0UmS2o9dTyTnl1
OhOmULlbPX4SLIva9cYBJJVtQM/HxtKecmF8zq8MkXLhmQShemsldUZjw5frcVJdsfptpNmxyYKE
CgIHOBdRaY6OEbIy3j8TDxsx4t/BxIS13k5pS7G2dSizEw/jxDBOoI4zJU4FVATfnNSe44ZGICDp
cTDhcbJTbx9Lgar7cWsrTEFTO4L8JcSrLn6/UOybDpvWJzwKFwp6Bfmve9PG8PTkUhrN4Y/VtVhG
H7B6UASLOuTaZbHxHreKuFjrvkeijplWfJO4eg1TQEJuKR2oLy4WxBXIF0O748oI+5zO8dE9b3JG
TPPZpMim1cM9t6Hc26C4awQDQpRNvS/236GVgasqux93APK2FSz78bXCwMPebhfzyQHpp51nPrDd
WVRfcKGiCn3EC8AuCDXAmgruRQ/oteuAks7jH0j1Sjub3Ek2k7tjgAiiOmFTLlQvbQfa+w1OupEZ
3nnB5csXcKfXkADEq+JGoUDkQj5yIgURv8EXFaQi+UtY5wq2xKxCPeuLIkpag4GNTbz0Bmo8vjs9
5Zos/iHCBGPvmU8DPfJ5ArtB8KBhtLl/MXBfHjJhVp1oVtCqKBAIkDnqNnBfIPosNsYeNJhbBZmh
JgVdEWTsT+9KZFj8zjnpSPgtXpikb1XnuiOl9yd10h7egVhzzg2qE5KuN1a6OKc4MI2jgc9yMl3C
N1+wEb5fnXja45lrgtfefOiEd3IwgqnNfyGdrIyjCDPliqrWrD/NPRQDdsU6J5dn+rzlaBHjaHme
witm/rp5VAyHQy647cWeOCbNUdlHckS1Atl+ZEH9OOsMyYUG1zlCLFnEbEpgFuXx1RaVbDCg01Ob
Y1MZSIm3GHlwF63DcLAkLs7JDuNlT6ibmlVBOAE/7rw+5i2ev+2ZbTsElxMFrOLhJ9xdgDfx2aDU
8hgDzlRSi1N+hRtemW13t/Msu8xRqDfu8O4brtCnKfXQ/rQmWp4wkeqWfci5gzTptbh/1YeWuBit
5sZUfhaQS3T3L+/UNl1ocY7/hjzzFQImadOnainlKv3lSYYS1lFUJT7ougp/OQ8NGTHvATyEbCXo
wzwoinA3EE6rXsJrPtA/yB6qV4ew+5hyQ6JBZerExWiW3ykbN8BqwvsTcW0ecZVWYpxs1k2NSNTD
zEr9eARuw0mQayvG68Ie14I/kao85T8n9H3HoZT/5WQeRrWaIH6X2br1T/E927w0vLBnZoEolxVN
okeZ1Z7ZGvWTaIFsrbozB1OASZUXWlLnzWM9X3YVc2oy7GlxYwjga0qqrAqt/CsGD2iqvRE9aDuj
UtQwVTIPe7L4Tk8kj/TKftA18IfBTjCYPC7rRFHJCE4QxaeVs3TiT6UoAgAFqzS84l5uOyJJNihv
OLoKtKP/jFJbw0rOx7Qm3IpUHBcKfqtuM8lJfPdA1w9HjhzBdmyr39ebwhLLJdzFs3MTvyHjO+am
vF4NLfAn1ss4wTj5NXELNGXhVcMZk9yNCD0YdOcSEoHlhp04RwC2Ow/xvpIxzv2QMOG2+PX8da5w
SjF9UMlRX7eJVzDXzCrnKVTslvmTSXEDHNwBFlpiUu51trgxHyu1FEOw4XvRyKZ0C+sGTVSvqOnj
n3W80LRGYzMU7tqOVyxSNtfLEb5Tk0/He6OFD0XMH9aj6qqYfEZcM+VZBTqhxkUULQWLXtF5s0PU
l/Al2gvqw5S1bPNFk7k+qlVy/GfzQElxManIv5wTTf+OjyJjDFWU5zeduPz9tzeDv4DsedcYgW0z
NoqMsNE9FCpIfty+O99a7mm+ooWaRkvoz97H3lPYFW5DS8e8kphR0b0sdEJvJZ27OfenLMbnECmv
cuOZLjJL/uUvlXxlk4SOb7qhG6WK754NlkRi6l/SjOtlGg5J7Zkah3unDRhZkte2/afxW5Y3dSd7
juf/Wbd1pVhk/sWXNRlhA6Ny904GTMAj7yCGVq0oF68Jyn3RFxmMF6RdAQW3fk0Q0Cjbl9oxZ8Z8
BUT/4z1xDsXMkJoJNDUK+8o6v72TaDm6uaeJyTwJjCayVgyXU+THZpntAKJtKVqSRUtWTCfbkxSK
iP0DUpI+TWn9Tk1DYTXA3hRaeTM3IpXYu5FVmJZVgMPIJFcEBgSuTtNsb/P6j9nGz8gzvbTL2iSg
bCR50QSTOIXXxYGojY0FCf0MeTqiac2tbTJIpam2XGn1hNddWHtD/2DXOQaTPHkSfiEkqcY4q/zo
6EvWxeE4qxGxC87uSdpmWjt8z2A8XI5u8PkD/QFdIMrRO7XvTerLLiniBIDT4Yls/Bh4u/KTjiAl
hAUJgSfYV7ejIlObnO3RKRyKKbHJ1QmOrVhjPcb5TlULEdyGEoqvVFSc3+Iazijrr0ESacoq9tS4
q29ACTRQz4otvfx4gxgCfOdmByOzvDpCz9k9sO7xyMTFRkh8rwlKw+/HJu7eQMcYCIrWSWQLciD7
z1drOEICFpm7gepHdEUaWH93aImfV1vNipv9EYAaJvGYX797TohRrVJ2JYtoXXkjFlcXNUSLvF8y
ORK8RuvCUt173g88Vxh0jGgEkhSscfj7T0Cj+fMlRlkTum7NYh9JKRxhjNXU4cZRRVIMz7bTl5mF
c7ItA47y5MCj+SmO867IDHi88AkTmzdPzfI/2/hmqDn0ILtfw1m6AnorGxNoDq8tf/tFZLn5LuBh
0iN7olWWKk5GckCHX1vz99yTy1zP6j0n7owqzvSJeOzVwOxQVXPMZeAkfX/UH+5pgMVow/Fk9+8E
acRFsc8QQdJoh3YmiC1KPWtmbj4pHidGXSsXwpqHItLp2+IGm6BaXSNOa3Z/z1Kwm7giocA+BZ46
K2LTX40RaC+PoIAUXis0iCGI8VpqsMZVt9vZ+bbjJP6TofqVlth7n2NazAp0BJzQsS4ZUcGZ5aTt
EQS0HBEeq3TFabXuQDUj8p+9qwt2g/4GmKaFqK0rBmnHQ96aSEAVDsPAunb6qWydaxQnUAhHjS11
jGi0d8Go3t3LnrDeKFDZH2vRL9tJRne9cnjU2/zJDFKNM4kYIIOFDEk9cM2tCQNEK1ybc5stJUfV
f1ZO/jfYqOg5bOKZvDh9Yjazt7N9sose61msV3uQeGlC+SWUiYbGAjA7F70EtkKDLoZLdb24N5Oo
UB76twYV9cJv9gXXTH/bPGmXxCob0Z35yc7T3ByBYQHNRUbS5SvsTzhDM/26sSE/9molzP40pKPX
uV/M8S8OagH6M1/j7ME7bVbmLDxWa3gbk2H0gnTxcDzKHDYUfbDd3pv3rt3zDYzPkAZ5LM7E861H
4F41saI/eEU2sac31lU5n+r8ghzQpUqnLAynBjmtTlWsl5xyKg+N21ffYdqX8nx1li9ezgI5naLe
TQsbY1UDvEjAZ0AJ/tIq+EQmgzDVO4YbMZivVLWyMA7BfJ/TVYguM85m1iP1odDPrUeEMy1toOih
/2k44lImL/1KFyf75XYb9NfH60j5sVRxxda2vkNLoGwlM0q9JkdMx6noHYD1ijzNsJvbp3hLj1sg
tC3UF3y2ak5WNSRD9+/0OZ7uzmg0nlUW5As2krMnU35hPxjDWvy9+ltp18d/PlVxoYQYNirohDuV
3hOupMtVmrAJLRA8Mh4iUBEbEeL1oTC+r8JTSIgsGHkJt34nU4S2ed3BGwUV6C5J2MGDpD6mziDS
jA9i0lKw79lG1ElCYO3mboSVRdlx5NYFV+DjBGbECok6taEyh/vMvUn6nHmzTx2RrFBE1BRKLwAa
swO9BJxNMjFqfxcSP8vvvMUtjQK+DVVugqN0t731PtmMJnbKXIepV5w4AwzhmgqanQty9ANQHqsB
kr6IqP6bjj9VZk7qoWKrmMYVTyrgxNuCOGDY762aEuafZ0mfeSdIEWTKkv++pwoPAdbEL+NolTaf
WBNeg7hTJLdDLacGeD+235agtR9deHLxudZ1qtHBVyREL03kjJq/etczU8KoXAW0Ca/2xAuXOypO
AccvynlpuEHMeDAOJOJQcO8ETiFyEBgJye2aaqxXBSh3qaCxtpQsQ4inBhAPA5FhAcWVNMdNlwIM
JZHawE86WKjAMBCmc0NEbx4O/uAzNaWUdTl9CCzzxMj15+u8doMEdcGhzfXO3fkPNQzgPqAFKlo9
z0btveC7h6hkZxD59UztOdpo0NMxVkP0FLs5eIeLSatTyq/HgVpqmkKYBgSvOUpELVoIerTeA38j
PH09Z/c28zKjEwWwhy96yOBmufOr3UnDYph3N8d+EuiUpSLxNyj6xudwTqWFuAaQ4wvAwLRnZsjD
Vl+jERTodr4wPE2xL2Vn2rSB/YKQ/0a9RFVdSVpY6+Xa7hCbC+dFg5mZIGc2PSbCrKzYHHvT6YpV
B5kHF79MCyS9MB3CjDRvT2ef+YxlZGLg1jv7j5jT8Bz9WRCYMf8hKJkOuaOfIgHTllO8P9RDAVC4
a6NPgAvv9SOzb6cGNreInWPBp8SZ4ilgGWd2Xeb1OpeI4cUXnngMHGXBEU3N2dKCevgXKi2OAEdJ
uI3JMv+weGdqmoImyZxpOgZz4FXfJFzwnbUcIh+YI7OyDwSwp8qblo9uH2GqUB4Ng3F5CC0gIHok
tKy91ypZ0prFMtkHtBCvd3taQONNtekkj0VzolEy6JZhbSm0XhHOD03lAQ5Eb3JW9jMyluVigZrE
le8xuQaFg9La6nT+CTfk/OmW+OrI66OoU84lQy3SKRnyjBGf2iZe87MlTJq4GY8wwstP0/YvV89C
9soJ0TNAhJfHzPflFaJZVQqlw6Ma13X4nBF4z5SqPIFH6HFueKr5g22/Mf8FR0TgP3JjKwXXSGD/
mo4Pr8rDiLwsOksVHD0QzaQeabL0HuQeTCoTUi/jEKomcaTHTnowEuNb6euy9rhJQPk9M0Q4cg36
wo2HqNdPKvWGTx8ui6oqK4SnakO2j3p2QJouKpuXGbGHICnMPGsMrECj8xWVCXraL+/3QA2PBLAA
JELSsaihqdZYTKWDnUh4cmR0E7eARVXO8D6dJ+XyCWWx0Y8dkOI+WSPe9H1V6rvZBbHgpWHGJnLO
QIqWr1j0LvcyYpC5Q3Z7nBW/+gaIPjfBI92OrJugrBjF+maUUlogRmwUvHnfI1awBogGsRHPdfh5
7LynsssKo0UmLx/CgYdBb0LTx6+g7qrqBRnmSWtfE3AvfTLjz8pWPTD0Jrc1R533GZ//Rc0sZV6h
XBSkaC50fTQqwKES5a8eAVR023ozOktMw7A/n2hOI0SnBVPDv1WC2l2ibMd2oB6x4FtT+khTnO8Q
Ue3mZeYkuAeQwskUlVVlHwY8AAqCoNyxogvZm4+D9UMFqqo3Z92GTQT2QMUpdmstb1kPac7fCdCz
rhYgGzTDWXTfJSTz4SaAaz7mrwj0koe+Eo3s8XwC0H6/IMnOkVb+0QYB2ca7hOsy0CPZbzdOT3m9
1kTg+yILUjvcSQX3T4CUdbXOTccifymW22sphdX3maHZSn4Lr83LH1bBQg+geXdki8epIYLPFBFC
TJ4rhyu5SKaRaep3boBjRO6t2tDYhqfErEsfXluiW8JPa6J1UVqA8gIoz43V9v80v7w+0fTg66bO
NAovDEKsXa53ThphHawFi6qiwYsd2xIMTusg35PffaWyu5Kk+5RZPlOtAMfUijwgq91IvOLKFp3/
dX5v+nmFbpmmrTshfZOEw+0VnHBZiWm3kgDSyPvfKaDGIv43+ItS7kkJIcXl022X/UVIk7RIBXi4
fZKUdLz64MFZbl431lDJ0MpBYKwpUCp8gDQlG0weIM01OTC7AfwCaURwFgMzfgXtEIlqoGlnE7VJ
oE33H7xa+dau43h5zHi9aOaS4sRNA//fxLAWLlID6Q1t2wTCzOHKlRI9t8RDLFzP9lXBoNRDM5FD
pqYSvoptviQ5dfcfDEut7WbR2W43ZYk1G+cqaixExSgHA6FR6pvc7VDvQ6XD2CMX7tQGuhi8NirB
cnWdpa4t6xS/WZ6oej/oWnlEjs1AoyYviWCkq3xY2BJTXtQ2szvjMYz+Nc75psxHUJf+q54X3NkP
O7TRy1mf3G5I8b4Ul6neQmyQv/WA3X2EiHlY584iWupQA+gbUhm06lURBHknQ2X1+uzZY8bGM/SR
3cVd/xwo7JK8lvAltmYvlhxuGaXy4rOHntnY6hsdGugJ4/G9KN6/7eUD2bzWm+pu/m1Re2kl8P4i
xr8uoJwGKmX1DYf7PG4GGRvwx+syDpqWW4eUot7Fk0W4333dATUT6FIKBAtJGfkMEDHHekhqep9r
hWyl/7KEa4Yu53XA0uNxF20UHlZA3ImsftEXsbVqoe33rSaGDGwPm2EwVuacvJCTmVOHSREP5pZT
l8xYKVxJZ+L2W7dn0XOXo3f9OiAy4awl/5FRflEK5z7pNkidRX4xEuf3PnucHan9K6OWLEnGZV4l
mb6iuk2WYGSFtimgEDgx/bQQWMUiRAsiBAR5EV1NNFdgVmpEjKYfALrqOggm0eyZp08UOotlZsDK
YeGFRrz36Ae6yOU0XJoQ6o35Sqw0B+dWqYkmnRCxKQkIKkZlUBRol5SmzDmpwKXhRvlXjYdE7srH
ceocWIDhgPsv/ddf9q/XvxEY5JbSiOiCGKnoKr8w7DvxHYeuET5W1pbc4cdCJezdRyAZINpftSt4
rb66ncEBW8WS1eL0h8sJcIGx4vItuwp4m2jXg4OfOM8lklePGePY2kZ82SMTUAHr1BGcTtMpYKKn
OWau9Vpyf+y+cjFmHXFsZdgZtpXH97/TzGRiYAMMvTHzOZRqAjP/ZC9kSfxFcGbNqirtH0HDjTEo
moBDjh1d1d+Slau+lZsmmI8DBs2LMTYINEuM/gpK4wyVytS0/zptJi9QOoKT3dlaVRDTX4dl/pOS
YwQbF5JUp9PKuDoIFWxPLsat3Yi/ph1e18KQjBbnsdVITIhNYK4zLLogIvtE2spmQiKtPIK3UCXB
3kLDvup9oyWyuAIrFdfqIL4IiepbBr/IGWE61v3ZiQjdROVeRX6jXK4Vyc7ymOdtdWxi7FjYA7i3
l4bsXo71RQrA2i6Fi9hOrS7l42XY5lZy7FT6XdE2dRm+CMrWaJKrYOKlIpq96kKv+hcQgsKxxrOW
9xyVt/0tUm66HMG4ozz3DtrslUHuEQweCvx65gYwuUMdo6OYbSLReJDTWoqLvL/8I4qAFyFFDUBJ
Qtk4u40FG9YvMRa772RIa19LBB4B0dqGWmQEV2rPNFbJ25Xwg0khW4pF86fHBzUZstcgE1n4uY2E
Oe36sZ2osn1v3lH4B9jwbbGFSotIry8FcreU1IHsoDdqBSgF6lNgHD9240npX5vQo04aJikeVtRW
pmhPsVW7otRBH9GNL2u261D1vzMz6cxtIr0rS6iZVsafE0jG8Q//SSl9i2ydTrfI4Hgbxz4o21ik
vlkGoY7Z7Q8L35JIzSV86wdmD2qDZ9QtnE/5iSfNcdrrvnxDge//R4YoPgCjP84B9lLUWldUpRq+
r42iIWIgeYZXW7goaR1jOZs/k6xAHbXY3AqtCZIyEyEa9IA+4HYntfe2FcvBaxtYKkEwq0qlolpn
TauwItTHNHoYgmXNmWw67HE1Dw/m6/7pvTdprgBzzVrcSYlsq9inFmI5xV9xJ7NR/npS/Y4sf5vJ
CAv9ij6gylYY/nz9WBlDjHa34HS17VZln7777aA9dOZpqV7aHnUL5lujpMloYOqy2cr5qV2LfLTO
I3NV5y7TGeHIbv+PvYsZMPja7ox3y40sI2topE/Vag6+NnqG/AyI6LID/wyBd2W7hJrmSgmf1Qck
3A7svOlPMRvBkYOilWjjKLYT31uILCpbL7nB55MbiOFjgMz9SKx3guzl1r8iGLtobzt/g4agv+QD
kX5t4Ui6XnjWgTgo3vg/oxZ2m9MCxGYhMCtmx2kJhnzQDLF+5XzKMlBORnWVpAlU0cQfOwecW9EX
weg/wm9tXfUwi7iQPM0vcAt8/Pm9wPzL+Q5faGSsW+CTVK9mGkEAd6hT7IFRJPvuW+774/hfOAuz
h0qdRUxaKDL7Q9wT9F9CWsB49NTZVL2f4FuVzIEJX8WVdeSdEl34vAn5pWQ9lZIcrdL/GIimzUHg
stucim1oGAzd3Rli1+gV6X0S5pqwRTFDInLs8xam1V4i5rsPz4waIX8bfxlNbq0A98HEFUt/sPvc
sRDeVnEi4maC2dbSoGeIIqSPFCdFB0b/jrzGVvV8Es6LNirE2IWpOrBNzy5F+7o9so+u0zM0GDdB
H3t1B56Q7+QVQLpL9tytl+qD7cC1rGlGlQeuXcdqOq8qLmvwhfcvQukWBZobj8IjfK5jwm+2oBnQ
O0jmk/RsmjlEpjnXc02C3HUK2I6btc6jiJeNWTPydJ1xPTcL8wbDASEQve42P1zaURwJtAyoQ4i+
UvRnjcKNdiAfx4y4llPnBNQapsyyg+UqvS/tokaihT2JLpjiad8E1E5s6wAd5Ge3+qpv4W/SMO0L
+czVZj5v8adquSSObugoxwG4pod2RXZSSiicbr2pxEfMqpdinLp9aGdzrmD22CSuPvNzEzx89t/M
AnuYuaOxxeN1GPI8SBbtdVoYeiEmew+RVnR11EdcijE/RJTQbvnceAzSXiCME1sfDzMScHnAalYY
6nho45FQ4AkM/sGCVtTtQddAkRyCgda5InM+dD/n11rBYAo2MmpN1irB22rlbj/TDbz71XB/shPr
U27BtHsbOi0qT/W8lfPZDuQ7e7qGTsZx7tb78MZNHWGOKcCKKbar9iVAFOhwXNREIMwJluYLF4cF
p+sDdBpI21hjDITgP83eDWwdpsMWJerLQJ+x9lHyHYDc9F5YWaXAnNGBWU/LvC0Qb5x/sNTglBbv
xrEGONBxtabcVgL1SwA+pqGL5YLG/QTZsH/F1hcmbFAMX/13wYlKjjUpNwP08x6snvkfzaDQpxF0
IxmKxBgx9AQBBcgB6FQPX+IdK04/89voB020B39QEMtiLCrwlq0sojfTiUduEgrbkdLl0lkgRWL2
GsP0WyTCBG5IC1O/hpEKd3SyauTD0HH4hSWb7TGltPouNNOlxHx4LHOYLFpcD/Ly4QheLuMZlt5i
JjjeF/e66x/xMVWgTNzrVlQDEJw6ZuC053f9hWLtUmuf3QhCYcUEM2Qgq2dfg0hySFCF5PLdbodJ
QWAK/vf4CblJ0RP1ho2dty9K1myid0c3h47XkNDCMs0AXGZAaFu8VuP/xEnuI9HMZJ8/LFGksUai
jWNBATa6FJKgJ5ypsKiH9qtjFZJ1F/n+dhjXsUMxhE2mTc52TXuO1x/DK9RAsyfLzUNZmBevHDd/
hV/VvqaRrnJmtxvGifTSJAZPcYwcf/0qYuOAvJPzPqdOiH/rqFpdf+vHiKq6Z8XdeGyYKqS0XHXh
9uDMslpkattV0Z2toN0yc5W4hJmKUO8ofYpmZH1IaAVwYr25l5yA8gNNSvHdv19bp793wUkxCgqA
W2fuW5DYwzHG3idoohik8OdlsyNXLy7ZOGSPj84ySWpyp1ONLrZS5AARNMpp8iukDexXCNUwdVnp
lGhOoI8stpDTBhks0LTaRnG5beUO3eZa1Lx7pwrdBTXU1GRs4FZALaljvTKpBnFw407xfIiGj0lN
5D1LQzAwsUAu6MP0XVa70pEG3FeUbrJO267797HAvyFLTAuY7mPGBcqV6iIAPuLmszTvbcmz4kwG
I09uVDpTeB6OxVEU/+Kr1QTAl7sz0ZD1pmFtZa3eCDJgPMJXA/mTYMrl2ppI5ASOaueV2YLGIZlC
do+/WBxX6JO8Xa3POLgrjX3GI/urBvoPHcehn0MsJlXjIlgO/MaaoTISDwRswIDdpvjxmm08G7T1
Prkty0MzHLWP3RnWikLYHwZ7uy1z71C6+7qe3kqUUDRbutkFZ21RnT6JQcgw84yoFr+NaJDEopvq
o2k9Y4/digbrI/nRZT2molgLVJyDt90+tyHObcj2GiSG0ZnoHeHD2vCRTo83nMHdkkUtcv4fxd0x
IHMeUvVGfg4V+qvcieuRUs50oWIHPkLI/kQsFWai2rR9gw4NumQbCYDRssvv+v51d4zCxn7JirWD
gRYdhRGnHp94C9XCUU/RcgEKnaxp45TeVZdRldnLJTnxUD8snzYsze8tXaAiRIRiYTTz8uFHPLkt
7bUfdPxqNT+e8r5Sxy2Xy570/9GCwxcHkM0s66akIULI6GtqZS8k13TJKLNAyQmoivdLc2wgiIKV
o/AaGaxpaKH7IVJQOIo9XWFslyM4cPEcF5Z2SkKAGuTJHIT9/LqyAu0bFiy9BiUYU1JPoH2d1pp/
fwebAUYa6VowA6o9iOSeo8Ov09cWeO5/2rstGLuVk7XAnL2HZPm9sRmfK6HWFfVT0vaqtCFG+Ho/
LoK5k7AiqqHQqKUie9mGFzIZEl9rZQORaSjrYS2lRa/BqeeIdjBwmQhW4DiAVbuNG1Q8zQqPsBQy
puRE9/binldBA3MlweMoq54aUivIWdfvuPDiKrg/GrvSWnfBKPiIvPJtQHdgKw1yVltwreBCPc2q
s+1M9Yu5nVn8yMUjOi18JlmWPwMVeaQv5s88lqCDNN5G2rsWMqKf6hUiu95M2kleTRfvkg7NdDW+
l01FK+4vbQRtcHV93oHNfIGZrAiTo6z/5JTkaldyuhLdIrZI1Qm3WLLr2djXQwaT50w6i9QRv2QG
IWgrAw8Pgnnso4TYOa99t45Z8me5he+f/CycRiLAdBC++7ewofAqkbCYFfOK3HVukcuDXCGv3uK2
T/BxyaYTevpWXyLguhQeHkCa3rIhwCq+8ZFXFdnpyA/AXV7owYiD6JIjpC0GjXhCyzbZbQ1kTTFT
lGMI7QucuWAiFCWCjQRmialDTYfgsXX6jvf30xwnkRCuYCL8jldKyUeCNDPKriRoez97m4GvUrx5
rFdtLzqb66snXEhEFWR4eNC3nkm62J/4roeCdFDAB+0Domu9S9RuyNNvRHm3K7kG6gwPgBzvamUv
sEjMSmvukAfwCUt5diiRzIODukYBRTOo+0e1UuaLAXnlac2SVwMVrnqsVS8LXq8Kty3hSg0VoGqf
Bh75q/NaTxWl6ZrcDjxwwJ2PiBLgZVoKI+oAhBDG26W5rop9+rC3Tu52FP3d2YjF9T4/YlfDopiZ
/E95Mnf4goh7+ZJyvEfkxZPzUl+RimZGLrv4hkUr6Cxz52TZULLp+nZuSGh/hC5OszafgBewfI9D
bSaVAO34exAE/QDBHO9nyc0o4JEG4ThNhf3mm8Tr3AhMgSurDnuu7axhMkF34N0FdDZ/He8Qrwkf
4g0m22PJRDQqqdRA8g9flikhd8Ll3JVPL1Ri4A4TI26zKyTYixwA202iTs7ll2Pcx3b/M2wrDqCA
zFC+sa9ufgm43pdLYHNwkT6XqA6EJNlo71s1FrQsk8hyf/z2gzbfOJz1Pnv7OPo0Nhz0uuqRbNq3
RVOcK+vsCAHwnmUD7ZSifgJ9hHv8e3gqZ+pVZuN6iaLc+0++Kr8Ho2bM5KADgCC1kBcLb40UCoXQ
OqCPl4bGsLt8aYT5rd8PkELRUzIrMw7akiE5semVA0LIBZe+nojaMP7H2JXsOx80APouQ4EwiTv8
ZFNmo6zv49VPe52GMKZ9RStzlAyKZOivSck7F3FavfQDLQSel1vxAIy6osZTPAZiga4OAKhREXwK
4o58Y5Y4uepmaYRsHkMx1iSm4swTvYG8TGu9hcOszRR/sJRA7W5vAh4tAu4L4vtNtoIDxWVeew9R
ycqzqcczF2vxjON+sOkaqZHX97a3QKBAutDRGpyy21TtwHQIOi2IJF3gAziAGFZLk7iga3aXxrOW
lI/tsfoY+yh9vxWmOFCuOj4jxJi2cfx2iP6V8G6WDqQtQgygoZTRHTGMkGNFZaRxxQ/2DZiz59S8
0i+EdWVh/QAjeyuJu9/qpnEa+/kd8jdJ/br6gZYXwzsiF9WFuesxFOP5lfPNBuZcarrvOnHFXI84
6eyRS3PlJ4+x4M9zq6zcswMp2TBKuhUcKbmsZmH9J6IdecVANsUBgBwGg3lJYBYvCLFryfvQby4J
hXjC3aO05Q/SZfuwi4gvqi26N/Av3lqS1r2fqJsZ5xLbvAPUNA4LC47BI1Cs4Z7YU9V+IDGzmgpG
qNRxxZLaHbdRUpwjc3ACTUvwQGTBUu0A6LRj/CB1KrPcb7qgef3jTgTQ6PS9BYsX1zL1lLdQ4dtj
M2wgs4VYyoxfn1C/t2zBv9xKKSc5zD/o9lXQHywm+F+ZkFYLj7WEBlEMFskLz1J6+bg0BOAdF62i
+yNvMaOrJjrYXcpYd/bmFBSHIIeBkrv6Ba5g4443Qmq5qQ1FANGx1F6QB+PTauXlT+JfJiFGOB8q
6YE5Nr3WSzJQ6JkzR7FITG3vo3dn0oCJDNXP35fXkySddfAgydlJ7+DWPO3vDeVce5boO49dHFcg
Pb0LWuoI/ZEbM2r5alpJgq7ar9If7dcAEUKrMFNDL6ujZMnhOwV2Sg6pE1XMl+PWUacKhAjrE/JM
v6JBCX7j9IPQALO5hEImwr8KNY0dNUzmCOD5AgaLPgnyFRF4oiE47Vvlk4Icwp4Bzr9eBr+J2VIp
/x/pp/5esT33vjsdfDupZ5AuxuJa3xMgP/4Ax5bcB4pnyPd7ux2+3YMUD9gPPJC88OYo07VtLdF9
6amZZg2SiKXAtkQ+Y2s6SdhiSaTCqP8XjW3TlXEcfkeI5hTyYuZM8k03dAmWj1WI3qcbnccnosCl
oY3WTr5wQ8aXbq1Eb2Jbj4vyqtQyg46dolqNYi5qcwapC0T2nRDZPAQ0YHMQLhPdUc+qamXA8U63
z56dfrhXOxm2aftLmxBTvqep4O9Ft8Xol+4NXpraZl8RmUF2Fr12/kz8uTa9b1VpSL3HUmHvJffv
I56z0+VM+HcBHvY1e+8XPHNOu/h5w7mYKS0+5O+L0WY49a5Gy2lcD48DM+/bpu3KFQ5NJpOc0Kp9
F8P/0IkFs9P8YwuWnChePWcL22cvNmwddUn3rr4QDJ830ITID3aVDPfZrfNAC72xyLRrg2SEdv9D
8R81CAK7xiM/Y0qhQWEWybkpk4MxmlAOl2h+HM97bZcP0UVzsQUjAE6hFKxGissnGXJKKm4wGdBl
gEmCfA+3EAc8uc9TOIqUTifnMtk7zgpoTNKoIFe2hh4XNpVTa3XVCzhgLEaEdwYRT6qBDdxGJ6V/
YD5DlWfGDwjbAruF2evcJEn28+0SQwhUFRCdZpI/x88eNgC+sMDGj35ugrubf1LeLAPImQRRcjb8
FAQSt5onPfI0v+VNuF3i+bkIECzGcP/NBaOQ9NAkoV7G3Q3rS4SxwFghtGScn86rmnZAvq6T+SOi
f9FEL8ydeTCrT4EvsOcILiWr5ovEIVNpO1ZZVY7kIhHYVI8bc8p8opbGoPj7ay8zeRms+/izlJxA
5+isvwQPyCDtf/3SFBZpoEew2J46qx27qc0k0nIaacnN+9PZ/AQ05YYlkKbvz6ruRi6QRsWEa4Zr
qrOBHekvlcKj5icJ3VPfgwTbx1flEnkU7EHERnXwh7ICPZmHhjgzcIRB6shBVFudDLxkO/xVR0l1
GkBTy6SZM2BhQSB0zv+4mTXJGTAwvREiilYnj9hFJLzDnKGQfg8bQUAYit8O6QIJrgQSpIhftXAj
PgLM769gEHpFb35TWEkRgV2IZuG9tLVM10nTO2PeVZlHJkg+Ic0MOjBEhuf1/Rdv1skWMp7AWCYA
SnEeGgYbYQl0B8dQ1yD1MoeSg67egbu0TV1+HpfIuJ3L2qzptQ4GqJPqhqu6YlXyafqa3xCXxTl9
COQMU3VxX63uJtmX82ywRM+6HZVq3VG9LF5oLJeVFaY5WkXPvUvcGQ6LClCAN2A1G6DEguwok3uk
S6WE/KByrAFF/TviBEmYW0BCOd5ZqyOTK0DAkKtCkDnq3rGRPlWeQhHIzd0AetsRl7xKeJZaU3aC
i2saitANhgp9vtHMi8Yhn+hd1STZyw0IZxmHdcIJg9w+KX7E+7mZQkZFE8awQ4dPrHmpdMd0yw1i
bj+bIQpbvhpJIDlGsi02bTwoyd3UB+gxLSeap3tc/m5/PGXlrgUVVgj6oK9B1whXT1uzdrJI90x1
2HPAHo2z5AoYDNp4eMWELEe1RitNXZ0SsLbYJWtG6na9aEKJSPBcBTtz7jBVi+Tofu8yJR+D2C4d
BawXH5VAEJyx4zPt9x4DH0DAKHQHOEcXv/UYBFcb9mk+VXepO8SZHZ7/IHa+he0lDa+3BcHbkdmh
6UqnHHH0qGrZlak+kQH+9Hkl5xbrXp4S0yK6q4aagl7eiThTdjV62ClL20pGbXoh771641MAwd8q
nin7w5lPVZW9gLkkLf2e+lvb+u+JkgA6d6yWxjEUsVxE+MtqUYl1ZWftIra0Qel1P8MmuUvXpubX
kn0w9+BGmnU1usgaa/jNf6PWcINK8LDiMYZaooqHxKxFwtw8pJcPz1RV+eYDFc237adA8c2yGnEJ
+W61IFoaL6oLCPsEWb2tCNo6mm/EQBHhFL0uF2fkUSIZdjEB38RI/TAuzOjpn0MSJuD7c2lAdU7y
w3MgPZcy8AGA2APIvKHR2GZo1bq+I9TpyATdWMv9Q4ldHI0CEJ9Snq83O1EwJOb0i6ab8wtAIRLS
Cg2dKYcHNEJ3zQy+Ek0p7tmUKvVLhR8PPx0MRiwPpX5Yw2OLIecyWnS3HpXmDUkPlh0XNgepKNAt
vKl99NYcjWpmTB5Xs2qDxJ2qOga+S7Tlw9Zm4Eao0lcdAcIoGVsj7FpDj8b3pBNI3bzc/1rGo8vz
P/5YSZ6enzQh4jIXKHwu1bRdJ+G8VSza9AnYg+B8wc3WHue/t45uuqx8kkOrdazI8l0wmefAFEjC
dT1wxsr2y9ZqXi1jOwb6evNi6MChp4TWr3UYIDqMFAR0NGGEEj9T4SHqtaSTfbQ4lvqqM8V9e4UO
HHzV1cK8F1jRLz31BxLHi1jyGP8BiMMStp1atTK/FkSs5DYwoJGxaTaL2oxN4BvT5yO8WrElpkRy
THJwFwtuav5zkr30bZR7a5RI5UpteufEsCwwJbPXG7nNznuMnT1FalU8BI6+ChbeOmFjY+11CZ3A
W/gakwz/pOBrsm7G7BruJg+4y6wEYl5B5qs5K/BZsmcLPfaOKSm4C3KVNAf251WFt/2HzqGwFZSh
nWXsXtjXkkpdIV4bg0n1fj07xpzBSnYngiJOZBfNtA683Aba1mIJ3YLUO5EJ6NvQqpaAnOf3NFXU
fjkN/15SXsP3b41/s3EbY6x8F/afokrF1xlsaOtRrAcKTFw0D+cjhTJ9PUHRcoFRSCnlSu85zMLT
0WLEfdTGKuqKTgj4RZ6Byj5C81d5bNvTC9CiZwUQ4i6bH+EU/PTUbtkv+mw2j7ZDrch9HoIsHoI1
39pC+UOYft2YDEGnDEn5rSEtiv2oj92TzUxRqCdHHF+zCcdxo/cVrtrka7fTG09hYM6EOEebwb5s
Qog8Gd4BKY8QLZnuzSJMONvv/vDAzcTmG6AGk8mmuqF1CPJeNRDdNrS0E2/6FPH16EsjYRK1+Viw
2cRSVSEXVUS3NtEjMALBhXWUpHUbhs26zeK8qaaMrJiYlIadl0dz2IqfgLzaRQekp8rk4Fadcu6Z
f1OPWtxpKcqJGJ0vujpAuujBHCvr5J7mNYp5+kyvKJsraDavQ6U/zhPBymuycTpOufbKy4wgdVMF
jvf8THBHp3+zKjIkRxUx2sMrOFgi8LJznwA0pdGCjNwf8VtimQfxkTUN3czZsGvuZnScxdWyfeTU
INgYXuL61403UJzx2858Z16Z2FuY/85/poRf573CAlyHKleRHTSKJAAlymnWHgrrAuGryojfYB0m
QIRdAsNhTxSbRiTvDg4EXp6899XPhk65MmoLFIcfLNrs9vrE49lYcxJ3Noeh3kwHIwVisWVxrw+K
Jv/HbkTHTwf0bxMCZT5p7vNP2qFmFsrqIjSXqeFc7ChJ+9KAaqM/gjPyu63wzSB6Gkfq7/cY+x5d
m0VesZBXQn+srY09A7CEug4WGX+S0n8c3/OTDjtvFYLjhU2mQWvS2UqgMKM5dD1nncrGq0ogbSx1
TKUiSqYdwYCu6XAXUhMm5CecqDHBtDllL5Pt+QSdUmcEYGBVytK14koce+Q9bh4O52nnDpGD3l8a
Mn/9x+KqPHv2XpGztXp8HBhF4HlqmeRizo8K8a0Wv6BZyqtgRVEW6ncJllskYiq+otYt3vWnco96
pq7j2kR0YokLNkAYfFaFEuRlvwcPTpoHZfi6in/salVWdBWMxmWuQ8kpI9R4P6bwZ9DcHZYp0bPF
JnRUVod5yh5lPryq0wP7GirtdqcO1wRGM71x7pBxKeCJ7QfETnKjuZ9sjsLnIwINwflNdZMpElP9
etuLsdafwWhT6kmYi9dhhv1UlG0B4Y/GOGfSXwb8CogUxQ6XOCHvGhNJRFZgtAkhUEe2IgbF5NqP
y09+AuWUmsX5VUTX+wWJ3CJTXZILgzhqCyCYindiJFjY/1L/LV+igLE9cbgzyhc7j8w+cMHyrCDv
YpBSGabxXHhq7KD2F4zrCC9VTyrYuy1b4bB/NbHAz9CY3ak4yCdF+gIGbVItkv9VRGHHW0ysqDKM
C9x0jX5YyX06h7jQBcwMd4ik1InaYKGeWVTgjfcG7gtjdmqhdnYehv9MhyavYjD89J3x41PWtmOU
QN8NTqUBTRA9iYGcKHf4pfNxyQYCuHXvf7JMcuc3HwTlXSprmTMMvC0+J/q9Af5jiJzUyZlJzv0t
4KYS8c9e8dqOuZK+Bw2+auXakzJpI5ujdl9UodO5j+6BABWDSph9PL90KlMc+Wwcteh8C/CVCrYO
NSAiOq2JZAsIAXKFyZBCTZ9JoLGQVFwOeDzbhqAGw40bOzyck1S4PPRwaWaFYiB2gTnzlXttW/gW
KveKadwFPjRNFa603CCFq6cNQ20ppwW7LrAsqjGUZRN6xZjO/dEHd7H0kZEQvdl5WnmbdeRleOXg
Kg2HgNRhJK7BHg+aZbFJdwNL4oXu1iUvvk1G0Bvwlrbn+KlRNGA66RfF6e70oQ41XO4MhNgYu4Si
DbAxlKHa3Pc43PubA10tJJ6ItQRrqaH0rQa1+euMo8YnPn+0Yo/L39e3fIhGFCSoyUQgLiXn3ApB
cE27wEhrJoh6AgyaZlWve+ViWDMvBfHch9WQy89Xxy0nMwOWbmkBLGFuOPhep0ghvvftn6hzVC4p
mU8HuN8awoZo5bce05a4KUoPuXxP7KtKyN1RGcQzestI8Fq/TBc7PEPyKx0b3bjBp8x+cBTLTvQM
87f1b++Pkkf/r587QsVbD6BhVrn08J8QLNxBK8GDKi2nebZ3ywfdk9gZWaXksJYGzKm+fZ0ARF5m
QPI7w0VoFffuYeUv76mQzvpR/tcEoJYTFXx86p6zNbD3c1E3A5doAwgWDc+liIEBPdjtpuQte8En
UeDTf6QPDrsX/pfZRGAGucvc6eioHkMvLxW7liEOag4ppU1GSR6dQ1CD4Gsw3faeIZfAgdwjr3qB
ok8dI4dBW8IJZQBuOXi+26x8ouizdetA3p8FdR3FlXcWXKqg0EmsKi8AARw9nO0NDMvXZ0jW1QUy
Gc0q/zwV2q7qDqSDqUaftV6dHfXncEaDGt+oUU0VuIWtINdL+PcfLAvnbIxg14x1jRu2I0uG/5Wa
SEvzdEYqvlwm4AfRo6YOXMdvx+SjMPc5XZ6qHDr5cLsOSFFRp2AV9EKhB+ZAExp9Zo8A1HCXuPT9
x4pZytcV8siczLXFdjwFiXPJyS7gat62v3XRNratCSHBhVE1mdcB5N1aSzf5GWMpVym1nUHyB8c4
O1ovSiLzFqXdLFyna+/fxQ02xwBMADJW4LGfVG1X8q0YclSquzDkaFnQPWWP/kgHfg9n2dSJO7Lk
gkHTn2NWPcrnUBNqm3QbtMaosZadgNHf0yUPasqxBQXvUdsyBJj+przv25IrsOE8aCWfEvPjq64I
pBk4gmC5rMNdpTrmI8hMqpbeMUdDxRLyoooafS5S2IRZ/KZ3u4rwz5nDQtEtRsZ6tWrgjh9hd3zG
l9xg2aa07XbNw3N+DWy1+KHY8NmNQJlYbJFlyBGEWht7I+Bf91z0JhZWjxS81QXWR6kiabI6CAYU
sqJ54IVtQoTJWQerfFlBQq0wGx8ez30C0LEtfnrpBPRLFySk0y8V21JYJLdMFFv9vROgJE40263J
q9IEY3rVWazpotG3CTAE4wfXU88VE5UnLS4kiutDwfp6UUZLfUZQaOiRS8bJLFcVYSws26puJJoc
iG4Zor86BW64lLaLIiX9z34Xbw2/E7+wc5sNcPiUwTsK0InjZ6DkEBJYJKP1hMYq+vsUashaRkYf
WEfHYGTzSiibG6/v9Co/woMmxNc7jhvHr11gIHXVnmpFKi4B7nBiwfgHTmVCADs7QCT/CzUPVKsq
bT/ZEKcIOz8ALObBiJdL9Wo3nhEiNDFAskz/nQRk4M6kCNj+EQqNQL/5fsp2rQWq0fwElmQi8hi8
FeLEkw35X+XxbGMk2//qXvurowPJ6/P5BzRTEITzpLp4hfzxHsHqh9Ko6mrvlS2dKODZQx1OgQ7o
so3oXcvGDB/aW2jdG43TNX+2SQDr2QTfbEaxVYDLYRC5IjximiA+Y3MENjHnxMuf8ehCiPcxYKI2
UYuUcRi2NsD2FC5c5S3NCiZQOkSSCvbYUmPY6jjMzLX8yY/mKVHnh1+e/w6RyUKROoqUuHu2RYQK
iddwe/2SoCQ0kZqiaCCrH4z2rqiIz3lWkEbPCyDASggyKzpfQyvmhCTqtKRid42QNxKvcGxR6vem
+fzLXHzi+vzljSc5pYFbaa3PtGBpSbaGzp72H1OK/UUbKUtkjAk8NtnNbiep5lVlNz6Y6ykfpV8x
NAWqinpEh02geqxoyanNW6aPBhN+IsddpmMzrvUokeWOAFD+b0iBIyLGhlvwpZc+4NnhmWvi6/Hc
R4aVw2fJ/ETuMVRE7TcWoYq2s9dVoC4AyZs70MT285SUvBNWS1NosS2VazEPw5C4oJpnnB90TkUe
yYBfksY4L0h2SEz2Gm9QOF1vzMVB1xwJKAUz7vVeGOp3r8wl0BYNu9ag/Yi3YJiISuTN1XYzocYz
F28+Ygfe8EP6taWcxpUFqeNi/26c8HtOYIrGaPOJRWi1xxSXWzwMPThLxKjr9ogo5/xPk8PNhRal
TIEVmYS5oD5BD1OteJy46URWD4YdpZeNepnRNfZsyO/pTuO9+eWNj2WzQ/X+vtx/a+8zjQvX2ss3
t//EmrpSE51gPwosD7BEXA/WZh5JqKt4Gt1KD7fLg7CNbpN0YxWY3cn3qUM2nQUt3UQwCTi2KT88
NF9P8IvtfhUssFc8X0OuLELVW+1G3FTR3nwlR1ODuWakuryZ1HFeljbd6XDpqp5udqHN/mPa1o2L
TXOYKuWpFMqSSwKY/N/hlALFZKyXkxTXT1LUcrBUFS/Xm5mhpPt95R7L0oPQldGHoECA2pUR6Gt5
D7v/cgr1EYhCfha3zjRpLVKwtWVr5cHPdsjN/YNo9Lfz6e1RpqSixMcfhMMivHNfkv/LALCPKVdp
y/B65+0dZMQYCIsHn1AXLxwAKFHsowLDilRF8BKdwph78l8SPiIqmvaItbQjjfQOEBOqSzJHMuQ7
XsHgxdTZfzon5X4HJP20tJnMyY7vt6rC33QL4I2nZyDg8wGd3xcP8IE2BANtmflvW5q3q7XsrkUi
Hpqx1wTZWIv61uFSGhBOq2PI0qXw5WmPbUP7ftBzfymqWt/ao508v3BJpLI1Xw0d+qKX1RR7nu4H
oHobcv6/benlXt9AW6Qsjbd0G7nKesyUH0lvQ+rOKFNbVdIc7KJ5N5U6E1mHoOjwKiXujO93VmDg
aIW/bLo79Eo7wvimGK241zj3R0UGFUYz7vJeNq+W38/B6dQ/SqWCSVTeyLfQlOHTVhfida8KnlxB
kLdCoRSh6NY20NvztAR4ozajheYMSAZBU4tkW+r86al4hS9ClGn24JcvN+RBF6GTd3Prc1N0f/SD
dY9cObujb1SVt4cb2D+2zx54GoG8GwJtybPwNhvGx+iXuRdNzttgrF3ctb0G3PHDuTDaKGX00qw2
Z02iuYzbuoNIrTkQJJmgezABvksDCSvow2rUKAVpwCGxFIgoKIzezsX2MxufyGrMpz+BPIRzH6G9
O54TuUmjUs78RgqC8dhFlZch/swCa3A8JEmu8xSPmwntXI8OIepJ96Xm/3l/G94KLlxhTl12Q0Jc
0NZNlppQAQD8xPfDsLcCAkR8VqyAvJwqHFfJGbVrtI5IIwe6m59VIsrw5BAles2Q9FZOy4i8BOz3
42PuydJgjbYJcXpMOZlSW569p3dfRNXdnEYVaah2M3AdlayGFWdw19oJUactu/ZTQ7H8ZsS1hEZ+
FR9XM/rZQ4Yq/NC/i9VrLSlvy4OCHD2jL7LjGyMHcPTs9cJEXJYedWURitdmbDEAJmoX9Tb6xUZ3
+ZgYSlMBiFFSBJoVGLWqWpH9fFoyDUG21uPquDrug5cgsHI6lYvpRtav5Xoi2ultqEF1D7qJyFks
EoDF7poW8NRtU4Lxhh6g7VoLZw91Wm6Qmw/ykBXzQsyKJL3wqmwREP7CXAzHXF5SvUlRc66j+VZ2
ISPyj5prSF0s/yFSkMBCLnoLSlqf4KZM0vchItbNlXOHvzr3RwAEh/0huypaqm2ssLDSsl7T/N69
rohVyFmoNt5M86n+2eNfg0jsjpvVgr+7ZGkmfrSC1SNrei3YyPCbOlcvJfqQM+lFH2kiP9Gj0T9+
UY32GhdN1yeju3IFBAhK1ox5cIuoOeyBtVHKbOIFgcPZMjYPqu5wyRQmKpsocxYSS+IfQiHN/Ue1
hCW0BmH9Z4WCnyMjr5JS4s9bJVQVINSTu6EOFS6Pkd2up2Dvgwez4o0dQqd8JXZ0wvgXDcVzLH9u
h2d3ayRGxDICuvIsF5MhKGSdMDnK5LEF317MuUL0CYBow8G1w8B56aRlZvey14SC+YZ84avxRqgl
h9CgJBX/TnFV1Z2YPLM60x+4Gu+PdoWH6wopfo1DhfMlrmxIK6wx4WOlUymANAJK6jGGV2CC1/CX
jdmmhjFVoMgvbGBAF4VFu6NA12ZaAMtbnEJ4qcZGOOvqJMKq/yEn9ZB8zUBdV/U9+nITwfK+cdeK
z78MQiXD67rQjwRm/bI3th6Q5T3XdDoPdvajZcr1nL1P7aXebHmZtBiIy7AJP9wKuqoi2D3hDDrL
KcQG/UsNvg6oUY1cXpd/giYCo8LfpoBWA7U70lMgLk3B4SB2FDJAb56eZYq0FpqQ8cy8hMsMSSoP
dFbL49ooeGvuwRvcY9stk/F7FqIL+0+pH7u84AvERZGSfRcl93s+616F17ieBHpOfHYl0IljglQ0
IOzHAo5Ub4fgjaV1lMN++kBFvaf8Adl8w8lyDA3eKGoFirEEYHrG5HJAv4TBTGCGvINOLlb2OHsH
HGNHMmNkfRKvwvZpHJ4OVfCC6fne7S/Ee8VtKt4pNm1H4p6VSkKmfp4tMwee1YVucAzDNsjXCO5q
9P8mWgcj8E3z98sP+ECmsCPySV0r1OiqJPxTrmQoBTRCRRsgErtdKyof7NKtzIbJndOuqzEzRJoK
2SjUBGrUZqweq0A/FEtGhpaNvk4NsRi+/DNyHMX/8+SoA0sJj0ZntoONQhcoAAaIzwP3sYEuIoxf
HOUR0PeJCGKPObihbwhCUOQPHxb4HBtN/vSyn8HNcxNVEIz7z3meM0L7mN72DaHCTJmbqRBWZkes
UIgQXkAeq2LU9+FgsRdY77xhd76Q+WoVa9ExHlyOXxa3+MrmSAK6shZlQ0gmqFeHJiytJhNqxWY/
2UvcXF9XDz4pJaKoG4gc4Uapn1mVVfawM9qTiyARdBjkAcX14BD7MNsZ1iJyfyy+tYYWE10UrAlf
7XcL9vcB3R5NKGtQZCIDNa1s2SClER2mvqGDx9ID9l5ZqL1zozDCaBfUXIUg8V4RbOs47mLA7Thc
5cyNd2aF8ZG2lfawhaCEHsIU372pHAPcOM2brVdLqYY/xwnGHOp5GBk71yRnaVW/Z68l6qh4XVJL
jmnwWzoBgemZ7QJIWiam+KFzVE51hNvN/hhUcc1vf2XcKcqHYM/1/C69Rhiw9KFB29nUnf+e5hg5
iPxhS9F+7nz9Zc218ZQx4p27TPmeBVq8TwwPpBoHUXZJW3xRVqtWiBJV+bGBB01BLY8j1jxlThyo
bl0GeWQBsXjq3dPYKMJhmC/ziBNW9nUSlvxkYANifVPYwJ74T9BzsrlsuRxiU85UhXqP2yEVmzp5
2P22IHb9THbxUW0KQfsg2cWa7hBewOnAuhti3jT+rOvHKgDhsGiKmbBLCia3/UrH0b57CcQdzaxP
EUoRBUSsuvIHk6KkKMngBelmcWDE54csQirXzSCT6cwCxJ33EZJquQa5PM/tcFb2evdOWKALz6+U
fHhlBUhi2uTmCUOH2aUOi95J6Tv3QofVfNoAH/5pypTaynlfZ0Ydk4yygrEbwIlCoLJWBTHGkMlp
qg0Rv3FvzC3Z9I6knLEbFBgGO4A2/SAy80zdVDgHap5K1pCgp8p9attZ4GjSidTWAhoTxqSbD4qf
dSNQkCiP0tve+1XEtMAHftwq9AcCowKeoMUPTyyTYW9VRvulp+RCWU/DYVvfG1MDdvQR7a6j5XO7
iMRHejnOcRcHKitsGvvMsQ8L9fNKyLDGKhN7ThBU6HUr//ajninv0z5JgaMqcnIJ5QZ+vw00HnF1
N7D6F0ZlNkVe8x2Fc86zCYwDmSzx3VBJ1pyNMMD3hjFXyN/XpMHxxjvtycq9//xaWNUeVtCnWjCm
BYANjWxQXI4u+l2b1iaS4Mzs5CPVR3Hm+IZ91OSHDTSLpQp5qg/LA6yLw5RYwfj/u1VBS6TOz/km
pyHXYs4IpPnaT8zssPH3n/vTQBSCp/3LY050M67xuHluRDtyqapwAjJrhgbl6iMuqj2Qi8wIG/3k
ySyjjMvRrhflmqQ1jgbwgnQzFMSnjxlyYZCCUY2yRFi369MiVzkWTqFAtN7XolRHJqibkwD2wPoZ
BhwWqYoPVgUyF6wGpfLWB4qRGjKrKaFpd7fuL33kHB8RA4l8chA+9TPdnR3IzwT93KhHBjxtursH
iIJV9wlMggZjgBjrzOiMVw+7ljAoJcwaEkLbHORnm04hmdHyksXnDS/luBGpAa1ft6doCg5yWUC2
WhjaAXvEQPeV+HYb2NR07wf5CftN6/wym20s3vOsupYW8mrr0Yyn6jK1wnHCMHGRt1+DHNFyoWi0
WTbzpJGv+V+GjeEchjrRZLZ8skSBpD2lzoEk6V+JlgucBDLu9CwzClojmcos1l6NfbmtRy5taYwl
zw//mwfrnTKXoKKR6H6FuZXH9HfwUnZQHVelvoLSO7d0Zpqha73B5wkjSH0URmPaNqaQ+0ZXD5uk
R1Z5Zwjdn8R5zh0IpAIMnU188wKnHmeTjz5SJd65xcrB4QCzNn3Zl4YCOODl85QjowYWp8qE6ih0
4SYEWL0VYOwlPjzQF6FhOzN4e4Dv4iOVDL1aqsDJzM0TcruWKbIDGtXgn7B2h4GkuGjQxxPFCDPL
A4CT09bHf21u5WaNSvNTF4wEzhNUXK2CtDMF+Li20oYEr24LpyNOMHJt6s5U/C46nVFDBXyK6Nk+
wkv1LQ9vt7hpNSnr7xwO1FoUqb0cYLk0Ujt+YYi/gJvGXwNiy0ZucGrDeZBlS5ZIa4noiD6ylRxC
yjjLALn4R59dQJFBs6KWY18o+8ukWTvpJztUxpt2xtf4bWvVdQ2wjYwp64PrvClOzGohswM34J/i
nOADIQescrSM8yZk4CFbEWZqxzigLTNTGeIQP2DLikrTECRcKaKVrFe2A5NfnUmAJOHosbZtoYrL
jtdNj36E5Qz+tKkhlLf1709bio7R8fLndw9VcQiE4PEnuUFWBpj4PdxvY+HonGnb0qHmMzbAwIYc
UZR+8v3SGFN6Kr3ucIR5diXf5B8h14sw4A2f/Mfk/E0iLfCk0l8jpTXg+6U3uYP280gyTxZMdkkS
5YQZep7VeTyYsPah21/0d2hCFirXDQ76M5JB8wmZVPhiTsJkeb76Vpnbbf106n/3remK+4E7NZaJ
lfMaQ4QeqiXl7oLEIHrU68QlmLnM3XSzOs4Y6uTJnV2dVpwh92PRlXBdAT5pVGFyRqV+t2uzdYB+
XkOd+iSr59qCGZuenqY3Y0Ny4ppZVzH3P+ITrLsZ+FYYCm6ZLlUy8zQUMcPL+pDL/oEqBD3Fo11P
apKM3DDClJ+SZpAw4sm0bP5z3ONhwl6YoN00M315boaVPK/mWV6EiD8ggqw3/VLNxJwWu2SM2qqZ
2S+hPPAAkXjZQ7cGcg8oL2agSZJr1ALVWWog21BMgC/CF9axG0Qo1/ihhX61BpTqwxRCMe8KeiCp
V3s2ITXzAOw+E/7Ur5hVIl/tSCC5bl7L9HZj1W2lHXXaicxnIF5xTp9b0CVHxfJ7V+3eSTRNLw/e
BPGxZ2HKo7a7wVIcKTd8GnkcWB8aTVMrqLt35QlsehHdW71/YGB4KqwbBxODVhftjVv+Uco7+8Oq
/yIx/Zq3nykeQylo4WFikCxPnAgmVbyH0HzSJVgY8m5QKLLmnCgmjFehE5HI6Y2KUiv/xJeaAgpA
IFEZWqLFDYlwRiRbfXlSwljFFY2jYU1bwXl8MHUY55SPSveySCBr+NknKKGEXcLYP3lpxsCjnSca
XoLZWCOgtPUhPDbq4WyEWUm2DKXbZN/KUEwhTJOlHeRqdV6L1pSAWrtcTOeNVIrC7cZSqla0CxDl
+HQ/RpHmQ0AdTnv8kMvhkG2dYlXo4wBwTJMcgrvCpJcRioXuwhMFK+DqhemvIs8IW4NZqfn1YFuC
iRVWxoIot9yOvO8h10z6nRL8N+O25WDbolyXRDhfNRzeJ8yHBwVgQo03yeEtGE0xsKfymUekzFRr
5049iCwsyuX0KVm0YQk5i6QzKF0JnxNL07e9pAvXe4SoELjgWFs4SmVlyOdZFmQIihphAh4oobUv
hxNibZJmLKm0JFCXyAwGLk2QMDBE8lumQNUHL7Z/mW3CdbgKoIshgKc6TKwzZ4+O/lXrL32yGV2c
P4mLS/SOvROzEAccpePNUT4NC6rNPj731rEbN/FaItEVk3azCqFkt9gnUjILbenoerslsOS8Zmhc
WeQi66beK1NqbIw7N18fYvvJUz5GYtS8jFnrFuISQVpzMe3dBsgzInv6Nm2otx2mX6xxRE+RohxY
W/2tlVHY+1aC1X00T3YJI5lUPLuWn5EDg/O5BbTDXFo3SksjIpTmoq2zi7uYv/NmgYIF6/QIJO+6
KpQ/M87diMfOZ6EF3SHQY5RVys8snUfDwicVBGBtrlCzmp/NaE2PDlg3YgNURNcv4IOkSvh2xgZC
aBawXkfBbZBV9xjPVSQVqtyhM8MedqZIQ2iTf39N2CsQ7dOwBRShwc2TOCcZ63ZXIQyJlIkmbOqE
Tgv5hjZmd9GyrgoZCYDkSIdSTTTT7MM7XhfcaZGNSpmXGITGmZKQDxaDMtuqcGc7V1LF3cD2L8DF
WIsNfGX/TVbo+to7l9ZkVj6agV7B0rM72QhuxZPHMm1tnUUKiG4H81qmWLB/gweWkC8S+3qrjdrD
pE22GGPLYPLO8N89O61cijsrQACfXIUvgap32Gk52ds7IiJ0BrpbOaEZ5OqIdlfIBdE1Z7VeuiIX
wcdMO0LHbDhHY+Za4EpBgQMbsDZLu/UO+Cvk0SJdtriY3KW0nTuPT220adn1WZQ+cGQVQwdAfuOT
DwRKuNCwjwJILvUyNDpO1FoXnLPTGAGDDzIcYodP10WyJ1IEcI1cX4Q12NfSUTsv9Ild3Q+fsS68
IkBr5pDTBfNThM2TP9Av8at7dWPvlx50h9E+cNLhWHH5/mXxnWP2dSVoZd6Pj91RM5UcLRCw6p2X
DN7QfpXfach3Lm7FApF1xXdTDgG4QjiFzyhNIyF+Mg5gMV3tmKP3KQR5lAvYMDVu1ucmxyimBZQl
2djFgq/zOcQtxAp9WhFxUB9amtaJ2KRfV+wng4+h+SKocP00idGEhsj4RXwol+kRHEtLCN6nsxEL
T4lfaa7JsYJ9M+aoL+ymjcSfcITI+7RJSuFFW6Um9JGLhcK5omHQqeVib/kP+QyYSlnxgcI5A21x
rqs9Qcavgm6JJfxdJyxoDXQhhKxojgy2KAaWj7qhH+lVmQCGb3+hDwla6pL0CYaUhQRvqXWUiUDx
iLph5oBLEBUhlMSWt1FpC+EDHGAQbAWtp9Lxndwn7mvS1b+c0Y8ltF5H3dv9u5Yb86cOBvKnmr4u
UhNKemcXmEQvy62V89V/UlzmxePw85h+4dgN4JI/j285gQIHWa92BDxYZ8tTb889q/0GT0KPTCuC
lU2JHDPpyFHktOgDa7UTB2xgwmo0bOTM/xCcGjaArh/tU6mKQGv77rXRo1krfAUYNHig9byhHeos
RJfm3yoZ+czg09asTEEZEBl3dT14Tne/ZpQgLHxJYts4fD5v5GPYuuuQqbx3AH5TFVB1JTI4+vNk
jJ/gVUD3l2vi47orOOmwxSE8vqwUfJphmEZShWG5t+eKvCGRdU6uwWm3g650Ul0K1oTSlFrepDFr
4LUtdUK0Tvrde9RF+VzaRuXHHn+ISh+vN5zVenDW3NnilQZ1/8SA7lFdKwz3AjH34iMCUxhjgiOk
+Q05DVlJFZL7NKSQF4haquq9TMKsRoQ2dgsy8zeLPHG2LuT/YE7u4GUVV/zaV5h290y8dFz5rCC1
KX7U4hEEe3y5AjBAdzW/HmlO8d37tq5waErs6LtE1IqRk9bolS8r5QS8c//1RPI5HrSyIrN7rpVG
qJuI5XhXTJCUD3RwM75ku5E77H6RAtVS9jdmUuuFbo7ObHgD89/8N+AKFWmhJz0LUPPs569a1sly
OQi19Faps+L+mXXb87SAIL8A0Pmys/vEJUtvVP1UW3sny20bNY9YWLzWbIDcLuklyVkmvCJFrZjO
GmnlSSAP9YgGvhTfhPtXhATBv66uB+XtOS5ZmuPbo4eq6FhgI7XFVn/3Uzd/9sxUgZR1nCGnJHuw
9kYKE/uzd76L7Rpil6JkXP+jTF71f/Nftv2WAvzPryJlIp95qXLDTLTuZZW9mV8/2ZnVEQ8SHTc2
9LJLa+93WEpj80QdVg/VFBV4gFimI1Ylndr2Xc7BTX3NqOl8HLEEzkxju0/Nox6SaNWa+gQfqth7
FlPEDjdYYQIrQSL47590ZVHjarzePZXD2wvGZOS5x1ADaCgee/KFLn4VQ7vTEM4Jr+LsWnc3yPx2
m9/SqfVe3ZFoxCC3IbgC0UPfRbSMsb5Pnekd29f38hArtbBNeEhHswEhHHHZyW5pwg/PpE9Yu/jI
IGQ4kAJP/oBaIx5DN14JVJ/qjLmlKoE76V74i1UD/ajz1zP+cYtlYgshtMR8M72j8EQ5jJoliaLd
9OBzskVB5mFRAX9kX7+JzPqbKLWZhvF1Z8AcH+Ozqhehrq9CN0ck/qrFw3pQzbKwxqu4goWTXW42
TE0DmxSk8GNWuUNR9gqLkb0i1oOJeKUHeExzQAD7SWH/Kez/ikXkootelUM1o4oHx3HjWIYMpnvI
cpZIdipmjTFRgBdcFdHiDMTECkAut3cFhzVbUPq0ws3RFer0bKmTvg/lLe/MzvfnUUj5YV1rWnfy
0WXD+e215Wus81atsAWpDBgaLmaxCOnbrv8Pl5k1J2bOeZxZzFH2iJKXSLJ+udrUOCstpZeta/cl
ny3n2JszAdMXPJpH6mxSc7CbxE5lk3zEQ3J3PKQ9M+JsW/2ZMjmzMqNyhSzrmV8C8K7ZCDE2ZDXJ
jkg9RILHka+MwlkDxliez0LcFoLbIZ58O01/6vUbwyp1Xj8t9ImRGX0BWzz0C7AtO1w1E5IVVBks
d2JUbMs9seRWsX9T3QjPxX3y3+BScy8JlmnouaPxd5Fy/evlC0FxSw+sI1LQTb9pjtU9P1h8ihzG
gwJNsli00qILslYJvIkKtKrB3RQuoqPGsTR1eJsQ3D/txYUMLCLMf+BYZRa3ll1uqbdJ0dYX7K13
1WSsA9N4nq+iFP+g1afPyTg84HFZXUzwP89g+IwJ5MqZdmCkbpX/t9jGNoaCbCld/fT52hzEP43D
iH9ACrKtJKLZ7DgfZKlFsW8KnUPcfB6x8hF0GTxQj/rq11y8MQ2Ix06CgtUaNGHLzAOfeNG9fQgJ
tM44H1zi6l4txK5UpuX/3Q4xt6n37gnbv6wTYEsFmqqq9uk6yIWVlJrrad1v6bJCXDv3MNhlYYMd
muKLAVAzz3NYoDUNdSAla9SqOSK6R+OqQptERIjKra1LUSw8RExvqlsdl13wIzsXhXnRt1D9C4sm
BS2NXaW/HK9/zZQ8a2KbxPo4H8UIVfukZSBkoi7jn0I0juOc82U1Za+O3kQv0YIBiC06Z1rK0CZ2
pwIs6QHDpPpJy0+eu5JQnSydgvVGROzMa/eRkP6M5Omwf2Sapj9lj/8JddbDc5BQSmf9xFGHopVZ
SC7sdIMtMnMnP8+ym2hOqya7IIodHu7NMNqrS0QhMoKwAbtdUOUFskvXvKqhoTm5EpYMWoB0umzi
wD5d8pN3GU7fyWC7M8Zw5JpCioBZMOOlAU/KOeRtvep3X2c9A3xLMdESLk1FALlbSAujvBxXssg7
wN8Ha59HhgfTnJ1RP4i3xYPIEikf84JKrg6up3c7em//m4CCp8FYQ5G0w4RcCMWxCcUN6yb9IqNZ
tC/AmgZNUIwOqADfvWxFr1AACsm3ylNOZnnw256dVJJ9+ZSGFcqIAk+/qyEtmUWvSJX2ha/3C/+U
8pmuSfw0bOAEsJ1TuvHq1mg/ztbGuS+6EswE+1Kn0HYr2F4lyVC5SnntiiD64NGTosMcGdwp7KK5
g2xSsxHoPfOkkzH4lMWQ8mFv8LUqqjLQChVAp63EUdHbBTQCiNAonIxEw/O112dmpjSIk5rHjcVa
fDbdMzbvuZWD68DdzU8pQc/a/KQky53B2zwOsZRfxxWYiJJ4AHoSnlodCEfT3Kq2K/VN7/TmwiiD
9XATxcUmbbIYBqmG19FLWhslGTdTF7WMgJNdMxsX1ChBZZZO+W2T+DkzLs6o7CJcKxdD7vGLe9na
/tO+s9w9v60qgIkJctVyJgrw7+imjSb4C6kzaE9UeMJo5gsbMyCCEMlsbI8KUweD+Wy8gghKb6Ld
xTl5uZOTS4mtwFBwLMnuE8OnAQi7NY5KR5c7ksDZav1RgMhnPRTo6N4yBkjIGyuYH7bYgQWQ//1k
RwagysDt/c4meXD/FGsvq5JhWEGZW087vv5qbK4/ces9U4IkO20p1lRD+SLr/QCT6ZACfyKLQKHl
VVeXYWhXFuIu5S+3PXG6v/Z4iIXcLz9PbcOeSVkbV/ZxzL2A/zXPsGwt7tSfu6DR6e4Oacid0aNB
V1VM16wH5OgLkWkW1AeQX3w6A3uzpgruvZtcVNN7veJCTs0jwEtt5nzr3GnOSIjKUiHmU8TXsVVn
6iZqicimOnCMO4b48EtfDgtqMVjtAXQ2l3lN4O6zkuMryK9T8kXS8puSmipga2QEv/tUbY/0ldvx
laMxqDB058n1WUREMN+lBUqgIxi/g1rdHvOdhYAbSlswPXw1xqQ19+2/WM76xlDBl0jb6qE4lPj2
ieQm+FbE75JFg08Rc4G5sQojtNbgbXnVHpxmlIDztMfj1D7+O9pa7COlUq94LmMOWs8dzk5v6nPm
k8hALUXb+MiuQaGp2QmvudQlql9ooyGFgGM1wns1BkxcZU4rqK2y+hWPhmubnjXWa7wOJ0mIOIkD
STCaGrkzGpYrk12VSRPfi4rreBb7iqg5CxJX9B3+g2axIpFUnZ+ceD0wwI9+wRTWYIflQr2ndcHA
pa/Ig6URt/BL6Q0UCijMtyMDI7XPr4BiUJThZwYljmZWHylg3SC8I6Buna6zL7e6rsT+WZc5fg9+
uBUgc7BTJU8dCYdwR0tE+KjEn+v+BPTbc2/ZE5WRegUvmLlA+ANLh9ZBsGQj9TEhFYssldjhCs1X
gLIjniezexd4iIttgOoV4UhhwL8ryPcYsszWudDo6N5QkpB2hsBbzCmW8g8jY87VtqJU/Xagu4Oj
yUyRZlbilg2wN1JeVe1g14EYN4Xb/OSqDeAZD8vH6Suy42YJx8IHsaE9NqvXm5wzSdXJlJANqRN9
uT353OX3UhR6ldRvZAeyeGsWHy6qwGvN+buK8cW8jZ5ShnDarpeIxKyyTQWLK8ZXbAx1TqCSyi8s
LU/O42HSY9XOn35xIdkcM4p1uhN2i10YIBIad3ikjj+/XD6yX+wD+6bDoHRii86IohRCCEsQ9w5u
B2xYFu0D+Rt/AEwTW6E4ai6D6+CvsOeAnk31otyg8TNfrDJUPcYSug4xzlmN72OeW9NBlNUA5pj9
ts2jEbPMqtNJp2FaMM08jK4cB605jzFHl4RGkGbWXsetTZ/ct64tSNjQLMUo5WjLn6KwJuol7mtb
AcsN1aYh/J5nT4uR4EB6w9gcGS6zCvdoXDG9gn2Guclc7e/jacY46DpPP9dJAYUfC7IEJxmTKtoq
lwO+c5LffVJabJK8b2bARW97drITUfstnDPKCCZMZtOXR3OcPKI2hKhVND284jF02KJvBDlfDfx1
tdosb2rCNCXa+nxhQqTJ9e2vY5vTJO4LmL/TLg54aVCmvDqXWs7W5SoZp3YKSfeUS0mdlbZy7ijC
vmviqIeU7BbcBqQgHSYLiRW5vToEWQ2iCQ0bwKq6326OqLqPO/TmKO7GNq6/iBtq8hD1qxcYOCRz
0+i8dht2l739p3iE2ucExN9QN40D54sg3YAe4yOgN53maThFPJHUIpGPi1hD4JQJn0zxZAUwNdBD
OSlgLWkKsyjVHQxd2r0Gj9e0UUHq+KTPAb+Iwdgz63frxqSKygFR4Lw/tWSnSPEZfv/BQynPtlJB
PbuiGGTk0TWPNtUThrhnD04z2FpaNCOhtDLayJCHS8fWu3aPyhQ8a2mNnAvYMPBQLjE7ooTGZI0k
RDAVxK+vKuesMSp9owHGm/tlQ+6GgcxsYM1pvJ1Db5zia/cOdMAdJPOtJGFn5QEmXtYcr5WFlrnU
Kwgu4dVPFcbVRVJdC5RKC0UGvueylvpANA0TJw3gGxRKrPOs8zcZA5OcxjKUvo752G+Ks36ZSoBS
PnWnot9cOCMn1oWOgic4P+E0ElTHa9lEs7wY3oWxbOdVV1yKD0EvBUUL50b3ygK7fB1VZmw/3zw5
RDvdCNnda0yHcgMu5dYzc0tn4WNSpgziwrjk2PzjWqvXp9AgyM9cWnISGZJk/OIXeZmzylB2as9t
aUH2Nix88MM2a3SlFhTwfcjT38aS2yuTvi0wEbKybPoQCLEeDanIsY5ZIOsEChM/NWirHZG7tu9V
w62nrzw4jRNVCDoiS+q2zoOB0GsfZrUhDxJY1eELYbADzIUthr6jyCwzmqchMcD0T+cLKYac24TY
lFXwEcn5dtxOuThiCYKtZ6o1kR0XxG2c9uw/4Vp55aYwkeqW0Ivnu2E7EURnoTUVQU0a87qirazD
WRfqIpRez/2Erb34TdEkIfqv4XhRGjZ7qEqUot5C2WTHw2nhIBcw6ZQ9x6lp8xvtmtxS5NJ/juSX
Q611tyUWhMjUg09pwQQOlzAG5CoJocOzygb+dJzI9tnaoDTR7/gGSh2QtQNbsni2wN+xxSb43RpV
1IkBTYP9E4UrRgNrt2DIhintcK4oiba7VPkdV9fpxrZIbLYuFS+KrCsY8gHflLdfH0n/fkmbkz/V
iSOVRsADF20MqTenP6qr5Kk6Wy2cQKKS6tqIad4wjr4ytFGU/ML7OSq139CHCF9QGAEXhVG47OAa
pIuu8a9vcIVAHG2XWmO0kGIfxX3BTp9ET7Me/yruw6XFVDBOB9gN5MAqDbCuHq73Tbrk0YhqZKYm
AlcRbaZd2Ya2wJgCLS8DXKsR5110zb9ZO557jFwvGWEreLupsReKr4g7wI4EnosH1W1ZUTjyK/Dd
IX/051OQn3Acst8D6f0DkS3x9YMQY6hyNozWoODdiUoFm/eVgknXylB0LTA7HGjgTyudMpOHoSL7
jcEgHYKeVkbM6xGgjxiqyvXkHSKyjaNgalYEjGugoUQ8cPwAgqh0/OpR0y//xp3+sFTio4ET8IiD
Z+I7K57Tczep9wc8qtDi8EZSmv2E5aJ6rCMKeT7IaaritHesnPAr9ow3912XpSYU2CAsl+lObAFM
m07N659YHHActCJ07pwPJcFOtptW+B/lEuRXOjYzia9Jmo17tAr4D32HWzaA8IaYgS8fVwOOmm0j
pAev7vSvVRGtBc/0jbtF97WehlzsRiJWO93snSdUM0z9wWjK3zFrXyYZNJJTFclqAXeQu1n183CU
jIaE6LPHWAbUrQD2SDFtaxz65jh8Wn+mybBky4iLDfrHixMGkrSQQvhBAvNZ3jeMjg1EvqoJoyuU
JWnlF0aDBUJYf95Q3RhqiVw9dXXGUo8eo9gmnc6xjB/5MEHX4GzV/XldCZykLI0mGfXs7Zcp7ofE
La0iJM8yJDUobzCEk1roo3zvltixVo/Rg4fbh8f+Xy1ila+tf0FVHW0MwERH/j7EbFIM+rUnoChn
ne388ffXb+g5ZPujsSUM76XzCKfe/2k55SU4XR5BT51NSmcmzMlg9ovrf+85uUL5I80uZfJoAVcX
Ry6AhEBYNPQNDpHANlCkBMzUhPvLe9dOOvYEwksQX+XfhNQai1T4y56sP9hZWMeXR33S2ZDyq4GP
Yiw+yTnlESZZZTK9poVLPurf5JFqoydEueiWKCNAneBQUfOA54pdE6xk9hIedNCnPk0qXTNVul75
TCbU8DC9tLlGthkVsI+J1bgn/jQPHVbUbPyTJGgbaZ+jQ4qS3QEL8HN21KtwAVl0k7G8UiZ/sE5W
RBHqRBxTL61MQbPnY0DHnQ2D9EsJobBJOmF7D1PSd+tHKSfIIvPjUAOlzj3x3TuQnLz+cbmlh7R2
kILg2x0RLLP+L6SfQbhcFDn3I/vQjqA6itP2xQRzTA0wKUKgjMTGILD9un6Su0nJMXlmgMT7D8OK
ldMu6xgJa/EcR9gL5PMinJE+w63j/Anwk8MNaHCnnTfLHGo/Txd/9jgK2QbTaoQoQLq/WBNeqChW
LuwMGBBQhwn3+KKeoNq+qRHXMzvQmIYrNbR2yV4EcI9PESL90Elz/CzZbb6CnTtj5pLVA1cYzAmK
1O723XAafrdM27nMkJF5MF07kJFeLpaNfJPd6zqlBHHTcRfcocmtTO/kk1bfLRgqtCAuTHrftTCP
u4tvZHW06oHCXMBCRZw5Um6b7YlP7TWxATJaPjs9V+kKs43ctZfbgQAU/4AGHEu7fFd2dhIjYwZW
4aoBVEAEppmToSzNVI6st0M31aizGQusC3OJW9GqxSlkrsGHlFX/Eku13ZXdSQe5rCmIJ/QTRDpx
PCMaYeqpLWSrMq9qE+V+Z2KYFtuUYzw5yhTsvQ4W0ENMNYYsT+MYZsp3V7dq+lb+GJq4n6ciMn0H
OYbWDp6PxsZju92NptCDZLl0XUJQtjAaaK4keLlaOMZ6FRs0RStAmBzUhXXQIseYpSvVqCjgPP0g
c1uRMASiG18L8Qt1sThOPrGEzDaD9VKdYLXv4x+GcKhciOiRr2oMFP6bZYjbvk4rsbc+Z1INWKbG
XDDy2M4jP8GM+s0R2/8cNra/FYdaRbOKlkWIzbmk0Lho7Jf0BAxaedM/rGS/xVjTB/hJBHWb8u5h
N9W6VjCtxAalSG2xyC1C6UhWvozJwkSYfU398FB3TZzi5fxb2qoeu3ctm6Avf0o1xsBL5Ff38bCw
iu2YeYv0v2350Hx31bDi18b9zntWLLy+WzWQ4X2nWZtNWf1jjTZ+endsrEbkS+AYB22+UdC2wgXS
De6pWPZpTUtUXcAKS9IhQgYxVOB508jt55uyl3cctU27QUg1xPWDhrkIWA+WpKwieyCdMfxQnO1Y
H10YFMr1Dk7E7Y5HhtsoILlh35AbdgbEkx8STRKfwLIep/+bRG4tRvphgpNXNmGiQaFGcVwhjjE+
Yc9Vq3e+dUTUDEb80cyV2IPbLq56OYYk3m2tGBdVjGYYA13CdgSqb9oQlefkGNPF4i09lus7SFSO
KRcniHihfx7yW9qER1H42AMYAhTQbjl0kSoDpdicyEw3AJ9EJN65WMDPjKkntKzGeb4jU0dvvhVg
NVT9uzE5WEU9NSmGiH8g1qDwmxdtPvW/ugOmrohRoA2Re7+tF8SIyLUMjUAFtHzaIgMuLgGhbxZF
WDxjj6Mc4Zt48CZvxY1Z8S1V2JPe6C/MmIybxxZx2rIPyGXpjHMYguDU9hQs66w7yWMqlvaoKF6I
56EBsXWq+72LwhWU0QfQ+S3QyRpPQOaCfFI17R9yW1gD1H2dMtKpGe0gT9Cff55BdlYKOu8aYqPn
8o9sODl2idx/NNghL+tbIzJ6szVep1Vm+lnmbLY11vH0EsnzxHM5dyoZUjy5217HC8BP4VOW86kI
vAP7LccoF+RkDNUuGF5ohncaCvxUVkVGi077JxxOYTKmGg+HfrMZH0UDYSeoTAW+Zjd0790q6nJz
n2KRhGlc+KKs+8fueCULI9vtocSk19txwlaWw9RcEDoff+OuhKJFYz9q9KQLTiF076W0hSkIQjYv
9ZqX6gAwTbAcptaRmOKnNEgI0ELWJHkeR9ClLJXgpx0XIggpgBFYs4kRYYkMGsPTTfNS3j956lzZ
JyUXjHYhO+cP3xHQxJUXfqBP8MRf8eA9FKAG79D8Z3/ux/pTuWZaHPlFh6BdPBiXVxf5/Zs+TpUG
5ywfV/yFiaxjJDmjWMzeO1XMOCgM7o3cW7v9V3yhdoazchPmp+8b4dGdk9mYKCjpxGRWWXwvsI4/
CH0sNKwShOXRLCl+VBpDmLh8HPVHtyyKRezR5Oo5vpbbOJKgggpv0wEKOTaTLY9A3SakW7s7Ly8t
j5p+f2D7PlmHT6rzXgYVlcG9FQyX8ymcVGEGn2jgR4aE3KE54rmTY8F4iHa2+ZEO3+5ox8VinpZn
lKCCVi13iiH6MRnqajN67wub794/XRPVcSRnWWRwbIsg2Tx4RmVDjwqX2ghpIGPJfHyAQ07pKcX7
lo7+E/R7IgzkODyomWK+TD38thaAuRdlrKw2DzBdZTe8kuPyZMSgK6OnZhMtgHHJOItDxNlxANoo
2IlpbA8IsIXAywgpWg1FEJIJPVHvxRUB2cl4WjmVzsBJfSFQoI548hNXQPTE1421MNpodq2QcM4/
D1HgSMmsn00Dj0ZNI36WzEHQcUQAdcz5jcnUBlyKFaUP4XpJlVopbvV8O/iTB+Ly+XioRUjDhMkL
XqZFhCz3RD+nMw8NtIFrMAGrt0ihiV4xvgmBHoc+1lhs1fPUffmfppZPHIrwKzpVcycrvi2UmWHs
cTp/Lb1I4jJwH1+vm4V7tpIqk+992+QbzijHfwzsVN7/YEZuFf0TdW8IMgrgXPBNraPQFEKhIDF9
8BpP5tNjD3lJU+sYnFqXzuu94V6TJI08BzwLM8oVFxO9LqcWT71Iy9lpoFOHaFTZtD7I2Y20XeQ1
9mgDHDjFvBS1vr84z5SC6h7KsF6Jt90HnsPrCKmZGVNnGB51sZf60+X7zqb5GWVv583e81J/ROrb
aHq2nipA//flecW9P+4l29c7dGIKCMRO/63hxHSAcxU3zLy3usBRlcIuezGdFZe/dkY0zmr3L1fx
lvcbyqpRYnSCCFOOf9zzs+MK9bHaeuuNjyqq9rht1sygf5IchcUzX6N+ONV6ZFPVa7lf+MQ/dcik
STMzfIicKuEPuP94I8tGBbtIgDEOrDkvT4T3K8sygx3p8ycDps8j6rHm5lF5KTq88DMkQRGRXk3l
nO0cnQuANIievb5jZXuSW/v9hC3MLh3vvFv+cp52dv3p0VdtJtwpvxxk5jtH20BiwtfDkcfL+z/y
90dryzj7Gwt2NED7KcBVeU/BPxbaxPnvXeWiPk6Rb9ZIDlxSGSHTjP+yEs+4ExuRtEx8QjE5IiyL
3CP+3sObal4YaMnvZxgLK1K6K4YxbqGgbVHHZ7rK4C7xoAY88uAC+Ul+MuAxv43NIfsLzd8kd6Zb
7jSYs8EUKSJVyiiSWlqpo9qm30NTK5fR2vrhI1cHbdw39FbolABDxeeysNGSTmYJDeUvFDsKJYlr
fjHJ8yywysZl7hjCrECHg+a1zsTYOLYjkwAevDDFylU9j4CzHEDnJfCZU29lO3SPUJfGQagt2rJT
LjUCASIXLjzT1M6BVf5s5NXCekYkVc2OsqhH2Jr9PqhonARdhSpM0rS+475uJWmaMTYRvkdj5sqQ
Uxuz6H4NMSfJAG4Pa9B0Fy+9G3YoAcuPFVBNFs+h/KRm0Yk15CowVYsgXZKgyzy0A/oYVtEIJ080
Yb4x9jlr4RIdddECRP49DmsI8hHlteocayNZFGvSjsrIG5saCpZ8SyL97oibCAYIgIOCmGpVozKJ
aPlSJqV4iYsYi5awXv3LCs86/25qYUytmb0HPfq3jarA3INJudPjugaV+tQ1lMP7SJHVcTLdXhgz
iTzg1qmdYKc0bRr79ARxj/KqkNW/K9ghCx6TyalgqM1Bce40ZqLpj3LJ6SNInYlZXvXKe70V3Y1g
hNe0PAX/FwZGb0LMVVDRQy782Ixs6gTJ3mXwePS3M+JvKHr6n8IeLMhSk5wb8P1/Zl3BEaieHfQF
zt+RP2K2vg0sAxm/zVnC/zcdwAt4ZrjiSxb0oDZv8xa7zWp9lA4iACJBoo+1qhq3H1u+NrluyFDn
rER2sRa1Feu/c49Dw065Ml6S4faaZlXESZQaA3hnmdIRlp3qtAJREu9KP/Pu7whRk2gx55+u5wMQ
16j4UDkg2/TQF2TIL2a6UslZxqDv73hpdHp82SwojwsIErySTE29BZ26HtDr5B9tFYD65yLVP9yX
Vwqc7vJqgXzbQUxNppwpv8m4DxnH/ZYrYZAhH0sN683LQAu7tNdU4bZuDH8RVFJo/m2bvSraZhD5
VWeNIBt96plwvb7pCxefQm1yd4Ma1Y2UiFjIWGeOrrd5lZJNcv03DZz/T1f8XeBH34mkoJJLd16T
O8KpAMu2tmFkUDGXDTIhOEwFxDlWPSjFT+5yxTrE15/gwchvyTE9B8576H89/T9BbHIbz4pjjwZT
5KT17yVIK/1t4eAEtcnqUOkLlGaw7d+Jsgo0CKj0iQ/pF9a4yGswtRvG21dse6QT1y2vGqgCJBAY
7HAGhsu5toLV6KVcEF49u6CHR0AqP4cdoj5Q3Er32lo2bVDVlkpLz0beEa4ACBecVoCEMy9EWHcZ
A4kqSFV5F3136bkHDd/JsibGdhod4AKVb8mDVDMAtR2Qo0MDsVzE60fZcuq7mWFWwgEpPjSEqoAY
qqTRddDt5s87uu44tXlA02TsaEwrdvJxx29vCFNcYhIfjstpy0Q3I0r0Uj5kzSOAEGXW2hGFHM3e
cpjwjipplEfWY0+wob1rCtofv9RxCAVIDZa1b04HIVRtuMTSXKaLnYMI28j/BoB4u9gsogpw/i+m
9RXwpbDOgHreH5Nsnml42bywuhD3XDZd6eAuTz/xiqWBe/SdWCqeCYDqM8dN/Zo9ajG2NgH/SePp
rs7F0yfJgbxv8eZ00TSk4yANeb03LusJEXQ8QnCW+htKMoDsi3mv9k6AvUn+BTiOi6n7xhn9ZOSv
pfC1+cwY8COyqM1w9WK0ph7tURYWWIEhdzAgM7bxRyKxOEYRs70oo7sYp7BKgNtSRUQxOIOtU478
YTGnAH7sYTFElD7pxwlmbOIo8Ddnz+hLFW2qO8jvTPzWlq4mWARs3zcxFr2cHtAF/morqxg72sxj
Y6wHNZizLRlwIngTguZ0+3JTUZeqt/QRBTSoLmtac+Vtc+6ySyMDbDmGF8aX0ZhiaKRrUECFWeNY
5lGo4x9yqRTxX2EYDEQBf4Zl4LUUNFe6bjwMObTNUVe75RFLAxy8o4UmvGhFH6sdmlYb4sWhHXOl
BP2h0CwPtUorwcCIvIU/6G/xieBWkU7rwhZQMtP2KolXF8cLa5fN2zpoxql2HvZsb4ysvLqZzLsH
988wt4wB1PiHoBLQB7xyFSFHjKFrZxO5T56RpLS1MLgbDdU2LnejZN9ZWZ3mNm7NAANLxRqXPbFu
/NF1Il7533i+Boh+jOxh6i/qlJz4ey2GYRKGlP0SfOCOcmyf0Itc9JW6IeQYGqDhUqM/MS00NFPn
S/FJppnvD2yz+UZzqugGlupqI0294cTQ9l3ZxPatuU/B+QSBAV/YS9iiipjaA7qvkHXD3SMvQo5x
ZIQylF+j/YvDIT16XL/6ltyXvHrGZNSHLWgPYEYSMGN3QWFk9+9IPQvKKDoHH++0xYO/dQ6RtCxH
o3KFpyxeGkYOWNOrlNhUNlGvPFS6MwiLlaBDUj9BEfLfl1Uuix9sFuZ+uTt4teJeq6PADc968/SA
eopHAliCtZbhW83ilLY4Qdo66YusgUfS+ky4h3KWTmHaG4tq55spR2iBS1Htht4PC7c4K86THOfS
wMlyGszRoQv3h4kku88RJuwzSwAaqFPHDeLa/ofguaHwJpMrabb098H4DD6c2F1TnPEhy4fnEU19
+K1LihUAWSaW4S4vyr64/ECIYP8b3qNJCgqFFt3jqRkDUW7L5/PHntMr8wsvjwPpzUXRuBFq8zUL
pLF6fy8T3cbPzD9MeA4FVwp57WwoGDRh9ao/mvP7pbY/dTiD0c2onpO1woXbAWO3CCY06bVVAsIL
6AthYZX2GDx4zk3LiU9W3E7qWJTM3rq8LMCd/rUBEIA6TK8G50yA8IU4XshjgWaNjhEyS7YhrV1g
mTHHFO5auVN2vTvUr1ri8GfuDGpHunnQ3qVqFtge3Pmhm7lEFI2DeQyZyHZygTzOwGtJ9VTRFGXl
av+ndh0LJl1CJv1evtnZ/f36qSHJz3XRjOQW5uy6gT7bvSQAO5K0LV4jnbd4RLx3mbk6kep1N5Do
NBUFY3dLzfrIlJmTNl2j64+5CQr8JeTghRal5OnhFxVByo82xyN0kLNh01cN3Aq2zFX9J5CZ2bJ4
RwtyG9gcABoNaj1HeNnlXU8M/oGWnMPgVLkeXTFSM69I57RFzrXkPtLXU6yiEIFLg8hpmyuc6HPY
f0YHcFeTkrHdxxMk85FBRi/xA/Ew8/uLvKCmu0yMqV9qab4nXHbLKMgMHuydxczlZmfj3ENN4bEZ
R7tKmI+OUm+a66JxNSmuUMcKRS+xmbCqTdE3B3eESI/6BqHcHQX+4zhpWsCzaw3ccR9XpZ7pdd56
bhiJCs3ioiK8iTXZ0D0ihrvcQH1AKO+y6KFdk+QR0Zbz5qyV/0Qe7pv8UiwKZfqN4HcKmJTJNyx2
MEO0f1F1xJL+D54wSRw7vCrB4k4WK2fx92/7tXJaOKf3IUIWUEtFpVKEuK5WeeTniY5aAnI7KJDN
b/i5wcKPRI/h3UmDcoBk5H0la0m08kScNDm2m9dV4B6fbkj2OlI4/hqeenVscb68+t9FhEu6HT59
QssFOuwnh7u0+h4pJAOK0M+1tFlNNFFRDPSHTkpd2+7A/e55cXl1TQ5nEra6cwHeq6JhOZ2WDTnt
nu/Qat/5XgHPeU+OonpzhbNYg/B9BM/w+Wl6CbRbNQz2fj+DAt9/QJyV5rlNcflKAvqGPk8nfx3Y
Uph6IQ14kGn7TEYJtBwueN1AA745xLcsmP6NdS03C68m/rTJU2TP759U91mNvNwMVay2I2TybHlB
1kK5SnPYfXwRl4xyUHGEi7rpA0RZT8Z8WmvJhuzpKlT/VxOWTFeRNDlWF6UmauqTnde8zPc1dWhS
KvU8Wc2sM6r5jeDmTS7cVDzFjqXdUXiGA3JjusOWskHri0GCJkCp6i23qavxnwVrY6CTfHmvvBwb
w2McmfqXOpsuWOzLvHD8BR13OdspkTp+sz+sBiz9FrTaoGszQgul5fzKnzHQjimU8vQHQQlkfR5W
G+qxynZATYUimyqxyraJkVdAuVREA4FELwnhysANY3kOowbKmDfIZWzixiThK0hjt3DSlDFHcHu2
1hOumgQPQaQGoXCjsCjDKSJ599maR1QoL2zbWNbSm1nCAe0V7A1fvr+scZahQ+nkicc747Rb2lfD
R79xXczzr9GfrMI8mRCVKwOYqmhDRxZOaPU59SymIgbvTo+CMy6UOT+tkkt/bSidBDI6mUPRxrs+
R2VDS57eSnUt2DAqlbQDSKi5+y9T4YipxDNvoBQoPKHHPCReWojdxIys/7GwYvKO7+84xgJLhHHz
tVHwQJOnqLwEoxhvsGgqpXCdPDREF3+SbAwu888jrvlvLd0cNPREgRJ/eg0JauY0Z6U3jUl+78EG
3nnPlApYg57Pq8LZfDDMdm6s3hAiIgBG6go0gCIBXJ43ZEI+WkMY7lm6N0Ag6HGAZ/dXhycmaPcd
ygB7Mskk7jW+YVT4ASI87G3+qLLHBfAIo5I9CH57Fe3NZVL7BoqgC9/mB2/67qIWDS4ra5Un2MRU
cGAD/+kA8BYVFAV1MrNVcbF7aP0Q5NdAyeRi2BBzzKmq4k8UECCU7dEPIYuu4cxFoIan5m4Lkprm
oAmtzK8eqj9fHPonslnGtmb7/KMTyAVpEAKmzJP0pISBeq8CajOb2Y9ku32bMG+pNiXcI+RyfN3T
qczExvbBNtYDBisUmAsPYSgGelYfFH7XPpo9LSb0HVbrWQBsgTI3w6BXQyiWqkUGvhMoHJqrII5t
2k1GqM8tF2MUTaXkMCBSWWGkF7LhipvBDIDb3fIm9XF4x7hBKoQu9UWoUI6pxGKmcD/WxBlGsOSf
K0oBwggjZeam8qSK6mNMAVRUbBlbj8LN1BvqdzHbyvLVXZnX0sasAakBLwNm0xB2IZVDpSL0PNje
eodQ1LQMfxSibAut9L4NBUBS/jjKPvxCXWOAG847TsUAeE9rbaQ9FFNcC4b+C0P21psfIgk/QoTa
csGj5Sca+NFH8x8/q2BNP5Sc6JrQk1pVNAzeI7LElRNQ7/fDRfMuA5Px4+HN4ivgn0DmIuEbCkyy
uhuvsQZMaBd1GzaZdm0W20e1uD4hiSlTiPNC2DKlcJ18U0Us4hctgZljfXReNoexAcOKNfjc4gY0
tDXtUVwbGJdsmoj33UwbHOIPGfRDXxhW5c2k52kh8PO/XZKsYluLKhi+VT7Abk1QeMDgtvX6lI17
pUUYV06b3FaqyUfCDwM1MXPE9fCrLw9IfZY46A/HPt292SVoJoA2LMzPYoeEZME5OX4prDYOoeH6
K8YnoMTBknSNdIuYl+NkRhnkH0w1HN8V8DBlvq+PTRZGmqtRH+f300f7FeY/d0wgIEp8yNAtDR89
dZ89A6rwIwWmQ4FgxwN5eO4Nv0Zp8yY/JNIM2ctLVTRa7x3BBxDmcjSvBet03iHW8hz0BvkBzrkP
h9d4s20Qq53k1WdBjlkWQ7myJJUB08P384aG3h3444cY4AoSz9U6HTprduDT0652ZwXAW01VtJ3W
HwtTJijzRKiVY76VdTRZgx0BNyNXCiTffAAk1Y8PWb7NIfGr8mLBw6TexQlHNpkKGbzIKe+xDUWo
HzG71A1rMqL8fJXizhcf63x5MotlJUUgPIYC3uSy1W/6VyepOLsNywju+hBj/pNC4RRTT0dromWH
QsNkPz83OWl3X6Zho+BjKV80xrs+IQuNp8jLvmMj5aUD3ZJjtrcVYl/JUPXha/katio7CYkLq3ET
pjroGFj0N/i3gjtBmdxsAKK60zndOD8D/jvfouBpI01WMm6Sd8oouuVqHgY8018Fw5zgvNvjXKmU
7j95FLPwf1LkYZtRmr5Ws8TGa1Yrrx63jQFi7br0OCBcBznxXQo6RdqUkSB1lFP8jWLRjlArJFzU
mnHbRdU//F6mG+MlhCAKBRA8Kp+G3AZAWRQfHsOf8ogho9fz9T8pO5xSKYYxRSIZUQiMIwuFn3c2
lsWPIqN7fTJlb7OHDyQow458eIqqxlGOR2943TV9PisbZdF/X2mulTAvdnX3Lj4jRfNs1uErLrVe
6HH8dcPiRu78gXvXqBdyNtLrfQCIGfoZSB8kWPnlneTxJVxYch/pZh9UkK58GSD7tPz97Y4RaM4D
VI+2KvTLrFXrBWwWqjLk/Zb6s4Hbop98II74rKOcz2AkN+bI7jlgf4ID7gTBbrSyJAqyf9zAPlzP
sTSqg9+PMMzJW81bedegGVUiLS+G5PG3R57tqPMQu6FSKI77OXgceEGSNB9WAdUhln3o0hZmaOXy
0WaDK2L4Pc4yl0doeftuFafUlwtE9C/Dv3Oyil0Igj8u/eSHRyLdD2LLR+zY/KtK/hnI/mJrRPL0
ydZpdkMye+3l4LtNXUtGl5dZtMD/5dEFObxYh9rg8YQBHZ9pmfpvCQ1CTASfktDY825z5VxJc/an
TB15nXwf5PDjLOe9FURLbXesWQVm7J0n9xKh4r6G3WH4wlP98PI/2EEWwX2eplv5PiVnHVRwN63K
SbQR4UK/x833DSDNB7HqflzGJHEfU9aFv5CUI8kc3NXotuzUjjF48J4K6Y+u4JvnNX99aPOwIWje
B7jMitQWsyiU93BWD8O6XYSSd6TeuYuu0/TpmkbGCNj917LzD1Tzo5P9RM6N1I9sC+GSXpaOAjMz
N1LPP/j+uq/S2clBzTOlkw40yYIBwzCQTCIAXPzfAnPwp8bpf4LOhVtBfhy8qhFvyg2b5xf+B8M5
nJkCDXsdGxYg6Ri16deZPZsMbp77NZCd5AYtlh2MvTkj76uRR9YNhcaPSdEpu77V1Ey49gjWFm5g
kdig9Pn68n8Rh/mTLIhgX6LdmZNIqkq3PrescvJn3z9Fj2pxPGFEJQlVNnNxNOdxMn32EKCDGh4Q
ctF3e6Y0RWgUgIc9tdPZBoAK3JMcScT/tItL9lrMSgAgcbHelKjz/7Gl2l9NWtrlQYbyeVFzqobh
yrjMTnjUCQ3SeRRYJ+o1uVa3q0TEsvDCH0/lJqvKiTDZPoDv+p56Delx0erIGZ4THMJtVEwrvJPD
OuW7el50xFcPV8EE09X+CeSCB/ZgZ0NF0T1Nb39wHb3uwlqXjeA6e4VkbayEK6lqwi3cshov/Qv9
fffvlvGesrWieiDNN2/o5vGLp1jpuSQdXgFP4YXke/e8EHHKnz0UNgqyROusdPQhSru6wnGjEZMB
7YALC+hPf+ZNMPdw1RGICkD7j5xdIvgr/AoXqf3qv8XSHd9/gLXxro7KdV79oQWpoSftBrwSwJNq
nCCwfl0qGq5h08P7Rd4/7oWf9IHrMsoR0sjh9vj9uz4/8Ad1WHPZHXm4e8l2PFSi0Eg9W/6EnqTP
uTNJzCkvaW+tSiszk/MAjjBgJqqPiqJ+/bEzxNUmOymmOGHmArOUHDQYZeLuPExRgii5WNCP6h9s
1RVjKX//U1q2D/ZSiLzqtjmjF8qs3QkWUPwAsgeImdPR+Q1npouk0ya8jhoLxkR6YPRrT3DXw65t
/yWzCXv9vBx7DMhlNahrB4QOhVZnpIZST89OHDbO3jT6IZYB6snMjtXlYaeIvHJxw0Wu1ju0bFLr
5otYRoDNHE15hzqiii7GRt4WVmumRs2Q1MdUgitsMUvYR8O+RfTpLOzXlczxBpIEvMBcY1BEyPc/
C67Mmr+yPxmBGyPdN6UH4BO7RKOzMpe66mVS9jlNfjbtwSS5M9gOAUG1iQxJAVajTozfsnsRCOSJ
a+JuMRBj6gQDFUMXtXcel2BIFunbmeRbJ/RijgjqEKANObMgpV6egoKUW/Om8w76rE3LdCB0cg8G
FEHc3YBMqOcj1r91mMWGF0Q/9lD9HLdR+YmmeWf5DpMvVKUD+ajc8AaFFgANVtYfbxLD3lMC039z
83LuTvcl7knRCfSqsrZBSFj2GFPzML2cl5g0kc53tRQscLl0oPlmg6XN+nNsyGcbRneFnBKLx7qJ
mQdcPXfBCx+EKpBfHPo57QsLt1vwuSY/3hAdte0FW4t+u3nHKGnu2ZQ2KIR4X1x5/k9xfHEoCOk+
Edwm4/7XkxL/NMRjwrVS9x+6lAf6T+6wExbv8n8Q6kRhsZoeUocW6PdnfPMqztNNeUHGaFyNKM3w
XKrDTTP7WXzqApME4BTeTplkk7/OU0pOJlf/Eelay7RrJANj7G/CTcxXQChHJCrTULtZhG57AA6j
vPx4ZVU2K8Fxa8ndGBHREupq0e93Y6he8UNqc6aEus1pW4OaEftiRx7iNnAHh47VQvKY865cyT3E
GM+OB5XYwp3163DnNpERQqzgr2zwKUTtt/GWVU4yCcgR48gIqXeYxbAfb+Qhg+pcN2A8/Z7mVWOX
89KC+wtQQdvsi0HFys6fSA/J935eSowTQGxlzPZ+4XicHqJRnGSxYVezMTzzkQZ6XrSO98vD8RFP
YPw2bKXE8cVlGKuL5ZJoiHqkBj3jyr71rnMhq8AT0ysfMuJO1FKNfAS4ClXqLetDqxdCrfDONtpk
RFJuEk7J3/nh06LuMb8RbuO98DNzM+CQu9Fm8kDYX/O7DQchbO5I9GP9MAFEkCE+0hpMeMx/deBW
vw2+TFLMICO3BT4lOJzPsIHxuzyLDnIFblsRx4BGjsfQHF1hTWB487jRCRnBzykznAbnISHakP8z
dIQupG48V45iD7OzG9i0Tu39qH5gPZUQJEEUo2cGTOnY890Dm9viqPuZyyCHl0JE+WCX3qkglOF5
F4tAXjn3vgb9SxzOojPxXItmHnlFyoIMYx2e/BrcC1IdG49ItqyQznOwjLTpigutkqwm+1iNU8U2
3Z3GoQcc1TqTdwOWDZvEcdIj6BZ5I0fsTnoqXoFzJ++skXkTBx/Lqepq18m//w4nY9xY8OhSBGcd
gnioSDEobNpKUDoIf023SvB5L56L80v4/Qu4FzcvtzH7SJP75uOtE5Cd9qZmyCzzo2YSJWoTk9as
P2jPMC6kDwPPlkrX32wp98nNFGizfDCzFoT/QRAM8RLmGoUzQT4GpEZPqxkF8fWeCTYhTosQDAv1
x0TSE21UhgFT/z9BlYUny2gb5wB3BVt/7p2ne9elvR7EB3xX/BZhKciVGPevIFTMuDuTTnNTsVDk
MaUoSEENF6qhAn2IIyC3InboPR0lMwF6CCC3WWh86ippMMqJ4+INTqB1PbuPL8Wx2KRzHh+u+Eda
iCfn5Oy4CfcrBjNJkl5okJBcnsvwT8S3eknrexMQorBYkoR5n6q1OL9Q/8UU9Eqpn4H1ycUeLsEk
tClYbsloVV1YkerBbtBDhds7X/yl3DvAbCdCwaSKNX1MQWx3n6f0f6ZXnPUyqOUsIduyoz5DEUod
JgytpttIY0kYgmTcld9TQjHdeq6xT+79hSro0gG9XOP9pPBUXN9gkOLyt8ePx9POJac5M6VP2PaJ
1H1LqBzvYfQO6Qu6sHwEW4TEPhk26FKmCF5e3sbVpoL2HQiZSLmGBHBMqwS4iYGJuo+B8+s8vlk6
y/GA6GdaYE0/JI6qvpjBbTuFWTyKdIpxgUKXYfmBDq0zMhL46Ak7Xye9eVy8ch8sXYNTzXuO18sS
jAFfNM7y8M3EAUb9/I51JYt3nx0mGtB2Oq1xt2fd0CQjgiNw/lyTb2s+x5Gnb1iuA5C/KZ2h9+SQ
cR/BCv3KQNNlHr7rYJtFf17EFyCd3oJ6EFms6CmNWZuetN60Bav5LgURyvvN5F4lLh84eFkKn548
UVD+nE31iQmB/PuM5JT5S2GblBouaeBNMn/+//LJSbKKNvjduTMXyNZCBj10kqdBSW2KtwQ+SzYQ
Zz83QUnlyeDArxYUinuXpoounBhez3qk0hz//GMf+ielpLFaeE8tMrTKV6cOF4uBh30QAk6+lD87
8tAGFcBQNM4hlz0MZNHrRmoPt/YYmZBoZpM0sBP0DY6N4zFB7KB+TO7XeNpGo91Fhni58jRRtxpI
h9KihQMBZ81mtOvJmq2tKbbVu08c906LNVyLwM2OD6si+q+tKh6EUOlfneeuKAiSazws/nZNMkXs
rKDhb1oK+miQblbMbeIfSrif7BeCVbK4Vu25BZtoozxNUcQKDIYnt/Z2nTGci+l7vhkM91btOBbD
DsnDdGjaSehEGMIt/LURPjMEyHiVWteePANPgF0Iyjl3f+4FGuj/3BtZvFqQj5PwTckv1TyUBDaI
NYNpY9eVvVl6dTQopCqRaJCh8T0KYkaT5jtEili4jCGeVnu2Pf7rsl4qawuEVc4kk7/GVxxehHSo
xqkCnL6VaCOHvS0R9iWXF3qGXHY4A7GSr/ZKgHkH0KXIh2SROj2nfhyJQlaSCtxI9NRnNyHdMhIX
12PeSRhnXhZrggcnDQilvZJRIJ6lUHgHCla0GvPRj2bp5rLXRE6ULg6XKzquAjTafKtJ13TDnbeV
3zm8h8yum3olsUOuxXwtJz4BpMGLyodHb8EGEjyx6/XIgoeIm+5xSxAKlP9vwUb4spDvg8DxFFRH
VLzVASK3ecbIiy2zdzhKvhNuSdrJ1hUOCDmpXKIglMC5ziFmb/1FQiF3JJy9rr3uaBL6ygzs2lHq
TpGfcd+4pYeceLjWMf9Qz3/cVmEOngoSctMqhri4/YO44VaT9jAj7UNPjzYYOjQ8f/fK+5Uo7qxf
y5QpFXgJdxsSLJVoxWfYbZMvoezg5KWoCuCQs1BIX3HKi3Z7aVYdvzadVaE3jg/ZSeAysrNDGUwf
IOhbpQzRNAQCl591W9mZcsxroSYx/7Lm8UPlE7G39pwkh62nH9p5zOVSysdtN8sueKxtHzrw4tpW
7we1FOKqlXu5/Is+IGkSwdODgEkEkzJeGLcDCvL1f8flaFvw8XqPmtydCnPS26v/yDhyflKnDXul
j01tO0mgRWVdq4lCY1kYVRe0cSNhZeQTn8MwrlcTlS4imXD1AAQ089sUM29vzMq4lzhTZbd9mU9G
FSBWlLkLVPEqN6+vW9oaOyOZGUAr1Cz6yJq72fohhW1iinSh9wRnsGco0a3q1jzxwpm+4eGGL74v
amW4AkQ2GdPvylV11RbBvM6GUqdsng6DsrT7T84o8SImSDct4xEa6z5oOx0gnYHY/5PvYrbQ2hd4
U+mGFFXVCuy+xS/7IdzdUGkb9l3bQ3oLzI7rIKXh3beW8vwZQr6us1SUaCAKICOwimhX6S086B+N
J23Qky5bAgRBJgIQv3/iguGbfDMYCPzwXbdilCla5FlMdXhWQQYkHvoC62eJT+Q6Lp16K/nVK0Hm
tLfxoV+TtfHnKEDypzfvlodnd8SXRvlL9+lnfYki/RGshqfreUzgNzEoWfhw5biNdMIw2Qa6EW8r
d0Cxt2CNFcjth9nvMu2Ww2qSqIUPHTUIbpaRny7qXalR4z74VntrXGxyEX7F31e6HaSl64JOVvPf
oKwt0WrO/EKV5ZpL4CaIulYioqdKF+kYfNpqExHBlXY0ard03hq0D9lwJCtNKa1cEf+flJRakqTF
GyKGg0CVGe+VCUwLgxVRaLdP8twCjNpPMXYwtyT7RK2lOde3AcDITzmoVBcKT9+E0S/JTtOWWlAM
a+VYgIJIXbaKqYQKAaUFMeIhm1x7cs6ckviYVqSSTRP2/5cQAJJ2zeuSHXLVxLqxDUyiE25cICs+
Ykp9eexHg5vXZSFuI6ICJihROpAaaFYfpwucwttwVp3d9K1YAr+be71xpqdF1pIpw2ZSUiVJNdpB
pOKxPCp/nn0/qaFXFotu/KA0DQMz/XRHKTUh3+G0Ak/YTTMLFY8uHYj3QAfa7gBDZSEVuTpSTeQN
ovkF3dbz81U6ICyChvaQZfqlqi7JYKvLsOsTTv7gnEKuRUqc0N6WaDuR6AjUUsmZQLUlPtUsNaDc
7tyj1UVw03yzZBbBa188NF4CrVfQPgXoPtcrrr69qrmGBLvKPq+V4bXSKBPdJlx+rKWK+zFn4iOk
W4Ow+yZ+aagZ8yqntp5+mfpEDbGbv/Kj3BmiiiLzfSJFs/6hJxyVX6TChQGAPnUc5Z6drOpzV0yX
vyPV05pF4PIRR1tnvF+bpjWnERGBEx7+SBHYAVU73RXxvEgF2Djl+tMH04qqbHuP3DyeATJHWEc4
QQd+Vc5Ike5t+g8UPYNx0lnSM5w5tlq0aGhglXELBZbdvG1vJfhI5V9uFA9nuD7Jn2rrOMn7EOhS
4Q8VAVD/g23d+WfttvEmpXHixYZv472c9Z4NgKcH2Flq4/z+FClDyK1Qm31gqLmRL1ciDxvTUqtU
uPKGiS4046qkfEJvK8pZe0YmgwyNQ6Zx41NiQWcaa58D9eImSKfnip2nYhs1oiTXid2lVsBRNHcz
zsAt9Iu0n3DqfpShB2adJl42ikfOBq0sS0sGLTeEQe8cF2yrXz1sQSEg5zQjQfbv9e8QfGpNvrMO
t6BN1H7zNT5xhsZqclUg7coz4B03YhrB1VwYMa4DE4Ch+ZsC9mzX4QmOuL2bi4TDtl/EChh7P9Kq
XebBTUIvjLqHnSdIjt0rC9bsOYA1F1/QtLrSybCpeFAGCeMWqFRr99Rq9FWUFxfLmy/icK4vetpu
+gyb3y6QZ1O1hU2kTqnAKvV/bK3q5jBj/AJj8rq8tv+7rC1+3JD0ODL1btbjW9pfX3oWbxBeWK6S
9wccoLSnk3JYx4znJOdpONQ3FLNowWUBrxK0DIALCTH/VIxjWhxY8N11ZqCNp9Gj659VNe7uhdcf
V61if6+xAdVCUTyZvLAd5UI5p5q21duXEJxQb0rzuPh+4D+TPVRm5N2XJtZsh3gFB0KxI3PvbXOz
3s8F7E8MtiLDAJEWO/wvnjBrxWq2yQor7+rx2ANwuouBW2sVn6iHtTxW0gavyNBqZQk5MonAi7w5
DjmOdZswza5PbmzuUBRPYeeOXWH6BUazVI0/GcP7qhrs9G4JOK0KEJLDOBk/t40svmtH63BPOTdk
hDlODVS3aV7XYsLJ9vxVKk/x4MkQ+s4dLRbAWZIzNf4iCqe0cmPmxMR/q25hgR8m0W+gJRgd9gel
y3AFfSU+42pIqC/fW9Kbgq0JPdBVqcF2TsTvac9U3tMStZ65H3OYtJM1sC3h48lOPpkY2MrdZAb+
uebQfaiTCjP+qDvCXKTZWVBlFzazkJOI00eCgWFTkPbAnVxF/NXbph0J/JMERkKnTOILF3A1yMyE
fU0V5n6hQFjNvyAL84BXY1Xp+CsHxOkoQdHSoavsLu4xDJLM2gxQQdS/u2o5qlbPzzg2cxum/165
+1CQSzrEmVMVM2nl+hW5EI/sUgzR1Ylmi6SWRz8TtcYtETzKyKIOHBEEBALaf34FKLZ3/Y0ooX+e
3NMDYWGIZe6n8BPtM7P4FCrucxIPo1raFz2bwYfvGxs7kK/y1ie288qa3zyxzAnYQs2BPM1rfVGs
C9SW4Z19e7pV9Qp8UB/U6tNavlqXi7JLcMdWs81KFNFKUbyRi8Ma0J/txDTy1keyFGloCbQFJ9uA
J9DqeOTfiXXlPMJWrcux/A/MzEH5bspAwkcWkJC4iRJYssULWCvYOrz1DYS18tlkbJBNkjKaqXST
9sfxJQO1K5uEdrh36a2BfYRTLP9tEtjf3S2aiOO+rATYFifLW3UyVHMW3QCtQhtGZz7mvN+M/K9G
YR0ntGQfhqv+PKg6yRB8UmNvghfwXW77M0tkvrgSSdc9dzB7H/gF5M+bg/tkgMZvsj55XvXfIQJN
TlNBeOb2oMF1eX5hUAv/UFFh4HcKFgRk4SDliT0ZVvjX1+rwaAfJPsnnLn8EnHfzLgUmNcrsAr2A
xgGrRQYloT+/dvqUg1bdKxFffEIhn7x27M2/8crAlBj3oqqGEY+oJ1Xl/iWlkQ2vocraTev/Gsjs
DpARlAvSR2bKikpE7p3Fe1jW+8NUglhJRxBYRmD09sTSGMAIm+3LJyh3Wt6ATEYBIjGNAcfTKa/M
oyNe03piCQVIX7ZBJ8oRI2joQAlKZ5RFLEe2dhcoxj0XMxLdDRXz64A8HI55wbzkE5MxyCLDdY2C
0jC/cyu04Bcm7OTEPiJSs5nyqlyB0bMrdHZGrt2deqourjfPyWQ+BqfgOfGiraF9hIBcHby7RP/f
Be6enhLnyfCrwTxQYc4UT5ZWtM8yL8SI7S0EuWmNSCu2VISHctS9lI0o2yrPUlC7wyE4sJyAN9ua
bPf02hkos0iuhrPlOuOLLBZn05bW2W6MX2rO2VNok8pLoLQSZSF/YaCdL3MKzuON6dasbaDphp6D
rLLOpcWNTQcv0Pzd3Hk9ADkgrepxlUEA5UmlbMPi5LfCBiKQiSAsRmE4Ao9ELWQtJ2gO7fGjx9XW
uVS5jdgP8bPRmTZ4fLLEb4Ugqm1tWehmyuZ63f/7YS2fr1MLC5G9u13ulyshSO7ORBZxm8tmiOrN
jEWvJGm7uVTqI9439zVp8Iywgc0fWOsvKvWyOYLOR5pWRl8hBUNjb7xNDiOMDcwOEpkSG3PZaATN
lCgWbMb8tfZ0GzN5qwNQNxzRcv67iq/raMwFQgW0K/NET0bGctQ6hcHsnrEIe02BKva0BH4EUt4y
3rFxthblXVAq10wKLOdZPTRUl9cr3IqWQq9TLLgu+BoS9t0RhxTaBsdN+KhHsZUZnxvl/2sUsiFx
qknlbf3tgb5f6yiVttwR9NJFBuxh5sqUrXn5STJPZIFilX7ElJ8ca5+7RxFgHaEgjYyu/M5ccYaa
1AjDUTI9qVB28DrFV+M6Y5WaS8YfwxiB2qMcVLxRX5e50BGUUEcEvyFtXQX7CEw9hDtFzCgaRapL
RpR2AQyca0t4nNO9Jjy2C7xgUZk4dVG0X7+U7G6urhQ68/6R6jAMe1ejovu+6+KG+rXnXv8A/2rw
mSzclox6ec/zwBVHNT+xtkTrIsfz/TYa/vmIR+osG1BnQD9NJ6lwMsAX/x6UMbYcxiaqPY7Ows4M
kDVBaFyENKGtwLBMXGHB+SoF7PgfwYReYNc4xemOgTr0iB7ddYZTZ5N9SYbGTYcfsz2YdDGV8Hnj
hduOEsUiM2yabfab26n4NhQbpzzkS87VH2yXkgr7VlNTUSnlGleFUgFWQIUH2UfPcVv5GoP2da0C
cWJDh2UYSnbPjlQorPm33+7DcvhnCGrySRdtCeaL9dK/M9KgArSBpk4a7VqCehQ8zxTxeTyqQvyZ
I2ciwTjcO6bazxcLsJPNtBEEX7I5tK2qnzocSOcZ7fXKc9opE2lNY+e1Vb7taFolNBhC95tg3Wbc
WtMUK3i9gar/J/7Y1t4368FvEQu9jrBT4p/b/JBzE5w6AsNiPhvP3k7u4QGUYrW2/ocIrKN5Ka9t
TouXFpYp9lRQ9nL0x6ZC0Nke+0gcvM+ncYmf5wPKWQz01chtp008Dwi2qNUhdmOsDz1rWuO209Ls
oPZ3EbGX/Oxm00JaXFH0vlvnn0bnuQp/43EShnQpED30Rp5sYlLAZt2XjXjyVqBuP2TsGKHe1agf
MTgNcX7S+Et+LEbb0s5ycSNzX6w84J2hG8sBOwKktmHSfLW+Zyf/Z0T0XQIQfxKnx978D4wdzCvb
JeQBOGD4TDMfnjGOKBcmGHRso2byMoNze0LLx7DxUWVnO74yDb9GAkuLlq8a+bnPDm+XKi6y7v0c
cKEK9Cz8iIJ4GI7jOmvCuLvE+xXhPTz18/YSxqmulxTIEvaZmJPNg/cLtFzA3rUKmiCPW14ClYXl
oYnVHZJiWv4pqhdStDuj4VaSRGo4ZgRLfRhZJmHZiffGnJZR+dqVu/5tp+sXcCSDHTDIl6levYiN
+wov5M5mP9CiJ0BrMXROJ3ews0MnS8eWCsocXLvRNAuKCdKhXPpeaiNYNExDYkLek95xFkHcsK4F
SPV8ZN24UcpJ51JRRn133yIOeceC45pBjoVm2K+8H3oDdC2jwDaftToFF7arlgYxOac6v48+SMpr
tjEsVimPlz1beXqU4/xcrj3giH3P8ebRA6ZnIJmq15YKN9DlKluwUg6SRddWEr4GwkGvw3uyr/PD
hnBYHgFts1cbAS+lDCcvbHOO0n7q5NRNdLRqP3JaJEyIARkbVGBD2C3DfVrZChToziyX61MqgQfl
cRUhkYBRxgoTrdxp06bv0nPSplb3T/+En+b7ZZHxK4s8fs1XH0NW2YrxGppq45LRB7u/8VbHo34M
3etYrhPdXBcTQpgf+wnQYFmVQjc0GYDSdKPwOa7pt5x0Zq1GUqU9TbC4iDWcAgfNjgeAef6PuQQS
P6mZ1qCePaDmX1BY4QcBCq0EiUyIQ2Gev5iA20X8OsX+MOqZEEC3wpA5IrVWmbzc78V/Ob26Md+C
6yVr+2WBreXaS7tYwaU3CJp1EbOPPWfgZqmpmlKp539gAAxltenOFnJN7jUdbkhDQjT2LWvMBMN6
YfzTmn2YS/pEqZQFiw6hMCgjFXZQRiZsU0mF5GsxWRiIDFjdFX+zj+9ypzsIT1U+2wBrvjTZ60L1
1YHQPhjfmU/QoS3TLF966GlH4Qmn1FEvCmp4mizdCXONvAYo3WhIuwf7zePHx6TlitlcEahPzn6J
wGCh/nVN3q24ilweGyBqA9QMXO2ZyFyHzT/Pe6AsfAixQ9lWNPFanGgEeF+ijGBJbqkDdAXTIz4R
0/sINv2FmHIFopJ7tqkIUVRS8a+cub0ZxSgvCaBxd5QAhtA3OL+g6yq1ve0PbhxuTGfaT9vlQbdF
3kPOwzGIeq/vU6JBC20VdawZnb0TXTFXaPN2PJrOIaBHlvT/eqQuV4ohdtNySAf44P6is4C3ldH7
xTMDa3kW0j4SsO09KroTwn1YsVccxeqLSj4lRoLkGbpKHDaOavnPY9keuV/M3ON571E7b8t5hCRA
NI/ip81313KNth6Jgdq2yhs8Ig4tzui9dkdqrihLovrnq4Qytc/TsUB50hBPLYKMWVpqKiRWKz2g
Rt4tCn4IMERmBCxzUfjrtJoVStxCP7KrJXwr/3nhZ5KOKP4+7n31dvF8blg28JHG9m8QN94NTBr1
4D6Mm9KoBwQ/Gkco5D1kU+AJ3DzKEow+DPrxibvCoSGxjb5kHiPmzrc858ioX11V448pVd2wazbM
oeBvLnBAm+UpzWENvGWX2+7lyZfesj+x0Z+00U6TS23w8xAa+M/NDleU17sbeNeQW/KDqV5kXSHN
87mnmYMOpyHVf/De76SOf6KQvduA4dlq7FC+r6zTdkvMtijkWcqnzjWp6fdyPDzyiXL1z2L1ymBB
55bdlsG/LPK5SgpngIrqDP7sfKCMJtxQqkdH7F3Y0YJ5ZBa42NciS3SLV7lplbGvcSD7TV+rjJ/0
5Z5ztGLcRs8vZ64WHvGhw61n1vF9eQHjmkNfI3IYzWOeBkBj40eKDrmOd/vb+ZPYYy0WBGFKqsdB
nKGwJqWxIxkcfInVUM6ROf+yKtbDJ38T6E4OXKCrTj3nih0AgtvPiHU1sI7ii3YXfpHmKqc8658+
wGDj4+oMWhkyW58ipyCeFR7f8k/+aoINB/CL24XELgY5j6dN9rhuYzQL73uKmmPPiFEP/LhAS6GG
ZkXetav9aS6q7BtLo6cGN6QqvHLzH83yd6mSi4gqSeQoc+tCKMpx9svzmb7G3Yc0IyYfEUf76yVM
V7h9IkmCsqnlNrONVQ07vZd/kifFVUnAnim5PlgoU6NxxqcLxaqFKeCnp1+S6nONTYBlBr+Y/R0h
qMb/dS5WVQBzMJYKhUYmLoVYV+gAB3fW8ZOaEYt9cxGjFhCqR41gmWy5niKyiNJkvUFwpagXkyfp
0G9bppXIZJZdsf1GQoO2OQGsJ4gdUgj/zeZuIXYzTbwV3NbCahY70bMrWeZB5FZj0/IvmBVrJkO+
G5uSi44yo6i/d0NbHw3CJxKbstVb4kHDWyWJ+KmAli0l9O2W4REtvdCWtlX3oR91/sTyetab4jxv
PhE65yA9zFS2AKLt1I1lRiI17lLr0tzWrpxSB0VNr32JgFkNny/LeXeDPMUFDna7TUXprxQDtDNg
quvKwOeVh+t0hHi+iPWfqS6VPgfcy1CirjtZxSOWAx0wsR47x8tJvSZMEoSEhftEB8q1V8ax3nRY
7WqrI9I8VeZCF/T1xlE5MNeg2Q3KEVkzAnLiGq6p/ivX5G8/OzoyDKq9w8+Ty1Bd6JVtFTNmA6w8
VS3wPZFMHt9hFHAJ8d7BWyk4Vt91lObr0vGPtu1mKbjPKkxJSvp96fs9AmxuBRWlK4q4ot9rKkmT
Vm2nLXgrC5YTcdgsVUomk6T2PelC3pbHUZXz5hk4NUpRUjUa2qZ5S+bh9BBF+jZ4HE1DDhycXqQX
Z6elDtsFevUsgZrC90fH+/zzs5Wzuf/6EFNeosElaqq4ZHm4MuOAqt7dNuAwv/x0c1jI9I/4C1s2
dLS8piGG6juMchLxXisoGM1QLBe4d2nH8yHpa3ucBBehMlyeMFoMogJuQrv9l75KuzrLZ5M/v+Ql
6rvSqHmuuUOGB/mPCxUgoyxdxvIqtfkhma1V8woURM7LTiR1Y+skAf2zvt5Ftb4HbIE33roFU/it
wsvz5qxWuIPyDTUG9mPv/n+uLguab+6wUvnwiygdhB7DECu2VYKpKsDlx0YUMNUvSRT+PfXGGn0K
SyUS6Wrh6zfHpIdsB9hiJzmlOk24uIFdNuMQS/b4q2QkVWxyNaAWbYdOP2FNogJM2iK7xsewVAzi
Qf1xj2Kw5B2kneN1tfDZkJGWHtmi2qiJNrwzc4Jv0330kQgLx8YFTzX8wDMIZFE5PB1b7+AS1BcS
GJAqR1n9OPMkPmF/GrfX6LzqsUTUqmfeQS3WgGdsdVHlhYT2HhffTCDQN3yHRw9S+pJCm1wJCtQp
jpYVMtr7pTltGdQ3ng2r+6SLnjMG0PFboHNgvDVb7dHBSFrQpWxa8f/elviUMOtA9XcwR2p1rok0
VV+pseIBiO+dVKI62QPSCxHWCv2oOYlUjFrmfQFFr5/znCVJjx9jOcHVBM32W1X+UM3RIQohPsih
yvl8XyeEqwQN/kJ7/+5iK591OxYA8WJpK0GGaPq4954jtAqdQ8P4dRb0302+K6fa4fYRciAXTkYR
3F0zGjgTO2IdEFsQzx0z6oWpcv3Gz9ydimZP7dDtmFSdiC80q8drdk3jv10pymvavKWsFex4U2YX
+nY0wWjNblyMOgnN0mR3Q0Ara9EQJo94eO/O7BDwVof9IYTKTNtk16TGVq8CeyB5kqAW6802tl4r
Sg1UG643iIwdmmohtWWNElAs1NbyDMf/MdZOmUcO5YCLNDgVZj5xxNsyfkmYH0LyPm2AA4Om7+ma
6np2VQHgxIvq1UVJ31bW6jK+EiWZe4wfsyi0YweZsDEl2b6CKUUlRsNtGfsTYzcz+pL7iavGn1Vx
Wtyag0yHiM6PWEj41jt/PQYPdCg+U9+rkNkSahieyOqWHFyHikVe1LMDDRNRTQTUJmE0bhsKn98z
BWOOHoTowazrbqe81TlqUW8k4kniR7qUlfASbxbPBTiuak9tmuzq+JTtvuOTBeDL+xbrKf9ut64A
wQLmYsw4k3ccFESuyY2C4zVe/DPI59xh49Nk4621Omi1CNX1bqrjWybwu2kLh0xwINeZbeUTqlr3
6lL+R/xNtZi0sY+wbkMxF/ADA6toWZePwTMgCPXMpnQvDYWOIXpnPu09xvoJJy6WRyTdCgwVffu7
iETZehqlBMCLI9DUxjUR9du4Djy9XZUijCeTT3EOtXvQ3sWjdPv2t6RHy1N6ia99RcPEdSrblHQL
ZHFDtYSCi7SgKm3BBeXiSCOuaVNGxBgmLsNLoxMvSH+qouwVC+NwuALe1gA0Bl2dTQ7NUW4xWL7f
hWIuiV1vDYS49L5EXnMmNLgO/OGAydvJnNZITNpR0c/aVuUE/pAKdegFyws+u7n41TvIDvm64HVh
mcSNgHxXMMMIF4WQPQlNth+wiQcT2AeH/6fVHiUzUuncauaJn4jhyZZzfo7NB3zz37uDP8KiWL3W
LhhAEY+Ym85OMK9uYB7XLLWDcZK7hWW7SAqB1iGCndZ3WUXNg+Mw99Y7pInoAxulm4ljO7Sn7LTA
UbrZ9SeOW43XsQ1fFrQ11Tc7gA1/uf/RWcIEAcyDPVNG9MgpMK59pN63fx+nmaXply5WbxQNbzZz
JgduUqo5DuzxAaVWeDyngBf3ROp58+350iXNdP2CgbhW/nhxFfnrItF10BFe4W9wTktrjFPahp4Q
JoA0MVz2eFEn1YY4wREYPNjeZYrWUjHsz5DyV2Lk2UHT1RNkGTRM4uscuBObWNsq1gIIuSx62/S2
BWN2itYaQl4ZntVXePrVIEZzxO/dOTE/w/78hsp62nYACurMfpoJu6+AHzicPdiRrCrCE22+3a/x
0I1cTzx+5llDZ+K0WnFBBjcsaxlRPCPZJN1nZ9YH2Jex6nZTKgM2lxpcMDSKq29Zc/qwhArIOUpW
hVqnVnpS8o89FLppEoEr9sIBwl7x8ptemPyjHGtIXxAzMPW87ctxLikfbA+vF+J6PFJoliIMkPb6
0o7snOMeMmiJHBOYqqYnFZVBTz+sjqQOcZ7ymZ9nncS0t6hpfrayKFM7WvCcVaazEddwJ1lAHR5j
8FGeDhEUOSWO1U/4HWANWCykp1gknIk68V6pfmSimmqnjzP55mKvcOn+FOJjevEgtuR6KQ0cW2gQ
kywYRo43m06CI30OmwAUfHGEu9+5wYT52LJFm6KVC2woZvMPeaWQNPkY6nj1JmP+aHcHr0DQo3zb
zroASqwsqrz5HH6QrTgh78m7c9wJuBk4bvQMGTov4A5y3ktt5Uw3HKEUb0GfoY8deQWmSwkOBVbk
QBv9O+iI/sILyIMAw96B/6yQWau2MgrK1c4nuqsqyEWVudoh8kmhNdFL61ySCLbFz8uhon0Z3qjF
YuUICVspYOXaRvjLNwS84caZMFLKlDVuVIm8ncUWQAoV/kHhI1rq87XNfjX/wYi5w2cmh8grAMIp
q1ze0/aNwH1RJeMr6j8XUDFG4BsFz6bFPRVLfMJ8i0W4CSC6rJnwyRV11xsfN3dfHzVCfgzZKgET
7f5mvGKEjzg7WaUK1LdPPAjPMQtkHEsdWR7YT781OrNa1Nr2gDbzscEwHk6PCygmRgmp7ZSplhnk
HuQBz1TqL0Gae4EQZXduJHIzl5Geg9CSxMa4TQrkfin4jENKklTSG3MIYid68PUxk7IrzrvYuZEB
lGUZHoNtVWx4wtFNVy9rvUkCt0SeURMMISa9ohTMlAgHxnT+mgMIt0M/1W2hIt10eAwdden16MbB
VtSs2Zv3Zqqo+aVVG7PQ9EujktTXToJ0omYkdG05tLNVfPaKyx1X7yfGblX5dM2usdOK+rQ7S2vP
YA11GZjozcZtXhVFVosA4rBs9IU6GSe/6BXY544WPUgWx9JMtToOh9nBmjkGS4+1uSnQtFUalseF
kIPOY+yMWdixT2aDNNSf/95q5LKTt2dEFfb4mEzaXeMNOtqPJEQ8fEeJ/4EGKgvuGGXElaoXhGsY
NqPP4HJ4fwSJoOa+TC2cIogUW3gBFuxtIl5rBEEdEpqdr7ELBYUs4Tje0cW32l5/XjalXNzUfANB
NCyD8yEYJIzT5mx0r/z5Pw8iUyqBKKwctQn8iKWBYGC0BO1V+dQm+04cksx5rAwRO7Jkq5PfjB9F
v5hOnWlg/PtGhSBGXBbdl6yJye/EyFZu0nT3+RLrXCdH0doo5GGL40MQZEKQ5jMPQge+NbfCkHXb
A0gyJBu45K3iMeDMgJIi86FKHim9vy0fkWVqvrKm4N4beuets+tOYvzO0HRKbYJ/GO+libumw+Rm
DnMhd+r4TRw4LfNdLIqKQF+J3UaHXcGm0NMqZ6mxSs/liggrc+gkjF6S+ZcjbgcYmcj8w78Ka3Tl
WAZW+reZzw95NuhWPH09MapwjBIlUtkdxHVqgE2ciNRgqlun7MLZori6sceulKllRAiPmJyAhEZZ
EnHPdoEU4D8H9QpS4eElQXj2nR0iI1cfLPj/508va6OxWbT62T38aTpxnh6Ux5gLf0PoUOz5bTpe
Tqs6TPdmWtOXkqUaZySJ17swrXrJN5wkT8sAXLbwnoT9jwTLnNV1wUwC55XmsQSaUTYhRdjpqlrj
j7nYe8ce1imvyvzf3/QXhwvMU2OIpiC93yAs5QHjjCjAAb9bmBxMdLCiEmzQOrVUu+6jDfHVXJ6Z
fn+tSyb8FjkH3eYEDy0aFaX4z1ibZ6BsK8WyGFzFlx9UvLqAa0iFf0UGbFAkbRbfQ+/5ioVz6g6V
ufQyKpTl/hNZJ97t2F+csQ/lKO1stBRv6cFwVE2WW7tZbqf9y0CmM9btv4/qrwMWJE+zKv5d2VUt
0uOau5khvqsZTEEt5UZcsYPECaCW39a9D+Km6joNkBksoyC7u+TD9kEWi8p3PrFtAhheBC+OjzVj
E4bI1VZLj+6vKAM8LhJCx5nLQszDmcsi/yq98VLGHNwDN5yxWgFWqGlDOi3Uu5r/0GO2PaI0IJBW
9+yKq8Ya0kk53xhh42ZeR/zPmS+ePLWCilRNnxLtuFuKI461c8ctQWV8ijNzZ91bmyzB4Et2GaRQ
95uLbUcVFlS2nK1LbwtqneH0Ofr6Bvaaq7+AuEkuhwGUs55asJKenIpkGD6GHJ/F1gncquTIQzrb
WzQTEIfDKbDPy49bbvfLYL605HD9TTt/2/NwjoeAy7KavaBxirDOl4R2zKj7fDf3Qws3c6/dVog9
DCVjAsXFm33MHaDneoOA14ENI28MeGYdhaKoNwR0epjiGi8OMNuqon51KihiZwUpvEGBS/VLoIQI
HLvbCYJNCzOEFoWNNaDxmfKPBZs1qEtaLL7v8yVm1stmwFm/E9LuR/QEtnBPlcrePTKIN0q+g1b2
o/ciwvhGAtMEAPPtKcqNtnxEqk6QLErnJXPQ9nD7eokYPmajP8G42oxhW1CxT5vMYUM4rtOmFpTY
/HMPBB0s/s8Y80RrAbIHLh8Oh6T/fVrkbb9HF9NKkKCTrzDTtKOEnyYlB/iRLNt3RwHwWVtA0b1E
X8UuY9HSArQT775KJintusd2XAXx0SVka6NWVzfaNvhCPbMw65i9JJhZQ12dkNgudi7068Jzlurm
atl5Vb4LRWKd5T8npxNbAUlCrhP7yx5d+yve/zXDIEeS4Y5OC+rLaMKxl/J/b7Zh7t8Hn0rBSfUs
8B9GWGWs6WSBl3FKDujuWpP+Pu5XvpF85Mwuo8WHr4eaeLHI6jQQcnZuko0VNZoTkxFe1+gt3tP0
N+QQiCgzCWUo24QCONekMUCgTo/CUkG2SxsoQOW+8enpcC70t2sAznlqoao6OQrK0asH0/vODtHv
IJfIe1trVdtJD+WyNKuABsu91d1C8sgan2urZiBbbwut+qwPeGktVrmT/dLXd1hhqLgrMoJyT+50
K/zuy4mFK628MaUe1A67CUbkkVhMOGSgaiqgfKjkrkZBCxRbSgDul3GOVyTETQGvmidhCpTd7tTw
uGKE7rlwzoORrA40d9yIlF/y16k+jZ8zPbhZnzvKF++w0WwFWMnGwZjZLIv0mx0LXXKfn2Y9s/Ni
4sPJvrSjXxfd5tbCBUdhuClB64MO4S80UX2KViIWYEB7PL8ImStDnZd1XGpWHMBsVCXxFvAyWnx3
A60/XGu66cKla8HzZB+Q+QOX4xPAKRewVZQnUeCF7ZZplTHKEV7EeLFMmllUNgpPcJFgO9ai+0aN
mK0EeWqogy65TFKZbfUSK3JipYNrwaZVSKn3p7hlZpr3B2FjGveMeuuf0zE4u1t+ThFUJQFiKlHH
UVLV4jZBe1OFCnC8VKs8p4ZLlrXsekQvgnEQ+lLbWkU+xROSZgKwrucMasNrkmukY0RTgGnLDHLM
CicNcpvENA+gehUl0a1lJ6TEa2o0KfoKrijj8UCL1o/qQ55nqGkJfmQZEnyh2wAQprfzZeaGXfX5
w77G3Kpl5ckdrFOqXEr3/Xh85AJdmjxKfKePbJ1m2TlOsa22SP6oHB2Z7lwNLYW3G5wuwwyMrGQn
p3FZUa3W/zRp/a1+UYNAg2eFFahjcWoO6Zi7W3s1z5vFoaxtc6XFEjIqOAAa4750eMT4F0+eRFCQ
+2kLUU15p6O1CgzV2D1XKxyd26L70Y5P4eEA1HguzQlR23gyyeHM2jqtOzp3UToR5SvSZe7rH8rT
+l79CuHpIRI5fxoAKQIYPoExwfvaUBp3PWofhXj/zj3s68RmrAnZ/VnFPePXRopkfjkyfr8+7KfY
C3jYSCsdQOkC159DsctrZIrthOOxKtt1BQCE/GrhhPcG03MHjtHPmFqPEIQP+lVbj1qZnmLISTvu
Q6u1nHDSKgceacH3rUKPznkd76CnPlKqVVxMKScpO2UofpFWser53dme0nKHKMwNEONkL7rEDMBI
GLXYKzjUsVWrBRjdPC9NDjwAy5k9/ghC0FyvXqP8pow1ht6Ph3FgymUKQpxcxH+6xdDPx/EkTk94
75AWKAOZbX1/0RShMDy2DsA9WhF88qJLyg9G8V6mwf185dPEm/asQfP4guG5y1aHHjX9GlY+0zH2
unWvw/3DioFVBuUpcQvfoGw1OCkqJzcE1v7Ou4vErbyM7PZCNb1LlHcpvb0YQND/orY5/zwbU8J/
dpT/U7uJwfIXIoLCkzB2E4FeiKtmG2gMhljdwhwj6FmJ5A2LAxlgM78DAihVF3TpqPPm93JvWiNF
fFVHe1m3Nok5+1qdxGBfaJFPz3W61JZEzH0J2A5vwPDwe93xoQFmxmOl2kqekMKGZHqZDgXix6oH
tIGj5bO9yJWGa9JBQhY+oo6Rz1ugkY1OYFqmiMlGGMuH74vQlE+uvP0zjM30pMiS8/bkpof4c75Y
VIvJBTGfMz5PMK/4IXu7NIhXwFDuOwOJAW1HxKezeJFOpwtTJxNj8qOqs63eC+YIfZeKw6ZQLdpF
JvqOtI045M/x+sDcayeGKcnXCtt9lkszZP+zMrqmmnWRFGU8bz0mBoVHMLmlY7IxjO6LNVzJXWsA
0Bijr1Rboor3T2xewMJgzgt+UxNqBuze0D2I67+UnzgMrHXiHyq/ducPpXQ/CQv3LcPB+ZmzfFd4
F+CklNEUBVXm4s08jm3T6ZwPdOC/61VZVrZVWjJDj4/KCojboZJROUj6B9TnPFbgHm3Dw0crDaY5
QeYYh9jtKFKiiIPCVmAHRkhQRxWAIodhyV9UBSG7B5EqUWDgG0ihYtPNt4TJp2LyKPTqmCrV0q+V
xYZn9OCpER85VktDthhGg3B0otfUTy1VAvjWdgratfIbm3QQr2K8nYHyITM26kB/rw8VUFNU1a/U
wl4nHUKBCz+dfwjgByZSrWrHHMJ2wvmZr1omVdGm8hN/fvv7Tzr08tbA7M91e57Z88FZ2TTwPLSh
G0QHMm6i5dDuVJ/YkksmjQIiRJbGvy6PxODlFKiWufPDg5WEKdajbtGENV6KVR4m4AlhHGVE1lEO
zIiCutUwTKRhEeJZQO4SuordUKUPJCBVmh24SDs8bCAEauJIprKZI2GQEfxWIqLMxfVl+yC8PpLr
4gpMKH2+cE3N0HAmLKpiyGCytviTs/tO/KZY4oSeh1AJwPyTU1Fb8cd2JDsKtbIdhOdGlyBMJuOZ
IVCpcfmxCD8v/e/vqQVQaOyTdUk84WwqzLbf7ep5a6snOEieG7BYa1nvcVXD6rNm7TAH+qW6T0hU
D5AkV5dsU4K6OhNcrOZirD7nrtbiU0Cy+Sibc7qqwTRTa3by7Sg71DkqaNbDlKvhNmxSXsDfDqnp
4fb+auhb3BXxGFgsiEdv7XDZpT9aqThfUYn/pd9eHxI7o4T3365tCHKStocqCty0qYfSlGY2iDfk
AYhPDTDOyR5iVCixLr6D04Ew1OMvPlJrOJHxDrECD3B4c/nh2t7C8PPKwcgkSnjOt+rtRNT4W354
0XQPfhgReh3NnfCQDmfL1wDdurdH28tFV0EdrUh0oTkPCssiT9PIXiPf/SCBFD65yl6PQzBtHG+0
cnVTJefpn2oT4ea5XDe85eKTY8YFMmL01oOFSEmZcCNIRxJ9fF6zkB0hLUbUAq+Kux62TPlcUnqs
Qt090cDT/iKduasu3SE6FqivatTPpSnULPbOHoOg7847xnTyvlV2UPBdbfUWB8o2VsUvcNWuK/LX
u+e8W6J+D0m1rDHKM2l8I5YivkFVepBHFIEYPH0KiQHMIyiDVVRGG4t6am4qQ7g06rSGU7Rhh/F/
TCXTuwVCtuVCe23wjSdyOS15FVeLsQX4AolBfedjeZaquMVV0ocRWSCjrMVqLeniAPics+yPo+Mi
KCY1ki2G37Lfy4bRwc9yviDln9HOp92b/a1DUyhWRSXWzUxjmr2qkqvSUqCu3E7shxYJzZ0IHUz/
9Du+bOoj1qjlRhCTHw1yYoIAAlgU6wLUY38SnvmTuQAUk2KXNzghpkzyPzpODs8llXef2o7hGVBp
CgqGPNNOWyJIuZbNHp6oUApJMEA8J+Zv3m3GMRVcy559xLt/g9DzSEof+5Pggl+uYPMoHDc5yB0B
EIGZG4QL/njzIhD3YmoTQJLEOfj7wRXXjZU7/ods/Io3O/W0lz96PBjizo4C/st+m8PJwlKku3Uj
FMCnjMpdwZxRjzDpvrcEHxtu3FWn2cXDNafV/72eBIjLG/l2NeVNhntCaiOE5hGVxP6iMW1vw464
bBcRKrXgUHiRWp1D0tdEGxegJSMGhLK5M6htNlzgvpVePN6LH2VqKa2HctWJYyZHx0Vyr9a0q2CP
zpOnKq/JDNAYJ3xkBuIhpc9A+KFAq9uoAGMN0cFR2pE70qtsLKqRn2JzGD92NNdhGGPT0/uc7Kk2
TTim2yLdhJn9RvVE+jH8+wy6pgEkY/c5LzbIqsaSO6hCONG6RUcn8gNNp2vL15nLI3bTbFBI9SJC
+gu2dgQVvj2l/uIF72mu+7oh9hPD+rxo3iM1pxp31aaKpBae6h4TDWoIsgCWiz+/y+72JnZaL11p
iqhNPZRivjOf1Jwqa7Gdh31D07no2TnuDZTLLS7Hv+ZtY3v1iyYwMyt1fx2wh/gXgQtU2j5IMqco
byikrIVY6zLs26Sm1Ia1i+Fc5jmCPC7bKc82P5RiMD20/d2B50vfkzOd+1unpTItFudQnh6eXBOQ
LTWU0/uKXUYCTgwIv1WBbXLiDBCIY2PNMP6jNbNsYXSv/Sc/sxgxVsS40AY++RnYNH4KYKRAg4Pv
XlSAC70mFdTDqrvl5bH393fxxNdTGLrEBikigeT3hghTyR2XeUbx99XcRCUz4ZAEOCvbRzp9b0fP
+FgaxdrJz8KHeWhJ8EHJfugMvsyfjJ5zHnZVjXSki4Ydb01cM59MTB9Bzadf0yYVYmsEC1jiMz2U
z/WFzKh2lXbodp3YP5UI3T5zVEhbVsdGRTZTM3FatUS9Ahg/wpFT5bLbTv746f/u97erciK0gO5B
U2A/+PHvDQFkDzv1iboi4Eac+0zRqHvejpP3Wf/WSLSBOLVjd2ue0WEjLdjT4b4+xCgDERKNpKrG
8NXb2o4NMel9Is/4Tox0v5b6NZzRBfq+t41Ww9dkxgcCsgTwn8gdGeskUXTmWLe1XbpbwzIQYTVu
2wKGNkm74oIQeRVIaQUXrEExoLVtauZkQcBmVd4EzGyeOtqYgLC6jRGyfOs1xGVr4Skvf+cxfsBr
WlV39D6NS8nRfA7zJVnCpOJ7W2ApNQGkTSbxhFCn40RCZ1AniaCOgXixRQBRyoY2RIPxqqTrQ03S
y9lmJ01NNw6C+RmJIQ4gvUekXbzXydfHkDic0qg3KIDKyHBofS0pVMXL/FjqsVFMlfgnGvfq6+pW
elTpLp+bMQhDIs3/RVA/KUVyR027XZSfxp4F2prKUKtH2PyzaNgxlCxk4WrVXkODkzcc/KBsmQ/9
a3nifoLfCZc/DM3ei4RWaE61U+B6B6W+dSeQN1f/0J3IfzaV3iaGr97CDDiQq/IRzKFGGpPsxhtE
dFdbSoJnxoX4ImMGJIbXG7xKg8QPESx3gWytoJl9SNHn5Qt8MyRHxU9s2fkFJDMvNlVh7sSIwZE7
fxiqJ4LkrhaSartGeUp51YPE2+L6cr22dTMF6Og9c4u0HPxz8KVvtz5ji0ZSKVIuF1YjnOmKjlgY
p4z341NnGvdh+2U0kKehRByouoIodPCiR+Q+W+fnkULcKrjHWBoQu0UQz8ZvgQjRLv+2VFfx3p1t
m1BWF6eAOjW8Kwoj6KIGvuu2nM5v3s2Zt7za1vzIuD6jsMsQ0esG09c+FW3wUUa6fknowfOGiCmH
DOEAV9uYiv8z8QNHsqxROwnYmE9DoLnEgaCxq8PFwfJYnoXFHC0YxRd09xD5Dlybnh8XyZMmCkQK
kT6abOX31kDErlNZ49s0TMqQGQrZEOsLyQhDCT46c3rkMoOlGAzrNR9dYKZay0DiU6KoWiadpSRR
YwN51tialvpaQ3lCvTBamT+VT3QSvK7Z7a+We1HF5TVZnyp1ZNQaNkvg7ZaLXzXyFSFbt3pPBDPe
L6SLouUCf7dQxwTd0ZO+RcEw7P997GvjXqzy1JTKiO9BZiIENKXBU3ldP75degA38pt8haNG7oTz
vsgW4bOJs46aE60PwT1EolzBU+fsB6x8ub514L3ZxJ229MI2sCiojyY4f6gts3wPGK4YLoUfNpsc
4D2dpXEpxO1aIuSNdFNfyvXZFwUS2LhxXoHPy1Xu20nATkSgllWSWokNB2/KYByGcR/yVmoJ6z/Z
yH0kT8ePYyTHRuL6v5lh4IzCDH7Ir16Tu6NGkN/4b0xlgFUAWrDNOWdaOD4tfzzPE2GjT/lLU8xM
38U0BfTGIKhH7nuvgwvvmyuHXCKCQqnMd4ZYOjmsigiAPkvb+kd7vGGDdATIMWaDZjXMj5+W7G0E
kUpuJwvr25y+2r/8O5HMp3T430RBJAkhBnwwWkNRbs/WifACOsvR8KcCPlaA3zstKWJr8NCzejJK
Xfpn5avs62hfaTJA4ehIOuay1gf+MMPWWF8eXNyNTtC0BH0DaC7Osc57B8puq4/HnWvpKWx/1jIC
ERfSxSxkJJPlgexwH3UesE8dC//GCyKByAbHmBQ+IadHpWZHlbnYlT7IvUqMQ6XMgRlvF8X0QtbS
wAGLkNSO+0HPSQNcsdRjxCBjTJr9FGAlv0E7fQQBbg1a7Cgj8ltx2bk73KI8o8QTS/HGghklxA7t
yxnBKtrFLYb6fl95cKeLLb56lN1/DTk4gjWncG1q/rS6o0dEhmwA+GKL1x3STH2Qx2l52syQNSEU
ZvvxC40RcZByplSUTBGMnwirrWMh5RWVoJiE3y/DVYoOUCUzY5gOUGfZ4Cy7nBKYJHbVrCuJx6uL
01x8WCc4L6UdYq2nb4DLkA+19CbJPzesHbegP09I/bm1BFt3RG+Sl0GCGn9kNWw6WuXoI9Ci7xl6
Lev3NNn2io21AwObfCYcz43kOMeUyU3J+lP/y7iEAOhYVBttjaY5ByyLFlSeYgThR16nfbA+85ni
AjDmIW56Fi4fE2UqlrmQCrJ+Wze3unYPrrypi+6/8tngzn9EAaw/6UtvDv22DwwsdOjGi9Hip43o
OV5T8zdLmfc/qkdlGqu1BX2q/sxBaRcLkHxOixSiIOvYqqbKElWvXg+oBqpXz4fc+XlRlO5i4k4n
xqheFqZOszhL9OxKfn+CO0dTdwFuW8fPipOb6NOphG88tTuGItKKOltdArtJpSiOJiY1GtX5Lyv9
VrSqGyNEWa2it0r2QeJFt1R/l2P8evMBKpCaJgQxDGkN2Z/2Vzl/ZiIcW32T+uajagzphudLyme3
xvglsvqFM1V1eJvteNweTBEPU0H4z2uMkbpokVa6GKxiTAtj4Q7Ix0J4TZLSVlcNDwF/BmDbJuE2
9HFVp0DttbYaBHVmvPN7V9RgY+yxwIw4sKv8bKnTDjsvPjj9SGolWgTd3WaEjG69HfYAq7E8J7US
nB0nQRRMNHJ9zC37KMZj9eiVLPBbgy8SNVKNYhdFXwB397fHsLNB40rAwOLfIcDBJBXxXJxpVecH
+GHbYWhhRF0T5URmnhX5Ai928JNY4bD/yRJG30XqXPFx+19H/2tZZVt+jYzdL/HfixofFLrAaUhe
CYeHaet4r6PpkmxrJTE93adbZ7U37rlUHaU7ZiBRXYWMmtEWWbbu2c+tD4MAXNSDDKylisthV4Ny
usfI9454IqKKSt0YHSYCgzScp7EAQID6o0YA3djc7/dppN0mLiYTwcfDSQ43wtCNntVuRSzYtuhe
hte7pAHx6jjMhkI14pdI1tzK9fU4zYF7d6cbdFVp2FqFrM9ipgLx8/Y68bkkQorlzJOepBiej16M
WxSWDa9VZv3qjywuwtii1pG+0+ruY585WpeBnVc1kkRPEVk+gVHO5rCwBs46wQa1Ribkz7CHs6K8
zREQyNFTfbXfXkaQx9mPKMII5Goj9/KefUZJkbUQnJ05vCtA2ABU8vqzd0Zsf4pR7fJBxZnlUC6V
Rhucva0VdKv1v2pMyny7lKk6OhsRT5L0xSe3MH4aqZwHO3EY32QFg5hhMQWVaDykq77YMY1E32gM
vDEiG9XwP7UtTbeT5ozZShOJwobll4rDkthf61YlUfCClkDw6bI61npTqWtveXVJV48Wqih1ScaB
Aa76cSntIppuuW4cS2VPQAIVr+KHMFCLBaPg2xuvTUETcFrdzpIJut9BptBwehntItCtFWRjBtfU
J3MpwssJgYuOhIgssOAjQuZImFLdewc2XbIfKbj4IOHqbMoJOdv6tj5l3rGCjP4qQPP/M2SxEWV3
YYMdiH36R2v2DjNyqL2aji1wGXJnn9UO6dm7NOxxqSQH8x561phTcdKj2toFE1+vTa0JLpwwSqM1
dkjURuDXjelzk+aFmqJVp2C7A893Mdw9SRy5qQgxtTFGXU9tKLxxOCU+G/8KellbeaJa7CCenzqv
GLMf0EysoFjwTHTEbWFPGibm/DMCN8ZAxzZPNiMBD4jUmDPtE6PY9S+Rl9hpamNgVg/h3NbpGirb
iRDIl8BWLWUYdI4ILWHQ0PH7QCoaxKnm4AvLSd20r14+SJwo3ged3g8K5JvwuJ3vlGSYYSDfrmSU
O19/UvtVXyYHB6FHoq3WcnkUndwwqG7FCOVYpoFoOH3tAW7CZWFfhqDIekY0t/Qeype3HkfYF4lM
XdBW1aDWITEgOc06BKsrg1KdtfBmaTwLVJECPYAy+d/wyUV29eI/xJRYqIWvfjPELn2TuI6pJCkU
PxZxo2f+9MwitF/hc0Kehr8zjC9XxRlmCZTKbSzQcwFiAZSnwIfZN6ZglasHjtjLpSjFZfcR0f7t
lxhgFa+MAYDs3a1FjQI9ieuhswDBE994gf9noQYh91OGiSKYfivryJ0vUhZUSlX8dGmSGFlxBjO4
1NuA2/EVLndopthG0VAfwyZ8O6wm7/dv4GWagL2SiXExF5jnkJ9sVETfJoWHSURN1BtjNzGUIeRO
HoDN+MJXvkZNC5/zPxRgIjte8ka9QChxttgusi57DqzaJpeA9lTJOz7L6obho4zKeEoUV7iWj3gE
mDmGVWz2ff/f+XYL/OR1v9/FMZOoKkv6L1ah23157Hb7+BEjG1/jTPInQDxn7PVyshxflBcQnOQn
lUji98ueQ1bQPVqRMx3crzR58orv3ism0eCYDeG3uNDzg8xn1UGx21BN2Pj9qPfUeFKoS8RbDYuJ
CGU0H9LVkLYmoXJ8KeKIpJ9JvAXbIiQFeKOdrTl5320XtVjT86mZL522M4pUDchwLCqL5xrJmIBw
r2l10bHIT2GsMncfXXW5xp/zUClf7EVYC2IkdXcwCMJcNtk/sKwFRNv096Zy14mLKkKOgBYi0RN8
BUhNvHRTujUXA3cs7btpHUn7AUVxUcvTHJq0r8LnX5xo+09Dw3uPhyrk2s/6lEcEEglts5YFhlCn
/dyPLyCuGjd69tXfIH7yNl0cC10lCqvY6U1kms0Qe6jse5lQevYOYRw+XoL9mDP5H0Kuz2kO/If7
aXfEzgDG6dJkCET39N2SzXqTcKAjr1JQ1uUTsc+UBSKY8swhNKYO84a2KlMLCfX2oSirWL1DD+3t
8PxuLN+YFaQuegZKKlWmZ86V7EgvPDdxG+dUyHHTz4zhPmQ4G1S0KLaYpGkTaNrbwrR1kkxZUv1I
rFykLkGhFr2nOis5b4w03k/D6O9oYxC8EYigrWhM3utl2XZHHctl0XSX6oIH4wSGgMsezkFUkm/p
FVc2SdE4kXbN0t2T+b35HFS/KrIvYD4GYvFNf9cSqBkNUSss6qFfldeTb+8IxG7E97g7vFuRKUP7
G1JFWQ/Jl7FJ2KlfvuaTLw/NRfnTb/FGVm6g/2N2tVpMIV804u23Yi80x4hkkdur+PZEZ1+HN5hn
8QDpjfOXgEKxDdfj9gpBr3x5tko2QPVkw8SAEjhQt+RH4S+EZ61Bg5bNw7bKBjua5E9gDWIo5Cma
8pLi1B1IdBPizsYG5Or3NbMT/5L0o/c+bcK5mwndNEvlEfe9z7rbRel/l1JVvEjiNFPMfu+HRscD
RSbeNj5SCi1K8g/gvYKgvAzLDlEs37xOGHLT3gi88uIFtNBfh/L7o+bw5z6b139aOr4ag6OgsYp8
gLM24nfMaoejMFC44C3cpuB1l41L4FI0HgoOL8PqHOuHLXd+AYZBmQ232y00V843gWTjMT2USGwc
IBbxPcpN8ppU1+nqUP1fZuc1b2TDa2uTbcJL5cRB3zF9XTE3CLF4xqqgkb9tY4Q+j2wdPVOSkqAS
Sp1VZbngqr9Wt6j5NlHZ5NXHyjLQ8xxWIBKfHl6s94CkPI0hwYi/UAjRbEuXNdpufWKX5lhJF8jM
PkKHVqlmgdhB35PIVlmkn0IsCGW8n2hRzU+LPq1PxchMZFZdEBfWm98M1LGpIbTf7uaC2y5r9B9f
/cdFosaZZd1N1YkRLWFVlmtXUtloq4kmlBwpOnq+BTjsyeBfqAYNAAq7Jq7hHdzqRbxvnOkHcXfb
AWupRbiINoqhxkJsaefevc75BTRK4zN7Qwn3floC8tDJZaRIgL5fEsqgI6Y4fiOd2UcckMHbCMNk
gze2cvek/jB6aMJTrkqtLw0EbmCSLI7vAvV2HdMkzFFCGuADVoB1hqJMUJyJs630ZcAC4yAX8jwK
BxpewQRR/z1FeEYbxG75L5wg+YzWZh+xnWobSvkJrGLpxwb6TRYl/XHF5HW6dHSiQnC6rvLJpiT0
6uOsPjS6RLPtGtNuzGOg3VoiVJWG93TxXLTPnsyeQA7eicEzMtLaGBM/PfM/s7EGniVH6/DLs+Sg
OU+mUd8XxrqPgm3dIW7QKx+VWhHblomSRaWJcmTK/+n9Myy3wa44OG24olc1HprM9N3BjMGk/jgb
DSLXjCgT6UKpVQYnL9uOll6z1/EqjqNC3lHCH/z1eLTkIUnHktg0DeyrCnsqX1weAKpu3UEKJSrZ
28zKxPx6QJxvxlyKJHxDgCLsimjPkWye83/TkeYH3Tzg0c/HedtIE/J6pV7+2OSSaM3OwaRYJyAx
jHM1gv2XCQkN7BfX+kl1Wt0YKhh92RMU4Q4ix6ReScEOnyerjsIRcxk7tm83cqAAbeJlDPRJB7fm
/Mh5ojap9sRzOJ5cOA53f9o9guidVVy13yanXB4Yh7VuAuqYgw7RTt8CY6XFHrSIbZwdnNViiaNt
nNinKCqfxkL6VggztWvyfGoSyNf+W9oVrOwFeRhjWY8gAIEbeSWAnd97vVIbaF+Y6quZwYi99Frq
teWQ1b9aqqk39WXgHjHI7/IErtjIfRZ9cvOlUK3OY9OvfnR1HmrgWBowoVR3HkhwtYaCas5gKtKl
Zbv215iXK2UZXbuTNW5oqgm1B7Gnah54VzZjlyyFagYoEdCObN6Ye/3EtlpH8lbzxyoxMEaZ+ROR
EQKXOoNxIPEZan502Q9rO3NipSDOKHNrr554o3AS7EuYpF6Uki9HR4RxOwfwEJ4YzbQZ1wWoy+pN
WxVSMcQ3nujESnAiNCHPKmuib//Cxa1TbXfMn+b1eM2a7aZVCxdQEszkE12OTQTEARALEhFlOHxM
2dY7v7zXtA9Tb8UldkbCyyQax4025VJdkTGNlf76kL63lzf0SA6jCGnf59f43z8mP0IlNgwjk3nM
GPNHs4c9xDhrHocmhOxgaTCxdDvmVNrhsQ7bPN4ORAGSDDuCPkMLx737cNXD33lkj6fR63/hsdKV
YWhFRWmf2W2ZXFBOU8uCydMN1y4sgRxw3NBol0uNT8ruQsPlYBh4U7b8kXOQX5F5hRXg4l77pt5e
Bic7BrdEwh0go21Gl3iWof9Djtv4TDXNDWZpJgCV8NmxAJfhZkjeoenENfxjDFnSwfdYQ2gqlDx4
pbza4tKoBPVg3nKui6aN/FUZW9cL6l26nnj7hvrvU7qO/Lf3qf/l0XfND2U9RpvBLP4UjFejgAlp
tFnnScA38bV12uKzQlqp82vtzJTBIiFk+eb18B3MVh/ZZaX7DicU3f20I28XuzPL2rl7DMXQzHvr
PQLa7YMtKFG42g+07mGJ4yyrrFUPb6XBPAF+B7F8Jgj83Lmn49gyUcpUXWhRVIsORqgzw+xx4J7X
ck2Rcm+N+Fit7/yh1BGnD002jIWNTyeuwfHtjRleT2dSOxBfVSTPdjw+0SSdBTwqSeRgLgnaR0ae
l8+WrK3ZvnZlBpYHYGQgZ9lw/SmuN03KbgD9oVgj0l40AN42YTLYLmVUM9DOGSzwFLOWfnRtFLXR
QrP1jlo4sTb0LBR1UwQ1EoS/70OSj1V+UfiYZ7qNtXFmGxiLIG44vZ3U1fKP5FAeRzxzY++lUDpI
3xt3YWET1h0Ia5Xw27VvzKPIOKLDK7Q5SFIoAjnFd6kGP73DHX8/4I4fmyE2NlydBRyQE0pWvaHh
jebpkJJEIhMgUDY7JwDYbiYEfqwweNMaQeDd/FjmXADS76LgIey0TjqQLlwlkYY17DPzB1jz7qSy
X0bbTbWlD/ZFWnx6xouJ3L0kVtydtu6mmKuog/N0nZv9sYkPOPA61+hXRSjyBKtv8Kw80vmhAYN3
sEPI1/1wlU2xQOLdZ3b5h5g2vwC0S8C1QGKGvHvzi3PyXISo/8rz8gnVEeGUatEh5SbsMO262SgM
KoYxFiOD2ucqZFelOoIXkhWon8xtp30q/dW1viouompmF2GynQMlwycjuZgCvbAndqn8idUfB2yg
RqeALhBZWxAPQm4qfPtpHwuSRVTNASyGO1arswH7iWE+SFzYpS008wNv7tClKCjrj6QiJLaMmsbh
02o+YOwpraOSw95irZ7ne/SGcpThDZg60K0n7iGeuX7kxy5BQgHgLLJ+O6ZRd4cZWn/A6ZH7inon
7oe0/83Xgf8iWrOTmxSL5NqOmoUUmxkwhdKswFHbqTz8Ak8xFFWzAFuJoDVprs+lf3D+MhX9cQ/U
Fkm19YLiUEumooFR44lkUhClRa8sS39DnULGZBfg2ss39Xiic6SbVLoFaaAktXwmAcEMxY7brAph
eP50mMzTGfYUAjV5nRwyTbENF/I6jZGYxoSPmFQ+ClipEdOL6DQShwEleUMnj1V2kKuBpLtXsbNn
vaAsUFga7ecz9jnjlpwLtnkpti6C+2SnuHDv+p5Nmu5ScjvZ/BmFK0+X02nP+FSFV/n0v+qSrQ4L
JsqHqLoV/oRuAlafWZ/ZWd1rvGNjv7eMTdonQmz7EgE58qO6ZoPEp2FJN6mhXjjpayfsJ48tEbaS
YEPqpA4vWfxp1Pso+FYhWyqY9HQbWE9vXzO5aM0kMvp8T+1Ja3UKFIRMJRaGTG/Upd5voqQMNpg9
vQ6yqjXD9vEYFUK7mCcezNqmprwoXtPYRu8/7nuJCL+pXBYO/65aGg3vqQejX9sIlqyPru8fJO4g
fbgpOPuQekSKD9nvijH3B7qbTdnpnyQ2ZHw//+Ug9p6rW1gvizLTzp42e4D3CblfmWOmUo19PBm+
c3w8tU3OD/Yj6qXgzM7DMa1wgvjVrsQS3LfhW0VDQuOvoI0waNC627KDtXEAFsgg4FT8zspg2BcL
w8m0h0dBzpO984AbzAj/gXilGjf/cswInyYX9MjB+Br4R+wRfcctk65N+QJKwuoUTqC5QRM2JXAH
2FRYTYttUy2902Kewafo+LJ+F4jaHJMSSOz8QRDB/FKV80BQ1C8Zx23mkyT0hnKY5BXAmX33PlVP
ojfspQlfY4eKtTZpdJ/7aEgvJ9Hrvcau/zuLLsindcizPj77xgywtDb4ybOM5HenXwWRHTQAuPO6
LO+d7yCAVENYym24JmO4ZF1piognG7uUAwXvSNee/c0pjiPia04cxpNE00VV/0Iywdmtpxl+M3h3
8wxca1Pl2WwLQNknwl/BPkk2lB0xkIOLngbuEEDSYxdbX42hqh4/5NDKGzgzrZRuJbKSNhVVcdsF
xsQw2rbBoCLeVZyEHdsWqsxTg6fopDV3Y6dxmKC99MF+F9lTxd/m12cY7hr7zdzVD6r9+TsYbNOb
nnfq5q0hVbHEB1IAP8qUd7w5vl86ODzYHSVhE5sXm3VO3OSb5ZsDhxyT6Vlh9IwS4+kCPahDOL/a
gjsJ0vBipjH1uV7BL1p4RggOmA/+9hkQX1m+tghEx2PTEM12uzqSnGRY9SVCqqMBnanzOm9EPpTg
2zw5Ajf0Yu4qWQt3MYfgV0G2LXJ9YlB55Rvl+BhsPeaNljAhR+txSQuz2z5Z/YzAAI5/MVSs7YiF
AwYj+Usg7gSglw6boRqr/q+LAQTYPxiKxO+FrLhWoHPvng+raFHK+L7fJFX49JY8w80J9QrkczQy
lx4l80MN66x+l7W43m4Jjosd8uRpiVKiddxDW4xl3mo9CZwJ8QdUylsyL5ajREq+OwzgUG5Xklxj
SoEDU1fJaHEwCmZwQ1M8nEx/gsUrTXsMONfjQLZz505w99HCcZYjVbNTPzI11gV6kBAJnrmUk8Kz
01GFg1To9YBF9YN7UFgausn/HVf0fncva1/CjjrucV+XTu76O29E4T7c2nj0sI0kYTfFL7822Xh5
50aeMtUZaE3KZa97iva+IryEZbkboKS2jqNwNjUqOfhaUe2C/bqcubdszS3gQHskKVDmJ5ibIid/
ZxtbUq/UXW0wb6J152yo9or8Q2WUMlGw/My4qmyncdiQFyq+RPVl4IVl1HDjJ++mbfy8X5IY0pAw
pO4DBxLCPtRFLZyGJY5unExgQG1SLGOl4P+w3woWCv9Rkhwop6cUhD58SO45XHc265VX3lpVMlP8
XjtzBuggM2o5QOntGgihM6LerwzBR854qDcclrZwAZhc3ZotPi38JERI69LcWR7gkCVB9eusTpKv
i1PwMNfwGGCCBxEYtcER3fyEJ/avG9EceZSHCR0pKHWUh/LPx9uuP7zEi7OyrmHHYpnkhSfOlWqq
JTF6+50UlSPToFak3qSjbwLFaNpUns4AylEuDhB56itlHZ7G/y0zCkoBO6BBVDDmU/NV6m5NpJ0+
hMPmLK4v+aCoNhiwKtudmy230g+tFeg+UscWsAc/hFenFdC+c4nImdtriDpwgsEDaJy+SdL4g0sJ
MHf7v+8q/AWrbs06sY6N+eBzSIWIo0ZbkNkd+0kbzeqTf98Bxno9Wg7yJAtJF6ZBNpwi0gagG/O2
4XttrorzcR0YCIe8zk2PzpEmlyjJVct81c6WAIYC1TSGtfHXZAiERnY/JnBXJX+lW5W728FTFyOw
Dxrc783GfHMYlBIlFROpuZNVWLp8DNv7IxrlIpB8h8hVXmp3M7657ZK2oWgkDTfyMVWijmKl5Wwm
ghFn+yW1iTwYHhopr+IvhOlYduum3rSaYaZfHHXYvjslZjuYlhQxzd8inB3kfezZ4h1E5BUMYNNL
+qDPMMCCOqagzUGYzTEZENJxWfIl2qJLPmxU7rkTDlDfPBC3JX80bbLk/fASAnLFFttHJbvJnCdd
jqtgcMdDrEb5QHN+70DEIIJv5h1luVZ63QNNd2XTYzpW8xJ6s9ZOF+JCDu5Qxvdu5lL5IvWcb95v
xrM+GmGOkbeUjlau96CIChUSfw/foCLf5F02WTS3CXNW6PWL+R5DyIBSFRCUturwUf65ay3QRH5i
QIirxUUrXpN6vYnSuWJpD9CGWfq0NeJXkddsqf4XsYY7/6xOGtHKMrMTQUuy0MPrsDpdKb61cQ3p
vtPbFyyCquGomFoJeixbB1PxAZtQvLY5lVCPLsjpHUnu4HhCaIq8rD0Q3cqOtDm9rimvNju1RaLm
x37uNwMez3VMCpNc3QAs6uUVi5c2jg1G9JEibXw9gn0tRL2Hh/5qYSXAqXGKxuDJ+irpzQuY81jm
VVldQ6dQsCKRsJ0FvHGxS/aWZpjK1iibW0PRKC//6hUhdvqRZiseg0ey/BY0/WUJvH6U0Btfu1e9
oMffBcggnePTx7miNvPSetISL3Qx74mbUfG+gQBuZggxalEwelfV1XkqjvItyvKe/G6o4oDiFmcZ
ljYrUwgStdj/TI4p5vBO+WIZTnifEMK/63jnHgBeCxL1Oc6UlFuzoggMz0OAPNbw79XJLxpcXkJA
tDc3Uh2zDj6/ioQU1lqrWkG8gw2XIrWeqvAiX9x3E8RrHUrA7VNwNUQIrfAc2n7v61ZOq/GIQyNO
8bHpBjYWOdVGa51mMqJUusJgSs/O1Wc4R8ClEx1axzy/HCRM5gH/p3cjfatGcxd/yGJ9u3NC5CYj
hG/G4SWoC6o2cnIJ1XoGi793aUokxFQfL4fmjSoRrfsJzwA3e5If7YvC4o/13PmzdqVod2i38gRI
4XP0dkgCdgtNI/quKkf9qnWfAMR3Lf3ecOhQDD9YMYdGSdgcHX9J4IwMoDj3KStgusk5JpwPrOWg
yN8zq17RhB+k3SVzStUxqdI51kI1Kl2Frcpuaxy39bAoRiRSY4uVNRS31t28+fXH62/LVHRkKKKy
EIeVmPUwR+IttxRSb9BIkPhh35+52csINbNahfgnxzm7LewKyPeppdQ7tNynub+azHYdG9j8hQHy
gYSbjM35RhBiux29TaTOIzal8YRClvl0Pg/k3knqNF/EGsx0HhhJbGyBDlozovIpjhg1R2f0vf+Q
txZ1ix7ApM7l0XZxmbHC5JbNxY0Wc0JR7J3/VIpZUYvYR3294Y6bg2kZgjDea4tP0s+AAAFL+OIi
7cgzBNSib56GOJwptr59dSfV5aJ04iNzWAR+LIDCr6BudLAmxJsxA7uN9ftdIwng1Sx3+HLvG/82
qboNoiL6rSy3PodZmqjN9MLzlnctxihOJL1DydO9CM7uuNDw60CdX+hwDkRtfuounToTGEOVjxLw
NTAipCmQeDzogX+khZ7NYHgNG5zM0WCPQBx8EJ4YLJNYt7X4cuY7P8E6LKbamnLhoPI7WnUQtZXM
mn3tKK7l+afxSJeABFMAyRhHqUpAYsTCmNL/AjXezKQMnh0BuTsUzTnTAX+a/X1VH8wJm7PD+sWI
AuLIx/UCmhJxLt+U2OStOSKgIrQGQbvmRFDAmtS6FIzWJu3oo2SEyjeMUTsikbdZUR4/avg1QGfw
Si0WmJRL23xiGd+/q3GW/e25euUrpiBXGWOQBwSS7XgBMTfDhw9XZmTrqJ3pnU45jvxhwO5y4HGx
tu446ZHMwjDHBrl+rQMbwlC8CAX5YEaqVL2+4YEPp1mD2ZtrfOse7RiSFarncxmyc3xlBFQ7jOoo
UU738+8VvgF73QCfMCQT5Z/aYQj/sxqun7vgnwoqc/RJQbU38BWn3xGPSZiiNmFnfYjMmOdibfDy
RlLA5HJ9F1easQpFIgXzsbC6M4uYUYLxhMtYZ8iUfdUqHffzals92dA/M6OqBqaX/Q7vJnkxDPhb
nwAwvhdjc0aPCRow++mBhb99naBULRPhJ9ZHfehdIIctftrKDgJkCg4KsnnlzWkKNPm5fXmpbEcJ
tDPY/4WHkPZwMfK8Eb8VevfoH5RNn8FDqG8di83G/qD73DrEbygBVvbwY9QZbIMIhNvz806lVrps
0Vh/Re2+v1tG/kiqkXIH8D7DQy21zyIUycUt0WyDv9a9dkbo448eE2DDIdyQ3K8lWOiyUYK7GjCG
azJO8Iv6lWRFUwIN1+whSzkwqG0ESdJvsXqFqpig0cLs1oRgfR15vG6TWRaY0s1GegaHcvAh/8CX
Ol8nGY+SZ4uBE0dxTPdR7ocOd1Xnkon/I6pQOhwIxYH/4O+max7t9/K8OO9+ZhmCaROfWcbvOOfH
HKXBAJtqGosiXqmp1duG0guJqwn8uFYp27XdggkLFwn3waDm/6haCi8H3c9WASvUZUrIgFQkT0HP
/cVnNexh311LCSoQ3txz/o0VQ3B9U205/EErXhLeCCpLxtawqSH4h7wpC8fZ4GF7C60/60/QCXcQ
U2HxkYU3XL4dA9ufmd79o5zTlBXyDebUsTYJwZwc1C+1cYri4jEJR6a2nA9wHSG2HzKAu5RB04Y1
IaAYQmgvtppegJQABxtdbixWg/Iry3iYnFgF9m198Vxve6vEjud2pAR1UQFZKuU4OXeKIqWfdLdq
YXCyck8uIRo74qYhB1Wjv3seIQUwZaO0Epp1uypEPG3L6/PQKajUyQ3JCYE+Ai3VuVr7g8fcntSe
H1T2XaHwQXnAgtSMI+1dsKoELPozweo5BwEcuU/1Zxv/6sE0dhxLr9SkZAhR9Lqm9/Pe6gY7rqvY
qDd2sPh92KzN7cMq+WfXu8A4TNyacIlJYibjyrF47wf0LqC71bm4w1CIRPO67HMQP+asdP4nz1Wi
KXd8DE+zVEy8OPM+eAL2VuOzQbkudSujjyMBOPlNG09gVOGd/F3HtusWB7NKgu5VAZGRx8S46yVz
NnUxOHSYlBGUGqK5Vc57DAHeIx3YIfegPeqLOtJ9HnVgQNCTaUNHEhEzGufPkLSKBewaMN1eTQTT
YO06eJfTzqmxukji7jH/VdruurJKPnx9VWBuc5ugGJsxWuD/uJsHpM7iLpnXDsfQnzhD3KAiUg/R
9dgCiXh0yd9fgv/Dz1OqFsRUgCFa/M/Fb/DEqsZoRIN6DS2qNQsXFNZ5TTP4vlEoonDoEKt1IU4t
WNulmXeubva+Mot9C0FpCfZRgYAC2ySLxvTt07g0F8K1bOfGeWMxzOHLolWPwuzrkshMDA2DBnGq
awyHXM8eums8EbJgWONBFmK3sjGk76rC07+aRdARnC5IlKQMFrQn3mmCPieBBdWmMohv591G/8Bc
lNHAoUJESJvtdbWSBBaVcNNrvEQDUnHN9wvnw0LUfKEDV8BYzQSIOQvck0ywvEwFh2s7tg3GQqeP
epOvKjhsG4u6OEkqD98vM6k2EyxaYJN55ALRSDC/SHfk1GRuLsK3U296kbdER/48rhQsVk1JVdNQ
FvMg7Qz3PIkuD9606tqTIkPdXZINZu5aOdTioOd/ruGFZh8fJCvDCbvSzasFA/Dnc9WUR9sZ5O2G
nidJ0cy1nYRNswCFltXMS2jfZDzmICEFkCpmzkEYD0P0mHfSzNLau7d/DAVLW8ZWtjVzr0hEDwLl
nnmi2d4oySj3bmDvuOUHEISX//4g1NF7HW1C3CP4Ul6zYBzw+lywx9a3gvK14+S9qYKAmGfLLwXz
vtZX3+UQLMBvGG2zJ8E4Vp5pkEjLfvh1Clx4oQWE5M+NjBVlT9t0p01LkykaCKYEoOFyvEfbhqiY
j5Tatkhp8jMZZVMolRqBjLHU32rBGDGsKedJG8vhTzjY5yRLidN0S0zBRUF6Q5AoNKwsO+2BoaYU
v6UQ60VLnjjty6HyR6VBE7PX/Ti1pqV/N9mXCk0jRvk+DSYzjXw+V9Z+0MnSBsF9thkyIk6ygCGx
C2DSbqTU0FqOTReFImeJyfrHup9SCRWUo34z+MTVGviQtTQJEzic4yVrKpstgTNz7Itq+HP3ticX
cP+QgbM5/2tKNDf/1RxVVlYlUiEAxvHuTRTXD0Q894ZWUyY1aSooT9/swGWE6rU+3Pb1kQpWNX5e
GS+r5TkDekllEQFD3TYvgAKOPNPaUzTeUTT12x1w/knHdpMxQftW/LVvWDY7h8GZ3wzFskspXD+u
t9YLVxwjJISK87qxWMcsXI3cswJFkEdAywLYCWY9ygoXbWDkrJp8tVz3pMuUbEaz1hqDQTMBCylo
p78o+XYf2iUGbIejaXmOPJHlut0LXj5tSOopCXFxe5gnolX+CB7/MQIc9Y63QTE1s8q0E3ojNPUj
hs16cC7Vl7j938+v5pEBzdysFVCmrmpnu4gUsLtWF+rmQQSxYXZySpTmKOaWhT1+SBnX+e5+3nPy
Qfq7pMGddxx3i7yDn15nH6X6ewVBSujaUTyPwvQY68kVBiZhiy+lAyYIqhRsiCeJm/pYCV+3xWpA
gqzWXNispB/3+RHOtifbalkttsdTgGLJsQ+QLVfl1I17517/nZGHH6V+jydfmJIPdfCea6NtCL0D
6t7Pk1qWi9mQPNHTAQEylmQe9kvWuaqVTNugyj4jmQRq62X95LHb9gnhc3/kogZPLrg6F7LEjABX
86viYymdcBdigQRloQN8x7D3ULBP7jon74LgMy2Ofd5f5V6X9AImqs0rZGdCZ6W4hskVZnL9MZUW
aFLGwGZxgcQozsXip/frmjt4tRjoVH98fY8OmX50E+k1gAyL4C+WuDlSHMZkR/xCpW7lOX8quZR8
Qbf5jJKVzHSRI7n1bWDqsiusMCfs7VUkdx6Vb5uXkluM1fU7g7bHlaWsburb/ld6Njd51SgdJpYe
RuFkYnR9IaKMhY9Xebgzepwy+SnPIzCD+ijzxd6Og3Qmc3eH6BcrpiH2DBLabKwgT6qfpxtE+PCb
3SNglF5BH3VttFkFJXbCuo+lrPDDRMOyVydj6nMPzgFxvfzJGIHtylfzSrLn7oPcYwc8/cIC+EUH
xcQN499NoaNZqMyiUbgX501gPiP3COjsjGFrjqbigo/58Guir1rnakPcelKlunYCDdbvqeYy3FH+
LUyWGhBEmHYG+/MIhvUQzmcffbP7sy3LvU7a1FNxizh/UHJZWtNPQDhD8S0q5MrpU/DrPsK4RN6y
xJRPulrtU0L0FFLv2VrYRbcgWk5nLh+YsSg8KeY0MNII9uV7+bffJw09BpR22BnVniLhro8Iye6l
kQ2iNM9YXVzmzJOTxGm7FncM2VF6lh94YYE9KSj/lXmSn1lB9A8XvXFC9xp7Bmm37QmvcFNO8gLn
1cscNhNVeOi5CNedHd+TqMUGpyYGefTDitMfvA/NUc8BHUdOjiCJvi5DjZSVpA8zZXVKOkEc4UoU
gxGOjsKu1iA5nRgjR3jPXilv8zvM7+WPoDWE2W2XUEsqaNaXEC5/Tt2/cMNMq37k3Nym1/4CzYqb
CqwNCe/SmwMOZ7/GyRUpEs23bym24UJqvYn1xFdR/bi9J+CrrnzR7+S10g4y4544IZclV41zG42Z
2Cfs9rGcIUYtvuP0N5becX1wltxD5mhxxilG0ydIoRVqn/9Oqj+EsgZVJBIcT76M4risgN30oICC
YRKdVsisAiSRzDSZIc5PIqD+GxHw/iti1uPQxFkqVlUAMuGTWhiRem13KXfhoxx6kxe5bYIvjchM
UvUqbeh7Ol7vWSkHIMTAFNUhsrlEx2Lx6oXUiH2rCUnOtHxt9wxmp3jqS2lVC2b9dXMKdSRDIdNn
Suwe7v8UBKCPh51JaKiDmBtdOqm7RjfTJUCeslHJSH3lyz5jND5wHiV6pCneFwFmFxu2RS2o1Mnn
QD5QnsvhLd7OMSEEJjH9lHK0wAT4PgBzU8QAGA/5VrlWXPHQ3melvoVWSvZ+e9M3DvNItN7IkiRg
4c0miR3cCq/v0rLPGOa140sgXrWaZKjPNN5wQp/XkJB+0U68YqCHLyoYGybaSncn69LJjws0Zs0H
ZAvMg5qcO3b+MDCn4Iv0dfRJVSEdL8HTDVYkwP1MdFf72EqiQZYhM6ByJWmw3uhZwOn7quqVivw2
jOrVv6/D3BH79uI6FhiIdYixsLmLXlLLBv0x+YjKG/UaJTjhmXcsmw+cYqvGDrSl90tP5Ilz8V/y
Z/q3ktksap/VwUbZUlNeW/Fthd6L3GUilOVsG45XeSmmJBrSp7yXK6psWAR2Bs5ArcJEpd++Im2u
iDAqxM9NtLjFrIVDpU+YqKOhu341VUXdqCQ8LmdZeCbDSVyyBPvIdxHQbhtQz41QY4E08eQvXqSS
wZmaLPyRzaZdVIssfIuapoiHlWA+gz9Eeu7TOp1ZgUKd/Dq1Vv8BBPI3bPqbSMClx8U4uMlabprV
U9BK9i9GMVLgPovSjy1pcufi5MmhkPavXg9KEVFwmb1Uf3G4LMEXAP8bUg57R3Ti3ILAYRzdswrz
IYZiPo8KWESOx7ctonQrNiV3jhkp+T16TXMH20F4Tk53u+PQyU1vN/mun5gw3WYUmJ52TbZyNuwK
GDwt1G2stj2QcNSoCZLITvptINtPoEp4MHlgVMpX/JjfHMD6hbLKBSE+ZZNOl9BG99FPLfUXBk2l
2kBmJ/kJ+Ktf8TiviQ5jxZToKQ85zX4M3cGb58goaUV8RImjcquiINSAc2sBPD9O+QjWBuf2xmDP
dB20I1Z0bmLuXAmFSnXQaxLsjBdUNYf7laLxkmGXSJj/XR5vefP1yeOLfBrDuMx4U/FMIi1VstmU
BI/QXWUs5Fe9HcJyTczi4mcWrVAGbOM0BzFSMScHGIXoS1rl1yhdjQMxkAmotnLJ7vzfG5obKCa1
815B8q2a3zdSRB9SUvEPH2f/ggKd1Ac2ZhrwGtj/qRnJPt+/tTKkEMJuNg6v4FtUwpDhUzh+vdgR
oAYWOUdXkLH/TDMXDn6izjrkCrp4ny+N0w27yAYn6poMTFcBmKgUG1j3BZF22h0S5KTnbu5LUCFX
bR/vsn1f/JxPHAUqrLzV5pdezYwHvduD3XPveymDFQN6/TtSiRTUizKUxuelWG9MGTrAxTAi2qa9
cB3gAfTLLiGe1Xz4rGniEfkKqm/9lvKSqTC5yv7W0lhYiuqbppX1B+p0EME56EI/1ocLEEnkHUrj
wxqej3TC+nJTJY5jkJXdD1NIyImKG2vhVw+DP3jJbaDLRXleAS4dd8H4p6+RpJ7JbdEvkBn7Tdwy
EL8we1IX0Q9sxfwKVoUZeItup6GMM7aBA0O4zG7A0z264d+EkeBKdRBHK/sodAjvZrV6omeitoL1
ERitxrSPjthdTeyMorXvMeLu4NCL0XdRFvKCFkBTx3dVYPDTdNq334iJiDEkq/7GxpV1Df2lqmg0
rpyDHYM1D61DA2ZlxmufjTcW11HZGWVNjvrDn5hYtVaUhRSPBs4L/y2HcZr7I4DBu0ni/bu3XKgb
ma9Z7b+B7ruypPTRUMsTk/UmYKI/Uzssdiq28/Sau+dsp4KcvAqHX4Jwg1yEB7tr4mturEL076pM
9XK0j4rflm9mVgbhcgwNMq9nsS0HWN5Oa5kz/dq1vTv/bDYgq/3n3+nvw613GMVxP8mG5lgiYDSB
jTcc7BlGg1UahuHcamrTpZmL79mZr6StHOXqh2isy/YH6wUia0iiMHAf+AJcEQ3ou6nE/5vThAOI
MoYqFFOKD8tcaXjoVBGnItd6PdsBWhHeIWdl/igS/Ozx99KI6kGggHrrTUT7WIy4JT8QKzhNRB/S
wA4c6yHpqUXh4OtxeLako+aQWy/2HlJ2GYGq62P85iuI2fNFugRE86sWxXbp+vkeV/jpvwfnL1Pl
UzS72exKSnkdmewkNoOeIDIolUsPiRbEZdMpAHhqCXD8yMlsMUJHqBLBidRgfs4C9MNZmHfKSm85
t0Uzh+QF82pLnDUi6NtJAtcnAOV+bfqXqJ/EqHAqNy/Od8sS/pAXjFx5lL703iSUCRvVPXuEDwZw
hYjhq7oJ7QD3IW85OCKjL4szOUHbDlJA3uJ8J5i5PWSO9VuWcs+66zBJlEzX+e8PR5chd3pGSlNc
exPgRsZzrSFe+nlJD5hZtQ5O5JHJJjIqJ6UK+22bbjH/xbuMHmtR7J4A8ikrSsdwqDpjCtt43ZxT
fpeslUaVtCgL3EVX3Fi+F2UE31LItLtM0vwB1RXD9Xse1sA9cPZbY/azeCBVMtb+b+6VNP1Z1mv8
rOCl9K5wqmb/d20EP/JQtgjY4t7/Q8gCykGOeqwQmMRcGE6lZ/HGSrbrYf5yKWmDOV8Vm2tc1qe5
BQ8EnkzdGKUMTaJTqpRTgQkV+/39N7Ip9M/Sp8NSXfYCBgPrrJ16/R41MFPZxU/NcnAAIhSzmDsj
RIkkbkqRbzMrar6UpbLz1DYrpJZXkIOWpUJM05sv1X+UeV6b09UbNFelUcNOeRLKr94nic+qaPce
4bTdLZ4kBAqIB870qMl0hvN5sM3r1ze6pGPTWZtlBcV32kYVAv33JpANevpf9qKZObjO6Ucyfgwp
QbCJrCIC7GxBZvy305hC8gd0ZujZsuhAiFPeqZWGxTger/SWidUcNgxDuTViz2Oq5SpqB0+ZIcJB
JH+sJBRdDEikX1mfyUn43DYr/aBOyHe0hdFkioc9CxLPJmN+CjQhgnRpJz3OdKNzpCkeEa62BMvz
uCFr4BwyZZHIcz7Zv52w0P/Nu3KrURNFIeIjnRE14TI4pv+gw1Kk1Og+PW7rjiJuIgzLFcrFKZel
q3gHaKDha2oDBrlWEmV7oN8/PX1sIwApnZtnhW4QUhwYsCBSfHusqlCEW6EQ1jD3FZVwvvENUh7L
urQLDLloBHjhlBs4bSzkkUeegvF9xFdFS2d7IKYYXlJY3ndVfgyo+nIhJMRhDAVsMliU2todl2nq
taaZjlo72SqAXKrFHP7prGwOoBfGiJW2ziBOEMEBwJSYSe9i+R2NXS7qM/E05yp0LLFGA8Hcc6ZK
HYij/s2OW+aOgp08+L03J69tvKifDWB8bt+v2wDGtswD3lsHuG9sD2fL7kyQGhTD2jBzupUg2Yyk
HAabjUITcaP83iTzjnKM/UL5ksl5yEVTv8dSfEU4tmr3tUYXrl6e0gjvr8BxZxtF+FODbcZKyBw2
rzs1tIFaWonmFRWWKA4siS/hSKSn2Vzg/ACexJuS0hm/QqAQhvOJyJgUgLQjHE5/IsD3YOikejHk
RSwr1YgMY+MKThL9AhwZrTvpTC3ZwQoz4lvp3LjrF+uCJCYUCs7RmhsM8J+rshAKPPRCdM7rpH3J
uPD58QhyTzhGBpXUQ2GTfQOMbaLR6gSUdjWW83eLy29PKFqo7dXY2L6/ERTjYjnQqspwlKGQ5snH
ojqPL5l5zHPKcPRcRkQRKlam8ZHKX0OJqwKdR/TeDTdWE7z9MubelkMl+UuvPOytlo7MDTbdEjdq
ZWyDG9Nyw4NPE3rdxU+LCnZt8Kk/9VZGIo63B6t0sDhCgO7xDLw253bI10114X2/1dsklznL89nY
vIdvI/UIvCW+uyCEFAlyXL0k06dznUrWLaPCrSFyuB1SST++9W7U3ob238QOtS0uvRFwOCrTE8HY
l8SVBpsLu2WaSHMNoqxP7JjZ9xubl/oyhWFhwCtS1uUXYuH5XpDqtYrRqUiWzcqPRsX6Y/E6d+Vv
sfYrzS53Xnt7CqwSIP8yHMaD0uDC8s95VKKNjdwf3iyYdyFbNiw9mU4E4dBVm3n80uDMsZo8pyrT
Ae8wyfo4+iCTLDFeWDNBTQ4ZBSz/kMl/cLfbUA0CUam9ik6cLfW2fSnRkwd4ICiVdYwvn9zuyNZs
wyHoPZqamv5YLndhrwDzByAOL82dB+NDL8lgnlZk7nUHk2Bs3ZJY1tXQnNZLzuGDZJKotJqyUhwV
tFaLKyRat+bBAHrNpfVvJpHTkehsK+JieuudzyZdYl1tzNwaOeYB+efxxgJwIV2XOLKjlbZgeUfC
U9N9qNYYOCaaHY4YDVEZ4uG8Sv48c2u//M+9ZBBC7fgGyJWMtGeloolX4nNfs2PZ/3GsmG1+NLml
6Wc4fX7ei0eZT+avsG951uRghKbi0tyZnJRamIoxUxM/k5698JQRsLZ0huL/nvxqkd62V9NuaQnn
1QT0vtfV14ap6OPAbvZ+ZarRBpfEf5RkKzrI4L+TDRVOASfTaWUTCANKe/Pp73FbGA/w547cUrKU
wBB2d3dPWG8370Q2prU0zK5lbqDLzGh5xQwADrZZXq9XDCPSqlGekZr86Y3iKl8CjSBY05DOyFhG
xqXJxzqbIZoU1xNLEgAfSRfvRKi/EB9vfZCO84P3Kzkh6eQwMpW/7ijF4cjwfPlf5rMYFcBQSxpI
tdkM0ktE79EUNJFZ/LXbGuT3lyCdZSg6J1kCLfuIuwiU1TRxMvXBCwKPNJL6bChYXRmS4y6jXdzh
f8CFOsX2X7xSea3O/hDBcZ4n2KLv9qwfPDIl+XwGScKgDDxV7sbzyc5rqCX0qC8HT9GXjdljoi4E
m5bGzeU1LCd9p3yKLOzR9vNVniHf6UK5X/h1XjreooqwvbzNH/fecX7Huy4D0BrQSuV0LzT2Hc7U
tCcTlj1QPz6TnERJtSEwex5aZf9tIZIH+9li3LvrycStLqTI+1NVYwIIFvY9gwQBwOWCThsCcM6l
G5GVUkDfp6pryK1WADQaW1Svw1jt3Lpw5LM5HHDF6sa2iSEXJ5BI/LEQNhD1bqGHReBF+uJyDJpK
AAw51i1GqEtpj7Ug/WpfWvTiXJNlWwsooMpSaEyCpcKxxzluAfhdavAMfyIC66tMRPP6MxmI1gvA
XlaH6Xh3Vd3nua275ZQxbnpqY/7+ecLhbcjAl9vwjMFr0p/5RSyD0flqKi+ci3Pxrd2oejxokvFF
6DfAsqXOF2shsPJnksJjj5ZcRkq8WAh8nP922wJsPa1xrxZfyXeWW+jggYCygAupodNQGcoJM9xr
QsSu9nJ8FXc1/1sKs/05PTLc5BYZZzz+DDHXM9RAc/gGSrfa4C2fwUF5qnt+ervgXrEGHtTXANt6
KKj0iUO2S2I/YO3YOTLVRuPhI+sCV6Ybr84l+Uv8akHY/KXS4bvdOHWYlXayg2eEUuprTAEf2OSj
rV3XXBeG1/AK52TvOkROoTj/KqC73YyYdV4qoVOhVQdMImmWg7VUTE0hIniBVLeiYvWu+sBGGcYI
iAvJHFXrtzHO/ICmtRIQ9niFmZkTVe7QnMVbuF73CLjW2+OSG4YqX44ETJdOZnVSq1rqIhjDIxTX
CDqoDl/B8bOYO9RpbQzWFGWgH20SuQbPrgd/xN7POGAK5JwnfCCSeZGSfXSXUoKziluL8mC80mmm
UJ3ByjCz8a4X6cxdde4MZvyxMiw9D4NAcXwlY+YzcxXZdbIPqMVMtRClHQZqj69LJohE++8dYk0+
DwY0Y4zQu52GOcgD55liA7X/gXwk3WdiDIXg5jPZEsEgVRMzTAI1cxXpj9LBhX7diN01Tp2UKLPi
KORQ9y62lLaQPLam7QlTtmueSxysNHTlWPkg+PqudVdspTBrrn7AF8KuaCKOYOF/TTFqlQXooFei
wKH7u7a9N7FFnPiirBsXtER0O+chGP38lPeERLQbipQwZnh9w9zZmFoaPA2WQNxFa35GTjUisAIf
e/eX0v8bwwh7Q5+x3gqJ/+Hv6mXX80cTiiT9jJbLAC7pCqMOVXQh8X0VWw05uK8HQhrLLhABNzDq
xntnY/A6VagE5eHPqi3xKY4Dq8zkCSC5v7GfBTAmU5Ftk7lQLLcNfIW8oA+Wgu1QMyku8bwAyfuk
N6iAxm68Ik2zTI+XvvDvvVOowFeZ8bmAMw78xo1WTXNl0PxpORKiFp2UzzB5XDuI9wHYMB3cNZhM
7aalkIF+2cbRYcWhRaqw9GUMavRds2KrWbPqgvx3adP/vtsSRz9ov0h70ZiserTzJK6QHdmXAVEG
V1ZSefWwJhBuNwzKNeRGXoH5+Xt8bCNLci4XCs0MFEXQbbMI5zyw/TyhedizWXfnBu1PwOK5PBJO
p4etdsZlMnrnMdKsb+rJOFdq+Xon+7z0x85oER+uLHsmU5kc9msrBb8EsSs132364s0QRCEPxhAj
bG01d9b7u9ohlKdOxpa9h90dhvOzDVysFfnbF3Uht3neviK+p/a1ghvgBJ4hn5zJ09eqkc8e3/h9
RVWATshjrb16Qs4jAugrGBXvRMVkJ5O6PJrc8lsOksEtwDhCbKAOGd9gd7WYjHoDUXDFVHJ9UhPU
2wWrZdjs6jnP+M4mwphgeEDekKitLG2HEXHmJfJDhpfhXG9+fA3Thdmlsx1P02bcbNpo/pTqCXXu
V5lMHEMRKIZo60k0RNRo8T3t6LsPohuHginlsPl46eW52uVYykNcJQgtoEVtZ4G9PmUGcOb9zPD1
oC2WKERGcpYE2GXZJk3n5qJAzqYZ3iazPMuVVPBQ+yZfzGwiOvPlEvoYj2nIRFw3geTSWjtWiD9e
CxWccH8xVZb5EC4taq2b1+SMTuUEORRd+tgY35859F0gjaDrUL2f5ozKFtLfUPdBYlsCeS+B9nCa
D57YFhf8aEPnDaMY89zm4x3zjT0FyZTyIDVmgn+sDcb8+b+20lYoPnN5X4UwPk5EMktgqFXPws7Q
sihqoomaQnDloIIii76obsr0GjJ7rruMBgdm+tHzbjwnANeYs2GjIsLzc4vXOlcMhp5qOItUSEOn
/RX1jXfKhsDCDMsgzSKpSZR979Y9jTMEWR3Ks7vy9mFOCuD8Cw/aosrMlz04BDtL0IBdADgm+bvi
kV5iZcnpMz71EgDKOVoH/9kAm0X4AnVFwu2UwvLTVdTg+kA9xiIngc/2yuGlOSMMRRqdEOUNCpDf
ZEIf8BrT5AIQ5a1JTfzcsPcb8t4ngkQYR2mwcU8mXeXRGVE9T/5W9L34VCrCDXKfch/VPDDYvMfe
UgArmyiqWgjVwFXKEKqUlhZPCfBBFWQJJBUfDQL6mhDmq6N34knS5hJX4FBjCoCechEqbzyvddQ2
BpO3Len9YyWwph9zFamAvZTNL/xfnULB3oRGsEUXU04NkSpqLhgPYc0dPxkxalPphk8km56cOl0Q
BQ3ifLwxEnSeLSk2qvZdty7EVSjpEmN9z1kA9m1d6y56oSm/0q7EAqJTC2BfMqp6qKjnM+zTKgwj
pTWy8jGt+j/Gpm1eVOTBzlUjqOB2KLJZkD/XqAZTxrEwNTFkfpKQMUJl2Wux5K177r/2GL2QAfuD
r8u8nuH8xKR1dQItRBSNRvOVgRP18prOv7H/DoOx9nxE8Ks1tRdp/w1el6uWPr66vnG566dFpUGh
z2NNqWyrM4qYMzgQ+oc0MByXHQPEB8SeP+dXNBPPqV/4TXQ+w6b2s61z0oyMfwicGbw0nCEU07zJ
U8SrDQX1Pj2I8SmEJOIBSBPhLOvdTpcpNvGceqIEvXVVor2OY0gs/W9ZCjG8GKFLUjV84uOvyTqG
OWh9SKec7VHxwl2h/yNizzKtP0hWWCsk3kxUtobUswmrBffNeLqegLnvZkh7tf4XaAiTHTy79ZLl
jaN3MBCps78z/Z0a8CmZcOfhRG6M7z4PIfZHFN1j9Vb38M1z6eci6oL2QBbSbxk0v4mNcBnPAUnR
s0Ou8Uuqq9dAxlJ5qRdZRVbZ5cflXaKG8qciFuN5PbNF/LblUAsKL9u8cEF6smfJxur3Wl0tK6SS
9jBu9S0syi52cWzl8AtZHCYYhC/PRMrXlwrOUZ0vkWYsirh1bwLTRTmUsfxSY2GnG+3fo28KisHW
yuc7y24lvMzejbuglBX3eML4gaX63OpjbM9dt1cf12003GBmuxTGH4hOdd/InrTuX5BMEwDCloWi
VbaLAoFJQWYCsSWdBNt0dwGm5eg1Zoismg8LGm0EgoTY1hW0V2w3Bn9iTBnJ3a9fjXTTrywXMe6I
NVfHOIvOH7glOSPSuinHWC+Rufnbkm4Hf6oqFTlk5AzgBPfiLcFlsRoBHY53DhucwqR0sWRkgmiL
WTYLDIyuUsI+GMBZnsx0QKspf5P0HWeSjS3Lmf5iFD9/G4dQC+zGj/cX48x+mMyOxkthYA+QEC+Y
+NZKuiZ2AwMyX1rrLUe36LWM83PT75cJMk95L96dElUDJRruPZ9pOU3RMJ/ABoOd3Hf+dXJ0GmKN
Fs44Wq+cmCtwzlhRZQbyH049+0TDGpnae1YTZ48UxZwkXUH5n50tkiHQvtN4M9JySEisQ7EEgo0L
JaBEqJWXTZ7mVV4i8pv97a6a48t+SbV9vhV4af4xu1MAf4AQYt673D5ydD0CsV9eJ0YQ8Gc1fUz2
Cg24w3H5KqsA9cdKW3koRSZGja1AW8BZlZyMFgevzA/8xbI1hs9jUKAbZx6dRFJwCg0mr1RFXbDx
eksxI0PUVVH3pDjfPt+LdpV4folx1uHZPzj41wqZ9H/I+tNuvC21UsVNKtACg5KEXKyvcM6a+i0k
t9DxjfXiHtxECvjPqzBY47ItbvJtFkfSMup9vxelnTMwv97aHVdZz3PxUuUgIkg75RJBpTcscD4+
tnLlaOmVOso0tuQYP/TvU9HaZ/QXin/5kfYqtBIXsZ7n4K7uLNAhO9s2PELuA7kAlM1akg6hIFmJ
+Yx2BLHT0cdHRe2hb3728DyGqLWCyH/v+lMKc/ftxP3fzuXl8rJfMXAShm+dCHCBFFUtWUip8it1
hX7DaDY2Ir7S1NGlYOzAp4f1ceaZaF80PlnVZC+DHTXHuB5hgSLZVjyQkcUieUbQIWaFQcVaZjKu
iPCkBvPdqQ6rMM3nJ+jUCx9IRE8dVEEdEs/fpwMQ7SGnyZKu2EIkR2aDzgqwo2HYL6wtvGfXBXLx
9/SCYyD7HMI+VWXges50CCzYqYUpZT+9in2vKQmcSp1Lbo/OoJHEiUEJrXyGxnYntq5lmAi1G6/8
OpCuLy/G9XA8buL/fnlXSlEvRF8DxWvfOjP+CxjS2ZFOMUeNvXWgfe7onWdo7wXwFeNDtZaFyOvS
011t+Rsm2rXjDA6iGAmk0L8WxiUACSc2osqQG65JlmYi/5Y36d3J0baEX+PngrEAwf5QGgCLz32Q
R40d0bt/wMjLPT/y2qvCgXgnF134uWkRg29j3349x5UWCimyUS98gGEPRKjWneafuEnZpAgJheZH
AFMfr7EOnDSswWWegsz3vwvzYINK4AFkzzSXdJo16ViWkN1yoUQL5VJhkT+TdrCvPKk2WnJQX2wC
LST8chd4KPiUgjCmnURhsjmeHRmGIoYzn4nEp560ibApHqN7inkOGmYvbXaxOAZzm3cgVWsaoOUW
CubOB1k5JCILGoq5PrJvWExcghQJAp2OhOz5/AC94FmEcBr1FidZD08sEInh4cPs22Fo+XsmR4sG
WMnffnD4srU7GkTFJTWzALniPyAHG5nWbwv7P3MdtSWySlPKFT2KOnuWY6dtsFk4c1W/X/vuZPva
AN+GFtpbItCi2/+vWvg4CieIEBZdyqaotIBINaJmBPvx1u4pipwN0dKbFVusKI5ROF4Lw0FGJFrl
Cv+Q7n39krdDzlGclNgakpUmdNbNvcA7CBdozheX2sWN4rUhFHpnnECQaNk8iEa6nRLGnRoOw3CN
iV6wrF+y3yDeXHrPP3AFxN7epSMVQ8uL4Yg4sek/2kYpFHeWVmwxkloTkZJJ4Y5yPNJCsxxH5C9C
bx9tKMHaSL5Ltjlfi1GDS16qvzK7Q7aASzAoa0cN+edGBqDyeKGusPRJf4htOJ0pRrcFulpXWcxC
UCHREH9P62MmmKhHq4wGoLrMJXo1gdR7ocAMTF4eqfTayxNnA640f075l1t4d2kMi76NY7GIIvTf
0N1fAw0x/VP2HzsrWQRugjCWAd88NEQbAVKeQeVlikC693Wh83vO+h6AQhCEnGI0/kAKcEXUb0UH
1xUykE/62dS7lvHskxy5lrWgiiEEr/e55goIhRbieeHxtbNkB/WgMvoORnBSgSYZisJIm72jYb3j
S567koBQ3fM82w8WwNyWL/mORqu9x1AaVGenLpQt1uODLLgghDGjDYmtv9pIYY64sS3z7gb/D+wQ
L9v3KG+3SxFKNieZbCT8He0f5N7P4KhkJzRQZvwZrKURlDzgPAvC10l0MEfu53EUf7QUPq3bCAc8
RuBw/BwvLA0UkfSFDDvj9b+3QhSXdmhfUt20kaHEEkGo/M5bElQdGjMMrSIrOilIcatXUb7gV+Rb
C70TrOPF04roHslmmHwhNHG9opq4eKVlA5ejk+Pt6Gqj82JuFrwp5Al/qA7tG734eNffFexvgfqk
FFcxtR2WpstearGAc2zi9CXohNZ9mbQwzeK3EnwXv1dap75P17L60yS+Jup91xwTjB+i96lccFHT
X2mum0op4/w2ieq1rg0LeZzTG64WQy70SgdSd/tQRgzJ3MfPI9c/4vOQugFuABDL64bF822uzTK/
tsZq4ijMnnQj2T4rupK1fnyImSFrQbHWz7L6epkZfRFODSXDziQq52WAZvHiOKzeaYdAvTMV2kAn
WFwKh8LbF3i7j9oTEq4AUs0cRDS77YqLZk5JCRN0CKcu37HdL5JF1UtDxtfb0l/87TMeoRUBXutg
KN4He3N+cUeIXQR4zJyJ4s4gVHQdyuWjLSgqlGyHBdO352wgvCA9O4MPwjc2L2fA/hRQm4DIBSR1
DB6Bb/UVmCFHE2jq5apMy9C/NxSDZ8lvxrNCZIUwb93ifBPmfFZriu4evMxrQ6DIFqPC+BeM2lAU
WqUFNsykHSgKMozA5NVoPQtFikdI5m773VxGs/UZOo/fHsJxlOmZqaG/xJaHbh8V/W1ujleT5l3H
KUyC1zwpASkIx5w9dYVBqI1kzuvsfGwHU8oLzSHnCo7eqv2KHfzAfDbFFp+sAi5ZTJzZbZy8I8ap
wmz7EcMdRfMOKktVsF/TsGRH/fXzSlMF2MkGlm0g3WR60tnP2i0ltV8gPUP70RZiOACF/fw6r2DY
8lpuAP5cwcKqO9RQgBLWCCommmiDN81lzLZuVTkmgNLCe8K8etNMP4NLN8U4UmPA/k9P3hUd8/ki
dD6sJrt/2HWz20Gc90rsS7BptmJXNv/9G4VAxdWUwoXyw851m9smVwm19XiEDUHMQBjMsxaXfKO9
m3s7clNp/mVtC2lAo0g7GCQfUrfL/2RYigkVBuWYAlYQ5/sARuububJm+OAvfaHbv0hiWY+j/rui
NqYEcKOc6NfwXLdms4xP8xw5zBCcxd6KSYfWkzCQ3RtG3BSlo3fISoyPwa4a52LWxej8lxmqfPEZ
/wfFXHgGZyWRjLiD+hEZrzggLNMWg80r6U+aQw3LIJIdFVm+KAcmBUChLSabxozC89pu6XPu+x6H
XlhpT5L0LVr5eErF41jDNMYgtzKM0FnR301vqQlH698cm9Hl4W4DlLfd49ZVmU00ZvY3qqeH4T6i
oQPywoZLmJECh/l9eJemd+YQmAWNZh7LL1sP3lHGGcXizXw0WauwdDa6TcakU5dzdR1XxuJwB+o6
Qaml9PNiIJgub2nHj4QXfEl+Shk835EvV259oFz7VZ9byN8ykGenfOZc9rJLLo6npnMsxN2smutw
pg8kpx9pcwjrm+0/uQ1gKVJreWLll6DIrp7tw+g6XZOswjOdDEDRZi+3tuUPVCJ4NnsdDDumwDyW
o0rWK+dyBE6bOz8GfwMpUSJReZvCgV639hnxwF/IsaBYqcGQZw71DHoW/w1jG8t4SSfb6knBfu2Q
4g62CGASBHcd68hMibh/uaSmKYGyHi6sA/WxeM/+Bkpk3LWf8ypf0y0A+1OfQ9MYTVkjvFYVbkiy
FcU3BKnLSRHrlWtX7VgYwrItpI6teP7VHOGAwrVCWoXEhJJw9/BgzgpmLYqyq/yZo874MA2toOt4
63j7+RCpuZULFRQ391lzqq3Q23ey46Ha6A8Ymf98phYYGxlMdKFItZMz7nnIst1KPMagN4WKw+7A
1ROimA5LLNpE0DCh8j7Ek2ZgROo8aJzyAm2F/4plCrEh54K4ZTIN8o/HaycPczPRyWXU8hc3ld5N
4e2i7oQ5neP+PK10bJ3DSoMwAEDnO7Jau+8VYJSZ79mqCPCZcGHGZEOfNdrZagyeeyTT09MzU2ex
A8GFVMAal9o9RqK4djgpekmF7BGvqVGCOZDjnSGSDAj+8PAAyB74l0rQbC8jEr6hadVzkIq1dYZr
aoTkv0mLyt0fvFyNK2Hcgc+E1WrWDFy7ugJ/ezGV4PKCCUwKZWLVqXWywraOLpJoOLRBX7a3aL/1
5b00IhNsPahHJ0gCnpmDcmiIbGs+CsAoueTgEoFTrD3YayaQIsr4VAkAOruOMZJoNRkC1CftVbU1
QjY6zsY/bN4yNPr+UctLWgJfTgd5cGvFUmEtxRoQZlU4DKNu9Z/GnLViA9phypL+x0EGYIwmKUQE
VjnfEjIOSnLNsX9GJeIf5PmPmg6WgaNrA9/8iOZtott9/P5zkoGZsCn3oEEfdU6FGXuZ7BUfThWX
raA8Dgv/4cw32i/cEMJHKMpS37iIyIwinRib18hs9IX0NgqwZVl6aHYWkHtvCoHrH2TrDmkHlYUo
ZsGoaI3cjCUA1ZDiuTEwFNnqYgNlKE4TloInEMnaJE/r5u/TPYpuQgpFHihidPRZggyaKPd9pSke
eY6gcb1V03uwj5OXbbZxZmeg0ieRUr1jJfB+q4/R8QMIfmNsiRXRfhoWSxWILc9YC3SyWOSz46AK
W5pd19kMHPa64vjV3z+pYzgf9oCo2Og+aXgA/r/yAwtM9VYn7iUGNwyywJajePtRRyT+/KB49dlH
kp3rb2lUzC4RNo6JogbfT0FdKWPs+vONDlFl4v9i7TxmfY/HyZLLBPNeheLBum4Q2C4e+xFbBa7i
ox7P508cSBgbHDSqiiSVEb9vmR87V3Jm+EqRGxqKFTk08NMBj8c3Ul1R7ADdlZme8HFC66TvQHga
ZMkfXYfqjHhbe2BBnXe/zrvIAq5gxZ7pt+CiPbMUzAgOzZenwUD/ISGv81zFfjQ8tbmpGMdFshT9
ejnjTCX9jLOtDtAbEhrMlYqEkf76BadTzlUJpl1SlgldED0972PBTFN2kaXviIjOsXyTqXkVE/hv
QKH/iYa7Ajk1qRd4GhTHK9Hs3s044FxqsVkpe2FMJAIZis9ToH0DL+ua3Jau+kPzwq7pdsftzyf8
aT5f8ZkDe8zys3JDM48H9ZwImLobkf4XnYvXuiPZJs2Lcc53ixm8JvkfU9esUcp4AjwsIRLscdvM
NTZTpXSLpJDBO1hEUCUr0YM3f2oBy7/0y2aCvBwHrSig1TOk9IxS5S8ynqL5Mpbx+lYPuMw139d1
EGAAkch2/T2nbx74reURn3pcQncrAjCy2uTIF2a3/V1tNxhs743bsbLE6OMpwvNCYzImjRn8qgp0
xkDFAftzFvdRos65pQUhgc4CnT4ke0NPP7F9kPY0nzk/rl7TOpN461vyG9oC5KlPyxcvBePSa9Bk
O/h6onnbJSydGnZnp4+VuV+NAteziRSNOwUq8bupeMiK+NfjU9yd2YvGYu/u0Rrz3VeOTmjwNbor
aD0DwE2mIC0S1KyIckerbiVaBkTlGA2kcYD3wSu1VPUG4z8tnYPYs4uctMZKJRwUxqwUVm0YXxgr
IUn0eoX36KQ0kM9sZbVBwT2osX6Qb7n02oF9k6Bte3HehvZm1p5iitlfk8CxIQgduTqXXzzGf2MM
HGmp0nfLD+cArkeE6Llhb644XQQ76Qcw3B/1IefyzP05PupQrOVtWOjoTOivRQqLX3ui74a2Jx+0
nT9jU3d9TymxIlJn8J3FLIuqGWOmi12PbNnMuHy7AcqG2Cs0aZzs0BtJYHffx3xrSnfz7yUapDJv
zv6U0z2ZX1X1M46EyOSqmomCNn8/47lntW9jtrnY8QXCoMe72DFILgjecHW25w7eWklDM+ssnX/V
mxtezTtqQeEiqW21gjIIXELMesMgjzJvm2pXeAaA/Zb5DeonHtr/d7AHpjor5dpOY2f7XJwwr+q9
5EtCMcoekyfcsiA9OAMgT62dHDKUpqLMOTgjS7ApRi2SwVA3EC2wa4TgWOrjOOXlxYmAzbuKk0bj
0FQ6BaiOhkk35TECTv2+Wx4VUDT5fHG2ruq+paJ0ZhPd9EYQf3bONCcwzRZd8RtpK2OqviEV+4lA
QGO2l03jIkK8qBz3ADvsTcBKWXW/xcln06pNSWhI/byH/69rWtaiok6x1G0mlW3HfBr4tbEYt1eB
8SG1zPj8S3beK1EWWl8Mo+2NvdrK9zL42JwJ9bHHHMAHU+EYo1MzQQYomAXoBsShg+pb8iZ8zWzz
b8pYWmdaAMiHCsL22Bd520mXrcFPfch8XKKWUmJQm8IEhUlPlkAHam8Z7j9mu+gwt4O4pWMpcyha
QerDOFLQ4TVXqvF6W74ywX4vpR/FXcvE/yQCtkOmq1o+xXfxcLusHvTKm4wZ2EZoS1QUbOmdZq5J
1E6sCvg+97fTTsvFIuiL00FiGLuwzi7I65JpfK02h2vFh7kjbYQlsYqFnUHlZ55WuvVdl8EGBmDh
OBQlTosJz9qhOijKEelNfe//CiPMD4iFKETSvyi4xr1hMdPzRfJ3I/Km6HLmqQ85mUtLqG1cz64K
j14BDgWIPe7GR2wlfZQDBoiLWIzDuB2puAUoff6fxn/Z86xHj767T5cPZWU9pfERksPthv179UVf
Rbgymq/wiXAL2ny/cJBVWt5J5qS6TQhKIk4AfhJunC8XLvbbpCso2KZnKARzdvbIH43CcxadD3X1
d4U61Af4229ymLjOXGUJJpmCDaYMIVC242aPf/8fClonoR9fujE4NG0I7ruZYFVnTEwtP4Fg+Fum
tmPrgIvN6lMFe3IwOqeZYqaqBEqDg38QxeP+kaH55ZxLuTzCUWwMIGyPCzAlne13Fkl3oTwmwR+v
MQDN1SLgHbb9ick4gumVXyMCNmJLw12y5oywtUJ8gDk+KKxwrebPAdvs0MjnDBgkkOE4oiLcXPaT
9IpfHxGrIrXENzwsBEwEonC+Jp6euGs8SZob1aEdGWah4WZfeE7gmdlSYdHXYm3WciSBTfIQ54pO
32uh+TdQnX2P+/ORsPSFWjejQhhAUnRy7JXbUk6znyTTjq/snKtqNfI3ytpn4muVHfbZ9gh4JSrb
0USeRyblen1TvQo2wx9TGgxzsmeO6dU7zYmjbdVcLyq5OdYe7P6dRjAIw4mqqEuLadGoT0DbwJ/Y
spe11SugYgITIdWUoMFA+PmTQbzFnKdZc7KNWRKMJXhHBsznzIt+g9oTZ84RMg8Xl2AWtxRhD+DD
+FYXgNfIQKgtvZfrV87JowOA1QLTlvUZ5erL+Hik48/3GtJTStezni7WJD921rO+oAaFif8/L3eZ
YEvO+xG5CjF35CIUvwC1VXqF4APNg2ZtMgUJ6fhTae7h1+RDhM35ZzVFMNdVgySkq/o2fGuc+/XN
/Q36PHOHwLa3csybvRdutB0uKXGX8L9wvcPbEqHeqNXhOdS4p2dAdphJCz8g9bshefkOA39XVjcc
Zc4NjF0rOClHXwJnDpAiJcfZTYCMIL8CPUqaxAxU5IRRnbXZJlxookOXiez+p9sKKMP0VCezSKT/
lxsy5NonEm+GQbnjZKEoyoC0HbaSl8sDIH9ThhGw7ryrZ4zb4UmkkgjHcctDlrigNptqSu0bxrlw
05SRyJGYZNDr2UGQaItHiROvNu+5Wtaf6g8xRLO+PXVFXf9ickAXiw4KpTmq/MXs512ArfrUTUqG
QTuoRXtDSswHtGlOrrj3nhttG0pevM7YyUDYP6FU4J9fz3BMwyko2le/bskyCPS4uU4lByznvaA1
GENQhiEfXlXylCSAO4ynvCLkOwWzJh2xbBtm24qaWtRAnKhrUiBs4VxrN0SJn4xgrBy3YjmDu7D1
SIBkRr8PJ5UDdvqzCfxfHBL64KinEtJFK5JhVK+V0hFigfVTKO0bgG0Mr/K9lGaQL+tvGEd5qSjl
V0e7B8aF++R45QzHGEc9r8Zf2aAkZZbC4YWhtS+HrkTo0mL7SUzrsOtDZiX02sbinUTaPyDUosH6
e7/wK+DGT+a8tUsQXd5X2wezk38uooY/WyFDU/EW2Z8tZRRNt2H4wqmDLG0sCRQXiYo/+RM2Atrq
tnZAL9vyqpnj+TjiqzFhUhk5tGiHet0QOaTEagmhM+9flifGTyHSs4tKtLAD3nErE72J28Xv4RaW
vxJGtdfNm21gCCfdz7/ljpvW/HMMAciYu/UtkiEnu1AX/+P7wRatyerbwSaqb5Xny1sfSGA3YZe9
OFNpc162qQzVgDPehcwTR9m9N+OpQMizWrJpBfuJMAt73pRHqlgLi18QFaPy2S+oy9KFyx94XU6k
UqtMjrDGJrac/Ob+vUNhNkQx6ppBtYdD0xZGQbWQYmcq/Uq0ItJApU6yv+Q2tHausPTecGg9ynlT
rH7bBvrw+rBZE57YRsGy2k/FXMFqo1x5qrx0kgjK30h6FuVNtWYOPNnvwRQX6CpKhBKur4W4ECH0
PKThBL59Mug+UsPyinpmu3V/v9mo+xoBMXvEXp6WmW6Eo6AAUEvOZesPC3omJ5xSqb4iTCRiCdkv
Xljhwr13581Ots0+hCSWUeaWCMpLk7v2Qih/BzJUkJVtgOovkMuLKmD93vI83j0QTpBgqZJpFONC
c2f9RPVec0KP7lgjHa0YGCqKPwAq3mv+jLWuimFKon6LEnzoTzYyeUfqRAoRQ6K4dElbdEz0F+zL
t5HHNEbp/xiwSMnzWbvsHIEh8pP9/qbLr1R73MJVeI7+AmbdKnf8qqyGExSrkdZW3bjq7Kpzb/M8
YcCZ8Vh0HvjGT/lSDgOa4yFrVeAP5A03q9+4GMeCiZ00k5tLHiy40J/5rOxXLIc7JQcNhlrj49ag
OYqh+6H8cj5TuMkNMtDFzN68oFHU1PCP8LVBSjMRj1VgMo88uYdiW3cC/kRQ7C0FQ2xkA4xWbFuY
7ioICkWGLsdIhfC5IDZ3svSphv8mRTFczMrRYV4PWrHF39zFm6mJuBKuhSNVgTgMVMvbq5xD/SPP
P4ozoks8vnrdineSYkYj9Oc982NbaEofVeAnXZdBxN03mhVjTPbYknBJY6qeNz8q/lO7xJsqqNgI
djG0GRBu5oFiI/czZ9eyeU9navCiclWzU9ab32p92uGcxgdm4BqTVQXSKm45E+govRX/O7/j99dH
ino4CwNb2ebyht6OfU7dOHfK7/kQep4b2RJVk4hBjD0LAdRAUIG/vxLtsgmZPQSt1Aa0XWHeEVnv
v0uDV4oFdIjT2kaRH9KjM2/pZkfuLigKJSqYXI6LOtVnty+z+qaGZa9r2vmExQ0gIDeVPBFgXDGI
VM3t+0t9sxs7CIEvfziVOEYjH0M73EX2ImSeYlHETPAJdDup//GYaNc8ql2BYOXpnxZaF+pJD342
kufbSwB03z88RLQxAy61RAXOfqZOV5pFs5F8gvLa8ThkbMW8DuvHw9X5oEPgiXorIEG9DTv6j+Re
LHIGAZ3EmzXQQLBLq2RWLoLoiDG/SB6fxIcaPRF2LyUTFK9t6OWH7WEfilNMkY/9F10jHYjskudl
mL4CDlwy4XfhQJESP5UCtWGJ2Dcff9KLFn83YnkJjaMeQSoJIGbi7EwmZ5OtGoMrgHO0FtZ/n9sW
RMwfpu2i413/jDPBm+pCdbWKUbNp8LRF32v3WjwAAS3zpQnkFY9Hjczckh0VlXZ/bNinLAOa614a
XtEmhpz/RTtGxd09rFiUQ7ck0R5Ncalx88z2mEVUt/rt9uHdXEhpsC/7fKprkL7xL8pAWP0iAFy5
sbtFkwcIMcTdtUKRRxda5lFsarrSn71TE8DZZQfLoO00+kizp2qbE30zM0684a8LMqQnI9ybG4Bx
gGDBFL/ye2ZxxzIo8r/+bFN5jZ+gRZOB9FLddb9s1w7u7713e07lvAZeg5njecqRN0gl3UkPCSRO
n2Y2C7BaBIjJhJGr6qjbMYtE7bf1MB4q44Hh/ASIHLdvFT5UTIdC5x7QmQ+bUGLIFCjEH4a5yoJp
iC4OwPTpyBUwUI4kT1J+Y9FK6qI2bBz8xiThIzJXsCKDUbUI5SNTPvxPDIVaATRF2EPqGkfU6vhZ
H6/WLjUMcdBRj7AAFY8jZ6ddAJSEL/sKa7QmZmLBLjwueL3XCanpYxDwBch2g1Cx3PV2a1EAyYBg
JgLOKqcr4SWwZUvFOpQCYg2kQ91kE9NYpDahfFCrUDeiQZmduyHlvUaSrMVq7Wwyki58w5vmwtyK
B69WEtOriMHkoHIUzaWVCwzf6J+IkruUWOF0xr90L0OpxUyLCrdp7xX9rYjLCe3YOHh3ky//kXPl
lbanbq2v/9ZFQYJLtH+HYyrcn6f/BR3L3bTe2PRCIeZcas16KyNKD+P6OSDYBV22/jwehvLRUL7O
PhVtnBwyzNEYDpRcfZd5MhWE87EzLSFPjdmBx1eGrUjEpbWDQx7YacIn+eTvxzgP2xhyT6nVduR7
UteT/ICR7Fqn0ZveAJm9BOqbfou1n0t7lTjkoQOTfbcCuDDhtxY01DXHnoJajEpdi1T/TFEAMdN7
OZlucp1LdjMMXGPMgzt3Rak5r7MkggebapQ4CKw6SjA33V92kFvjFV13ObP/LxyFzamAzZoajrTn
3WbzLoZAUeBW5b9v1PvpDQBFq3EN7s1v7lDJ5R2e7ekrgpew9QtqV4wzKBPwNu95RyT8b5uyyvW/
+LlwlzAS6AKAQAzSRLQJLwl4KDRTULvLx1vNNhCV34WtrJGn1C8KW5OL93RIUJMXqEvxuyIROjGE
Go2PK3mI6Oef7NfmTr80lkKW0iE8EuoY126PnHpxZdZYrIIj+eIy/l752KPdzuBfYrHqlNk5WmIx
VAt3q/JSYNo/CnoB7PUfvvJD5RsUBQA81bkYFsAcu5mBN7FKZ8QNAsllPpgxa8MHKEF0lOgLIN+5
W4mMeT26OpTSyxgH2empa9Sl6Me0/deK1YM0v8VWVzABnDHeCixcO9kjKDf+AjJxlsDXqsueSmJ6
9aFDyQ/6X3RZsn5S3e7A6ZFVY+k/AJYW1Kk7lP/eXtOYvm9qcxTk8/2XQSKn+KnEWFCVrR5OjpXc
ju62lyXxP254AJ+eKcoRA8b2CgS399m/HyRMqGhrEQd6eM0mbPdG86woW6ev6muTviLbeikjqzKt
3Ihlo9+2SjFgOiJZ+NrLrerfKB9LvAmAVLGX8dif3U58/kr6oBYMBBNKfbW7wZ4MzhK0h2NtTTwh
QIwvP0IK96jxcMpbAWZLaDBdTuxMHrTd+XgRRokMVu5iSB0savsrv1jXgd3sZnyV1tSdaVdyd75a
Jr59A3BHhrf1giB5TfM11jEWOGeTJdF4ylJB6/n2IXNAEIzJr69YUObmJuxrVS1VtIz730uyGrwf
JjZBx5BmbPypGIghY6PMm/ztgRJLbpqeMODlud5XyBpo7wxuny/RH8AIHzuYydpregf7VbvwwINp
3hjPRdjXRXR++cXBbehzrVWiciFcKEHKkMlej25AX4JJQpoyDqC/RNSOAHv7Wld2sUhxec5bgjgO
3/A5GXBaktE1ttZi+miGpn3CI8tXm3BPW+z4eqhCVOQWHmcJ5o4MO22/lJXerI0S7ccNridoOgvE
HgiXk1zBoWHWFYBnBqyvJSVFE4fQj03t0OdpYjZreoP9ozsUJ6wajXRwBi6CGPCyrfZKyx3qg5uX
wCsPyAuqUrmOjNwJjPQ7Q2xAvMIQBAqlEirA1eAtkMdKr7exmala58zxRyBMsIOWSz3g9rNrwqvv
6IzcttYD7txTv2DwSmqfOtG5HxPwVW5aQqYwaXp1lko0r148i+9H/Y3tT/we4Q29N1macgAk9Kff
U3HHCn6efsagDe+ZCrdW3hGGAM08Oe2vXwVXdZ9LanuM4Ht0uriQ9tqG3SgLkDcglhe3JhaiV4lX
XNfFATaB3tEFqBFp/4ONBNFQf5WUokDRtQFiwlb1Qzn7wZ3RfHJC2cdLyVIZYU51ZU1ocy/cqNeZ
H8TqrVn1b2uQuC3ky86IW8quHCCW5BlDKJYYQdu2XnN8Y3lQROr4q8a0atkRBTbLNpZZJlIyTfxc
d+AD1QnVVQZ94GwinwjaVEvurcP5HUVqxCprSJ3VaRAcfbWoCTrxtULCMezHPxjnqrrMMU5UljxG
da63DMLldagDPCYn5nA8RvCldwtIMkkbsZ0zkEpjJqI/Ki9JnW/Ch4//oPFls2VTFhlI1dU88YV9
kZLq1qs244ruREsL8xwHX2ayTZXlNfSMvagoyK8itFCwu6HFGzC9Zin/4sAYKKfR5F4dz4u/kzxC
D6ulBLzFMdakupJFVyakIswCLWE988EF9AUpK4NvHBfEAce+tnVy28g+Rv+zSbjM6S/V/JIGhBVi
vndiXRtAK6VezeDfa383f7kGyhgGq4hOGmLPTcgC1TOE0tX3OAopEDTwnPbLGRv8J9wmSrhX1z7K
WMU2JP9MIYuY6SowB98lp+pbtQFUgpYmP1Zf9rvigc514uemSPGmQBisV30yw30D3VV6/5V3ZtAP
5TqHH5zze7TI/hdeOnXsSHKs5DT4pk4TjDCCLcVH5zKBYbhnEywpGWjszEBeKmMBuYKJGzSjRigv
EfE4h5h7vkCKnDfw+eWZ0TLICfRwl9jMGvqKlXSv+RyGkfaAKZP4CvfhtJWPrLYFCfigex9F5b5y
2twbYNCwde5IOS6LiHmFylowSZ9HTejVsmYXKFtfcmAQ7qT+38Diw7jH/423FMLMNHx7Q2v3GQaH
jDU4i7OPhshGhOdFrvI7uw0o4nmFuxbG3+U3ojq6Bqej1/nqFnNnBL+nhThf8LkctveM9tnWg/73
+fzHm0I5qC4lNLtuPvUbGvcRDheBWbFGwoPGjgmBYqItv/oPhhaB2b8WCSzYpeVBOi/ARFS8jsr+
FSriaWX3rYVerzp3iPo//3wo0XIm6WTSSCaVfNPw3GnS29RZx1On9I6mMz6R1b5+aVA1SCi3Omnc
ApitF50oimqti2kj3C3rjzlo1NTGquo5grS1avUB+yn7PNoEbvbD3AA8d/CNaMpEey2P3UnH/GXe
z7SSVpf+x2YMYL30dhaHQ5YVqA4Z6v8b1L4cV9s3EhKFxNCGcS/mEI55efR54djmxM8WI6OxURas
0LS0w1fk2/oYR4Iw0MAT/JqEuR6irj+0ZiRP106HJLq5WryJXfGILev8o72cv0Wa35dsNzitrIq+
YyFQ8j50+SiA2CDr3I3g9hGfry9RBI343ZYzezxQ1CEjU/ozPPOUgMNnkALKeUaWOB0xPx5s/KJm
3aqoFR9nFsiL/yQfZwjaUd/fkq9jrjJ/UPhZmKypgSOZ3CE3rx8kSTVn5n2tlvyfOKw0yhgBd1bh
TQ7mrWY+RZbrai/tCj+5HOqYCwGLH6np/OCIomnf3Wq2muMMQZDTTRoCJiRU6wRz2xrdHPiTyJOl
oSQgYlRtVX7+3vl4E3BpcV/uk/jixPlI6btTjodYRVW0PEkD306WTxe9OnWFV5o3sAXvimKPZYrG
SLqw2khPVzpqEjrR8B/i9+VQpPzQSXsht7BbWsaMVqAOIqT1kNYbUHedK+tbgjBfzVlpBfMRZLeL
flYN+VvLlAz4soQU9k3QUJWLLHN9bJaycLduAKAFiXFqj2oTlClbYr9Jh7aja1h+7vQo42cScbpe
lJsYueZuCK/SAyBmhmNSlzHeMNtOUd7m/mrhOG65XYVV7wo5XtCqOXFjswDxMPKEqJriHxtWUv3z
3qIDAYS/f0wi0CQbomJZPCaDHxP2aUbdDrZw4UZ6hyZxxnnQSjS6TTYQem8p+gSACsp5I5RLX0dX
46YdR3XUbAKpXspbQMXmKmeV/VSaEUjckRDvXiDyz9m36ZIO5p1KDAi/8XDuam46hvHK7eXGKNpq
/p0i+YeotNW0oHiGFNUmk2ujeARnyeoKr+WsEsUuj6M0zQz1qhflLSs4GQuWO13dX2e2uCDUUzf0
N5wsoWcbOUHmW8/FI15cZMNe77jLMIkm6xN1RajJltNVQh2mJNqkh5PeOL7TiWd/mHtnSEGshnj9
ApI7kwN3QUR9jfEzTZqUztnOGMfGX+rMrx6fRMPfIP0VzUSl/hadj1r9DYZZ/CQzr+WAHiiT+61d
3txqAraLnZ3M0OyF3r82tPnkvic5vY7hJ6iy6H9gCwOokzmZGAFvQQ6chP8uY6bOgur8XmzDoDO9
RHT3P1psT7ZGYW09dcY6Km5HVdYPmlBscSk6kO07rVtvql13uvEqBJT+MN/kHwoJYN1s7ZH3wSrP
beYqP9UsfJkA88JcoqFK7ZfDKux5MmlpydvZj+C9wZ8D30+n0jWU2LODraYVgPmei99e2hvXIZRz
sgJ4UlvR3nAl8MAY11UzJx09xR18e6IsCt8ibmdhEHjjAMFCqf97ktgHfi6B8lFakQjXsYqfxcz7
9cCQ/hc3LqjrnPBn4ah/wGetz4kbMSBJV44OVOph0AyXXtzBryt3xebE8U6GwOSOC2V4GYGS0/mf
M3mI6yrUEZmriAVxpPoSFyLNlPX7w3ml0vFf/hwTeaTucNkq07yVXUqECsq7/EsvRQwHteb8euLW
FbWf7E5vxYY3Iuq2+0vL2YhqxPp/TFb1NcGqNQd/9VCUinvbhSRKwvgFbvU3foGEC7YmuRecc1H5
GXvmRDVLCpYu8Job+aQILdolsfBwI+Fc+46he7ENpK8StOrmKUvVPshZ53giusgJ655WeNSY0qqz
3WdH9Oi8+CmCGdxkTGYm6cUf29dshsVn7N8LYbV1TrVj0DlHXWdchwaSwh0M43uR9csZqz4AL9GQ
UYimyLPcnLKhpR5GHAI9TcSGYROATHvXgS3As4QkVAVgxRRlDqDkZSvspUXDhAMj3kS4i/OcDm/r
zBBMfC9wFlxASB4YA0010xg+/cPltWDgU5oXECSG3sm/95mBbRVi0U9BwyPK3kOWl+BGltoRd6pn
wdmwMNCpkIm+9Ig+OQJ3cri1afgOoXkgV1SLoxEeUgxzJPgrBlRwleVLa98QcbJBlqpbpd5dancs
9CO5uNtnWI13JRZ1D2NRcjIjzhL7N4k15H/COpLjHMAMvhYF2Xi37scNvhv/SdzVQ/S3iobTA9V2
6Iysn7Z2JiCzWy7ApWNYtansEDwfBZ0VE5Zjez8ocnf9dfXCK6nQACATGZAsLR2nje+U6Z/Enadn
AIwniUN22trEmrpfvMZme1PXn0tJQSAb8tVGBfK90ytMNyc3kd7GuyTf5BykPvRp34IZXaJweqLv
wdix/RG1KXb4R8XUFsHgHkpvp7j0Pcy/JB5UHu1JkvpfYpm/KYhTK7N89GFsFGpZK80BafhxE7JU
k5ppjb1UXYthNJ75Y0BOpzGzWrBxujttmvGNBX+/qNu7uLbQUrpFP1n86Pw91uPCFwSlZTWx5T0K
1DVuXAL7fnTa47lY3ISzGwLRHq4iXtRsC0X7TXtid75AO4psp0ioup5lMMFFncSBo+jAj4ujs2BM
3wS5B3y4NZc+AyZr3YqzpoASXt+OpFvJ4B8//g5q6t2w4GWx54uGHQuaggenVCfPtb2SecDaczEz
UVR36+Ep1HFQcpgkcpNU6/0QBaqMngXVY91mOdGdvCfr/ZEE8N+Jp96Ae+kj1sx6bLfjEc+J3r44
xVdsJkzFFdnptHCBaZKtG7IG0J8a7y+ylK8L+kJZ9rKT/kuVThYvnZoviMen5csevHg0xBcGFIk9
tf2I29IrQewUclAISPFUKsptKaRHePSdPQSRGf7Dlp3x7aYh3/Wxhku9YlYWHbVtgawrqT0cqxcB
AALG9A9S5vFSz5DarpFkscWQUlJMo7MFO/swym0U0prIfB59xHcKz1oagpNYZO5nqiZqC8XGZYzF
OhBlV8tTn3VzpA3/FVdQWK8X/D8otZFe3M1QBc2t/JVbS2kEGyOYZR328/UKSIDb7baARW7Khk+0
A5YMIIdyHr1hhQzHTScPxt0iNni/JAsraM6UjHhBtUlGPMkoSLvJKBsvPnHfdpe5rJeO/O2RnCCN
gQ0PUd81H7+tG6/JqWTWOb3ajuU1+8c4oYKUzGow6SPfXGDyJIjNl1xTG77xchqgnmLAXoqkn8F8
QRu2ItiH2OqgtEZPsXZ1VJhAWWvrvFC5mFjcLNdtqkvZPWfLnTiMjGzobAmmk8HtUn3I2rrrTDV3
CT64+ygvPBjv07nsG7ouBuyO6OQpHVXODgm5Hy2+3Fi3dhpOgpXrsxsN/y3qrjhJVOWp2/c8JeNV
0kZnRRMO1Hq+6E4gdaOkCV8EjMOitBGioqVGpP+It+B3hVhy53R4e/TQ/fOpCpRnmDGevoB1jNKr
imE11A2AENJ/Q1FGdsotZtECWUK0VMfcwIVAM/J+RXtCiNOnynP1VlhN7cmC90DeP1tIC5JSDJc1
TCyoIpdpyABR/1MxzgWdtcEZQtCa+tMN0v2SrYGbCIzpYLKNAhHOrqn0qO0826V9J8LGUK0tf18X
61Tg9LBR9NYJQnXc6riB8j0DqrqYE9O2vIH4T7PIj7P44rSVwMWoQk/4OI+wU7N91vmMOi1dYxoF
6TWvgaOGa74dJy/gpOvFB/dmyXoOp8nEbGeIZ/5f//KmFsk9KpXDXrM8hCScCBjimbSbPmqKNEg1
2iM9MI+iuX18kdXVBLxm/exQ50Hkx99KWAWr6/Bsy21YevVLxWzvYlGT2SZfbcflkcOUYhU5ZvE4
gFnWDQ+pHnhfBOsE2vf3/9eVAFf/IVZcPhUndJWsiKCA2LypA6EHvvYMQDljzbPGavXSTpwki9WH
ntlW4MTG2k4ATxGEWaOpwnmrLVVfudPJEG/WoB/vXtRvxBaddx+O2vN2vOAoFduRyfd02fKeXTex
7E2YhqPawbj3gWVIacjO48NMeHeto63BMUMxMk7Ex/JJux9+8G6Zv9wIZITj/gB2PNZwjEOeagkf
5t1UasrYc82N6E0bktmnEBZJCOS4v0iOAOfjlvoqV2J1x0TvfUIhxthkn8i+0G858QkCNmmX0Z8w
r7Mt4thVLstVrjfYCSs1Jl41B/MVerVSbeQ22NhJOOpyQN+TQDmP1kSAXYrDBczWzG+oIyVRc9Sz
8QOsNRLZ2dhQPn1wn8mcFnYZwD3mFqPbuTvLyLfa7ziqik2BxJtHVZshCS+JB0pEdF2/nhuqTnJc
9BG7RkWlKxU96oT38Jqq/9wyWYZO3FGZ2F6SBjQErSA2NJ/ARl0+W4XUBWWHD3uryT/9xYKlSAcd
EnfbAXSs6zHlsgQWjISOpX8sZtVpczv1IT0v5emhXvblu2LF8msIbiXtH2vMGgARsYV5WJDtLdS3
iXZiJcG1jO/3xwyzPnfoEkyOUdKF6Sw53VpBSkXa5YI+MMv/WTjdzKUpYaVHsMKvlI+yXMbUTv6h
UmZQXmVnLeT2SISh+qiQJh8rxpmEC1VSFYj1hjjWc2tAmWFaVA/yNsXTo82J5FiLXzHJVDrCTKDO
2f+3Esh8sSSVCaWbOb/qqZhafnAlcoNDVVHu+R9RHxuPNsWhP4Hg6KBg+ykMthfIRCI8FNTdIdDt
k9m4SBPaAt7LL5rm4uqxqORONBQGBzOOy0f3ABix6PtQxh99yHB0aiPSqkJF5lqGcyrhZi0rcDeN
XCu9J4TIy0TLSAOWnBI0lU4EGotegOJwVJio100zY4GFOpNCDc7uyU4cx/uIk6QuSvWYQM2YN7EZ
yLrLZk3Kkq27OwtV1ThyiuCYAfcBBB0fpb+HpcLqa5Tx0zEFwVBhUp1Q6vhAxFP1sOO+7lrUIlDW
DxW1YoKcggiHW1apCcTVGaCY1CqsLTv3QCqVXX0ZGVZPzWpgr9zJbudNbJelA0rvEBV5GPHDnfA8
cxGu9u2g+A4V7YuwtyDIowQNxkOmzM2RpU/uLItN4OZzFoScb6u0YcEee7c6CP5a2CR7+SL95K8H
AuZQg84m7jRlfatOCSGBbmz2euPk/FKSMQMkp+woj0Q0K0uWTJeS2vMSiHo24tT4w1ttcVS/PtE7
6kQ5toTBjFHosqBm0LbZs0MEsTmfjNS9U7tAKafMbLuo82YzAHBOGQw9TSAFCeQkOKamELHpI5Zz
lUPkHD4hVYqC35l9jZ/puL2Aoqe9V4LsGEiywx2dcPJ/Mgc+Pkj1+ZBmS6R/29ZIWTJv0BdoInE7
OAEnYr/y7/gPFZ38YH1psWfvj4sAyb861XZR9DkBUIOIKfl4dBq/7M0GbZbsukhoxTqdP6vPilUt
eRjZBpBhDwGLK+6OSkRk9jIxk5rUZB3cYjPuw+eEepfxQi/0ZfkSOupkf27+w04uMlnROSTPgSDb
OkXcPSruGoAUsQnJYI4c3/yVhYIjHGXbuIQuCZ3l4nFwgXXxwJ6OZ1HqkLMYKJf3R8rTtNnP9Kph
ZC/kq9FLp2gCahUFlyLGFWQ1tQuoxM85sKp8pg3pp6s+mL+8sOTTxw75sJ4bgWrSamL0xgbr/EXl
Eihfzv8vRyWub+/s+KpWI1i/OIklZPJYXlnTpN0qi0+zloayIDkoZ5uCYKpQAotmxW/AKjJUj3n0
cydP7BflcvLfxiidB3/fOq2xnOLA2A1XqugAF5RIyPGRGGDeAZ5ovLmnS5n+9upclk2j7Zqtbf8D
/QREosGxLJcbzVXvxyAEQY3oLeIv02TKa8SQywVWoPTPcFnDKV1NMMGH1CcnY6oXqgzMvZqNvUte
zpyb8tFSyawgzMF8wJJTWlA0mQOVH8IfLyTZ5NlyG4ooeM3fIU49xjlQsqu9l3Se5s2lwVeqxUD/
xoQST5HOxMaFyxPLCebrn1nzRUxUTz7NwZV4pY3N3D/5x7X6M2CNNElhNU3QWSS635e3WDCHGgSi
pCng9bT1EwWzlCGPaLIJulmLl6rDLQjKYSdpHBHgO0JPByoUGLGbUc5+WCzeeZkTxwDVjDx4VLe0
Glq4vizReX6aQE13D6y36U4kceljlxaSvwGRErJqtu7PL7CYM1iz3qbLhEcq/F7zLmokXxtwXoxF
Q8m3scNFOVlQvX23SCBwye6kn2MBOWdxMpZ5Br//lv67xMYmYujlgkw7RwjWQDSJfT65mTifSC3V
ErNIBXtFRPPEZEvu73QmDDqfQrPpCafJAremsftTx1sKaMXS+T2Gcn++JYp73QoJ1urbmawPUOAS
RSMprSGxcbjUpT3EDUvqw+mVJ8RMz6oSvaetj+J1XIYt5pyoA72dPwDSgniOqzwYGcNy/7x7r9UR
rtAQbeelLUJhMHQHpZCZK61ryVge5CiD/UfzJu2kYh/yrD5MN3oIefClj2fzUs1gRrL0MzSv7Stk
3mtj4orMjpENqkaGyNTZZ8hvCy61v9nSwsCnH9UUjkV7S3qMkVesg89cxPEtyE0rDsPyJttUa+qp
0W3/JsaAOaTJLNRpOq1jEseX7UXIRJai6HzmCSjQPYv+a275t+iUr7TNFxI5k9FfhY9c0Ih4n+v+
QAeeheS4sDoOIxhsTycLtqeSn2BRBGQ7OuFJ+EP718bi3J8L/M4hkPNw7YRzvRQ9KKwndYQeH0gv
L5Hd7epdPo+G6N2FmTmvn/NB/kK8S1ls1tGHZ01fFQ4HiBLlbEaMtRDUP9iLf4RMMnIC4s7R8n1f
GNZP3BtVYBTGTrzn+EQmZH2qqFpe48r9/wT5oBg9NEjiPYyYiLyat0zfvYge0aN2Nvurw5UYVgVB
y3antOX7lnB4JJeXV8/XqbiKjGOvD6H58+SMt3RwrIskk5GkLkoj/gD15gArnTFKhYBP7YOA5QKr
B19OlXiYbLGkcb21ge0PavVM5g+XJbaFnGackvSNFAaxaYnwi33CtqxDyib72/zGqoFYdkXe2zMM
wiFKCLvfCDnyX+cS0S3CioQuh9FSc6vl2dFpIF+DWU3SMabW1YhniW2T7QttcanP8FcpSJUy6eM+
0uo+xeo+u7zG3UEsaQEOeOJftCmhUUeTDk/inZHYpt2s7Wsoj36pRuyZguDstsuwBEtUURvYmU7+
5xhYuyhblD72c6wOPTiqNgr0JzIZXqNrBPMfm+BdW8mZVTbo0yLbGH09/lHxRQMk0vOnx6gw6qeo
4Hd8yABa+R+8wXTxqGa6XWU7UlH4SCCuHXbamvAnbPFeIGUAJNTBdyhj0BAg30gAj7tp8CJwY4n3
CpgFRd/fXkOrzK4eUM2LHGPZHLl2swetQAYjtCJsCvYVhrx3ScWYgOIwt3cUfZPD4ZfTa7PfnfsE
2WeA0OR7LR1Ut/P+FwssZnXXKHb5yjMIGKIvngXkReXcq+u9TET/tjdjr2hnL6ySYTk1HB/O+Mr7
27/a0Ziogtu7SomTsXL8JbpRwMJaYpgBlrpXoDuiOR+ujpERUvejKyNVxM+GXG6f0999BFN3aL6g
F4JpWK1cttwne6sTsF5ckJtSGgoBOr1LJEFiHpXGFx8qeoLyaDz8IFH7P/5RZ617uhkRzYusnQlP
4Fjma+G5D7rtT0oGnl9L/P+HxUlc1FDxac/VJSjl8ruFgdEtiqjSCTN6DUXeWdPZ3v21qsLNZiKV
1gVU/5rCWi9WXGxBctWTtsLVB/iHByHahGKTkKBp9cq1l1g34E1XENgHoiHmiVDrMnqg3DaRPDo9
QpXn/7gb76+uq+2GzbIRSC+BN6AylsBHB4VkIio6vK/tC7AykVX7pxF3bfaVKFXq3o2A1YU=
`protect end_protected

