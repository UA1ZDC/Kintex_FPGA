

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Kv0N+ODrJQAnD45jVEsSEPytnysm3pvAbJ05V2JaqTdEQNJrijqrY29nJXOyqQOIioMFCyAehxdh
SS8dEy2RvQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
wl26nrMFXa6fm7UAkMFkRbwMiWczBO907OqYX8JeRapSfb54ShwQXeaNsbVvqp4GNYQWgD8fiWsc
Rg1ZH/ALNgmzzsXH1hqu9qf40O6LpbgjO9M5gvRZkEo/Tsa2oqZnRuXHxvGdfSUWwgm16QfnXWFD
HONMKYo+TnX1BbyoHuA=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
cF9G3LQheZJrMO7arGfYkxyoON6brspPywtxFKpTvNhoNGqsA1QaxZgfesvqKSR6jIrBuWrdpeSm
PoQl517JxEpEF310dys+9f254GuonHdyipWsWNgWjbTCuw6rYLvLG1y7lYwgHlSqKUNrBaGYERTL
bx0Arf8JZijWzxoSQ9FVJxjXj/PfvGzrh6e0n/oHLpafMxMPZcDI+yx5HuAhNXSr705mAXB8bgRf
GS+N50n6SUyWqcyUqw3kHjqQ2U4vJW+j5ZC3mQaQb3xJkZgzHfCaBKMstoXIjqY6XkB5Su6aeqKF
tsdYwq2h1uyBfljsOFo3IsRsUpNIiryBaM1j5w==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
fN4hvSzwAQXVTyvBcSPI9qSFGq1b0QWYvne9odu5QkpUwhn44DFKeJSRI90o/blLQLnT5fdJ1IVC
mwqzRlL7DmT25nQgDxB1mM1knf9aPQaDbovHFOWTzAPBPJqGcsU8B7iu5g++kkRlIJA/0D9NUZP/
zdeXDuR/f3RpGDQ9X3WIBcSwde7JdAaZPxu8gycDj+eAg//eJ+Ch+IApwl6KjZF7Lov59CHOoVNR
udrlY4+R4MFUEO48SwDCDlqVGTYZykUVxSqzXifsrNKc0qKvKF4GbqbVHDidoVCoh7f7Jnj0snvM
x3DFGPDnokqNpDBX7xF9L6+GYPELuxQwMV3Yog==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
MECPOWJAU4w/UvBGQeSeElgdlWQuUK1on5QTAzUF7zMKC1Dzhpw/yWAmwgERdTOHF4jFwSXDGCYX
dcq7yoSgrYHNe1Z9FD7/4uOTgF7lUDYslV5k/HR/cVW9QWbwl5jLUaoa4U/BsWl+xPk3gCXBhT1o
1qrFxMGkr18FyvER+gYFNuGtJOdwhkp3EWSeT0uUZpww9gD8GQxRUyHQJxyLO7OrJ+p6c8iZL8us
t83ykRj64BZ4A7H8a4gi13wX2JOPHaLBMG6QaY9NxFK4P+cAlJ5tz1UR5CiOSua4Nbo8RZAnEv5U
qSe9Ctk2cb+fZHyT1Jbe89K38c/68dSDrW+q0Q==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JGQumRp5idVwKA3zzoqht/27epSOGyhvfg4tXP+tPHgo6OfP/FU3H6/X1Nd4Y66ilN9i+iugj0ng
ehLY04ISDe8fLdY/NaZ+qOkmAGDYirT/RxSo79rIeXhylLKnHv9FphaO49Z/wGAPNVJcMj7acDAt
BmSxt3Wb7gOV2zsovZM=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FGXHNsFzSGXjbxp7bvoF47vhF8reHgBm6BrifhO2QcSTwMmIfvC72GA44UQ8v8jHIWHgPlay/nGH
qq6loQoHzagZ/voRdMzWla+HchA2la644cxBm8f8Fq9WGjAfrRKdp+ka7tSEmDbdQiKs1i43XT8z
Q9z55GPf5g5GdS4wXPj3ZM9TkEPcyM6MWas1txHsPj+r/l+N/OJNLRx9g9A23yQcrqoY/ibZoyFW
/7no0S9W9Nh+BPh8OXy4CwqtsvPd0/Zl0/JDLnm5d0hcEAn+3TkTvrZq0NgpjAEEOfrxtp+HqvpD
SE2gPjJVpUBZWou1zkZKYyakXZCQodq+NDtzNw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20128)
`protect data_block
ymS68joGCzx6AWqkg8Oa3rCpSU1ysot32EhADcaHVZdvhqgznxguPtsXjCpyeNX1C9nOg0vheE0m
Lso/0aP26opEFAeYMoDxNfPwQrUc4ReHNUqp0Oqk78ppxfd4OYCXxF0oDJz4BPo5PTm/YZG8dq7w
q3FupWoy4raj+uM7ZPk1SwBGE4J/gYyuPB7HPXFeTQVaRKufhS0ieqasyeCmdWMcyzCmvk9EKOCz
iUQPOlV/bLXsc8xhVJGkVKGiwbADD2gaIJsp1Oy6t8o9+Zws/N8CVWpESwx96498j7aF3BPpVjJd
gql8XzLcSYK565gGWshp0vG/1pbPur8HAyX/jAByhveZuP0vQJlXpozSWu1LuzS6iQM26YjIAZ3b
eNCZRShJBaRdZmGfIAEEv5zlzFsYT0C0iRvHdgH3vaSb4a/Muiredo0y79akJPh694ORoPc3MXyM
NvKTa0dBO5AipyMPZiX/njVNvdDW7oW1ApmsYGp2fJ0Rs86GJun7rltumgf9ZtfXQDumrVzDpd6K
4mn7kfOG6LY6kOCzMXJp/sWf472GdATiDtMGyGzamTQfihB5+3/oiK88EoSiWxzQwBA2BxR5QGFG
0mNnsfeC/vW+co7PsLPMo0MBpQ6FIKS1n7JyiWDZPZXJecBr5rWGU+F7NPlUkVJ0PwP+gjHFIiFG
LrPhCANOgm6MMxbj7aG1jsq3NOrXJ1sd73lu3xi4XVNnNQsXSu3cGv/MIN4QYbIq60mtd3RaryQ2
RurOjYNE54UiurPAw2aFHhMb5o8L8OAG3B9e0mosJuoPI/zTgl1Y/UKXSPpb493fdANKUQG2bXpg
vesorya7rKM/mmDTNQN6PFZm1upM68+JQER45xC/eN137O601tHitbcGTF7l4GgjOkxw+tE2/qCn
QUfhm4FLRGCzRleYvpe34VhudRth5fn1+s09x7axJDN8M4R4DgONIF33KPUrUZ6Xm66Wwk8F11ud
RXd/A1jyK1Q5jNN17e+qJnB5W8x0AYFsWLrWtL/R9oeFD/3RMAJEi5XixWs6265VzGwv3EWS+B1z
Ysn9A+A++Eqq0C333DVdksSpQBqyHjKytLnRcAHwvSimg8G0rQDY13DHwdLctzQEqYj2MYkympXA
9/+JYqTe17NmubYVIij5SR6zHOBohHSkkN3jgZH39HWeQTbfUHOzqhf8NRH5U52qb9MznbZ+1h/I
x59f5aQ6I/pUaQpqLihwXHHrv1jNkLzzKDottXxALJo+CjykM55NHU3YNoz/e1pzSpaDyI7zaqmJ
zltcBU0oN4wr/YuP0mBNGtwhbDp2wt1ZB48obi3LLzsfhMsGmM/u/T42ArMQnhSnCwNH1Fe3t+wO
YHLbTGjeNq4ijmC+jwmrjDLOiGnzRFmBVYatSwUxDBgCveou/iJlbc8jpkW4KG1MfnOdSC7tnz/h
xwnAFHX0QpOE2bpTCrQevF6J8Q0siZXB0w+yERszrc9OMg+0V65KItKkBouyEiBz98GXoWdo/mHu
lTjO9DmDhme5AvdlXOi6ikkV+l8pyvjAhPBKZ8iC78ROpHTtv6V4BdvJANeyBvSVw2KsBFQzd6mb
RiGZ2ohaTG4jcdABRZ5dmZUU6q3S016j4PaNrj29s/WEf0gzo696KR8ZGFhQNHValy4WNkEbpk7N
RoEBVvdx7sTQioB68HGLM7QEBMzKVTvdvPRLX7EZ4NG+zTw2EKseJVRWYugW8tsHApAa8o5F9VPI
QRO9INfxZ/ooTW8pT6PyRP0H+hOKuR/eG1+HTXFAd/j+vTmQOVp1wdI6orsuILut15P43tfP/tAN
U/G7Y3jKkyyZBF/s2XDcL+FvGFdpgeIFGp2dQUWy211awBheDpC5vrEJ41DSs4YyIvez3EhgtJGX
JeG3asgGGBVL5dIP4iI3VCJ8Enc945gAN6le+aUJ0RjfaGqkXeH+6DUpyVE4U5MouZ2kACZyojSJ
/i/TGp2Ha02Ft2cR1oYmePzIMEEY3QKU0azgn72JBoqoVW+cxjPwBJfS4bBLUoJ8dsIJ1cZI+3GJ
C7YqseHElX3p7weRS8o3iusEqMEnRvgD6O8W4BB81BaBHkOwLAXwgLALlbZiv9wMOz0RnhX+f6Wr
ZutJ/Cak5b0+NK72UjhJfpWcq6Joh9O6N/rHcq+rB4qoLWQ0RWiBF2lAIw3j6QrzHYLRzkc6dEN7
dYRXgEhHfwXeXwQUBjH1fheVGngnvtsGZcBshljPfvpBnwWQoJ60R3pttijUoVXIjeJZBxctsH5t
q8mILtL8Q+MF7OF7TX1qdQ7y/1VVjpuvLjiEV8NeL1hEZjrbiuqx6CnONdePbqeEcveSR0tCoO/B
C1bU6LqSKeh94JgbjPueFGoInaytu4erdSFHcAvc2pLqpcINSrK5GdI2xohZ+Nkk5/WSzYgpCYTW
+7kbryK8DA6wiAScbrdf3tzD4nJJ9DpFq3SHVILdh16CfJ511U9TBz9D+fZgn5Xv+8C2hft/AZGJ
LOlSj1dcPuFPaMzt2QoQA10785AaUcDZMNe7m9wiM4pBb3KZKa2XjYXCiXzHsfIifefEGQNDNNQX
LWkEvNLlWnklKlJhf3ntBzyuh/rsDiGFeauSjPRs634tqPt99rMpsx1ITTeWpFv9pqfDEwd7Ytk6
NgY3Cs44nnex/oXjZniZx+3uTU6p2KWnkK8dBMArqP9JgmWWAkhqosNgWpB1Ccipq5GbpqSqBJZk
CTSkVnVRDgPDvGSNNE6DuNVWwsaJvxt400Q1p8QQwW28FlA/4qjPZCZYboq/4IpZmURfXy2vPPNP
W1Jz4lmumtmFknlE6BGhH64yKtFI7ss3ozhBwOZOhtcDnxz2bNRgLR5kxuIQAGdNoRl2sTWIui3G
BH0Vat0a8G5GWTVcKtV37OY8se+6zeSxdW2k8IQwZ3lWwHRjLMd+P1tbllj8Vy5qiInNTfZuIbIH
QoG3ligYVhTObk4Ox1p9GvKDqLPSMpBXAqsZRwzFkz4RVn5bLIBMGIbCjU6jC76GQkKXzJNVmqyi
h+IMrJYtze3DXy4hKklIrCc2WryL1VsuZHkQbwY1pPSoCUSK6l3sSgaZfGiYwY/f2rMuI51og41B
9Q9HT8wrMyfaS3wvglnmXRjJ7IRjiLxXhdehfvsBwHPMTEDK735tJw900yWJaAuKT1kgAE7ceaiY
MUQr8pvIn3r4bQgO1WjDxDEEThF3B23Q69SVXKmDqap29JE+KGrp4rLa1PX/ZbH6nm2U6i6gqfUU
mHmAbu+O2IrC9CbO9L/thSSD0+bR7F7+RzrFFQFO2ZMpoNMiSWfwjY0cp0lTeuECdM1p/NeiYnNY
wtwivmKD/jcafu8Mqrja+iiNPEP27W+XfAg/eSyl2B9sA48f4y+UUugeeorPDa2K5JwnZ9I6zOlh
1HM28pdJ4X2ukNCI9JDBGOEA9tLyT1YUODRiPP40F/ntfjs/2wRBw9D29inFVOTGMcHktPdqg8vW
Clm15Hc4g+J11iGsLVC885VpxCVjlnHt8RkvtTtlZbpUrbyjxBwvYYNrrSg60Vk2zEKTF5ceWZca
3TXFKszhV84c3mhSjE5AiolKSM+PU2pk5F3cBH4LMdmxs/kGKz/7hSm+902gzXk69HOvkaiEoZhM
ug95R9ghxgpI5ZQNLMjhyLPRlP1BbKSoWb3h45CSSeiEOiF4Q94vJA8GOxiNW0VWLE8T6qwpSxAP
q3d8NlWgT2DnA1QJOqFErlVY02GjhP9+1CBafw87QAepNL7nC0sqJDJq+cVJl91oERS0VoCE+vHQ
phYlrFeB/1zq3anNnjO2p30JMKR9rqQN8Yp0RnkUEGnjCgm8DZG2IV5p8mUZXCv/DsSK/kil22mH
VOeiX5j+Lvu1qpJVGqt3o5u7OTimqXqjR/9E7VFCtGH+5pNPrKuDLhCM78KS1ys7fdny36fhiish
NYvkmwXb0QtL9DVu5xTb1r6wtS587ji5g2286ByM1w0pFvnekyApCNlg5MemKm2NMI/4vALCU1im
i3yIrye8TU5uMY9cJBRz6xaHLYPBHH9I7AISH/LxU7MEHMUlRpxoBMAVs4rN4SUAjzNpCVlb4FUv
cDSOa0U+5R4YpUVS9wbMtkalB6zA6W8RCVRa4dUfqoiqkqAdKcKpf4YFqBi0cnKG3tfsTNFDt/x+
PQXxnJ5kRPbrtGfG0CAy/nlCTbdWAzH1ini088qYbk/VEn+2J44ulS2rb3X0Ha5BOkH23GHVx/T5
/vfJIIdJeKmiLi9cD0cH19eQif3wkt/fq7qSb0H2pSqeF1a7RzWUsjrjsnng81lhFqGijox4qSOm
mSvSVFWgSquFy7I41mVkO5fJ6NRs/tLtp5iCzvyRxFibHzXZ6JKkNQmV/QnxHJdyhS2DDT4DzPJP
WLy/Y+x91ZkoZXW+7VZsqzoJkmJsr18lVYJCzUnzjrRoMRNoC2AaX1N0OyXCTpmOHuxboB1jzbI1
trbD0x7d1675Pr0W37st/CygBsLOc1m1+9V0CkKu/C/7ikvRpCqRklzxUtJDeDJmQ2Ok5Vrj4J4c
4+xsSOh/TZChcDxS9ruevj3C2Na7497OzafHb+xsA0qHWZt+q2cMqwDudPJUSQPgUO9yR3dGNW+8
cv8oD2d/h5VugjGjSiNO9lyWP3eJVtYDx0zia7SbJGHs0hCa9+0G4DhNB2/S+YBT/nQKpGsuMDSg
lB072xfYjf+5URNyC9WIhx7fJD4pDIBixLPgzkFT/DOXDLWDLhkXvu3DDGut8zUoFQZBRzoXztk4
+0OvsyJ2ivSK9Nsaw3/4aOlDKeBxYUG6rgyNXUqJ7c/wZrm3oB9xoaJw4E6DtddAYWy+Wg6Nbjk3
htA6GQdEW5TkYHVLZfJNHJlRKh3RVMufEVItklRaZWNpatsZBOxiF3fJmXTwLAoOVB1+Dqc0U7BY
3ZwSgO6GUBo8PNwi+pBvn5Ky7lBO6dPHZB92kqA1Fw47ySV3zlwh8lB8rvmQgLy9Bx5NfUdfj1bh
bedyqF8LolO3yBasBHhcg85m+Ft7Lckyu3BtBW02Z1Q7dzQJlluc1f0JumCgVDSGWJ+nni3rfyrN
3pq2DBnTiJihJAlz/LcxftpBRJK2E+oQhNFF7iHW1nlmMp1EAq6BU1e2GM92c7q4L3EbLZz4imcf
EVO2EDUMMBoADPIII20yFxo7CvpLbnXesPdYH03Am9EOSpCSx89RQVlK5UgETVw8tpo0QzBoGJpK
vlgmp53iO0UFYWhvidZ60QCPgWD/BrJ5VGgNCMfcqRf1LsR2DJOgXSsdgf/rwT+qaH02n4QCfaSH
QYJwfvaSWT9/cO+PvYLrTvrrSlegEyR8ei0oLk85TIWuRqgZv3VWtrcjtzjJ2VgDj8cbzcoZJCh/
FZjOa7hfJF39UDDfzTtAiMWZvHRGTNhGboGXWeBQXlJ4vIKgNv0FIOVorOWTu+M9YN+x1YWbOp+X
tUU5XjA2mcut1RYF8x3w0ZV5wfGCPSpGgiO2ZSPiwc2Rv2wPLiephztxLDbThl7pxOtpP6c/dKwj
OH4vwgWenMMPmqK61VNFmtadLJcFSP+oQ7dUULEcbvnGvBNqvBIPFspx4UmBrYzZ2t214gka+jsZ
xMRKXuurOej/47f+HvPkgzbDx2ugQxqMZKEQDXGHZ/Uyu/8ZhDJaIxrtBDzuxEAWivH/F/LyYLdx
fb4ZyQocvBSSBNFYAKLK8sJx07db3Yvy54A1nthJMkR4Eico7QWgn6NZbotTHkl20GubqeQ2MtZZ
3X02q73TRliE8GXcZX9jJeBniiYfvAhFzVZ95KJBlnX3VFd8HOAIBRDp06rJaFmhc+79x32YUdMg
6K040yqGAZWYQJI24CH54aPvW9uOGPEWe9IZmkA4nz2ppoaHqtsK/mrhXQqSeCFgoOxswfVedJIj
1USsMEusjh3MhZsEyiuYiB9nq9R3R8jMaez+8iCRxLA0dLQGZh4YaWCrTWuR3LTsJ1xRvNY/4Kgz
BHllAQDfim1uLmvTpWe86ZY2CNCcmPUV2FmtoMmwJU/2f7Q4oCR/itVm6ZYpx5O9Z0ZWf1/V9vAA
XVnSWoI/jwiRt09gyVxglIj2dVBGcZILedrQtcFuD0oDet2oRf1iTKUvEtaUGwV7FCxDHv+MWCvR
2XempGoc3odQGH19OC9A5XasCwRthPqXtCB8C3kazQdMHXuhkzaHnUcxWZQomAhlxVxymNxfNmlX
ONdaAUwTqmVPyVS8HZJzUYDLtzxqR8KJeoRmeM2C+ZQXWk5G5aeL9qYRZnP/m09rSiGwGsqLyGTE
vC5iXHkgZo5Ny0dCJcVWeknlJY7rUMViUFx4DJIZS784cImFhvnDwkb25Qa5Y+a+JegshJzRi12Y
cWIrhHx+PIbsy2yeGCS1gG6flweftFpwzDVDYxC5B3qvEpM1u3oxhRIJIHkKzXXDjeKKMP/Mcldx
aHa2rKNjjGm9MGOLGyGLDAjJ07PQjxS8ukUJ9j7zJIB0qPiOMnRtV5IdJgfY8LJosrs+Tz5amycv
uf0EnnvRiFDouL1DcI7SieSaY4H1u8lw5UHBJmW0zrtoYV68e4euzqwfp7Fo84uQkAvfh7wyrViX
nBnS1+uJXXLaqhxqXxm8/j1YMKetb+pU7ztBcSJa6YRT2sakx3ivhtYZeNRG5lruiagHddShenXs
VLwqBj+6AAaB9rFGjDJv5mhPRAonqa78Tfqs1wVhBNlgCqRIMhnrm7o2FZW7a/Dov7W6TLJjb5H2
P84m2C5aL5sLXN5opvGdb+CUI1fIuQK/OYD0PZJZfKk5LnTUi8U3Rj8W/rq738rJGNOnW0a4ShuY
nVaHViwBzDdnAPXcEYZeosQfG1c7c4tWEhOOnt4nKbmWeagkB+Nm50Ox3oU/ihtOGKL5BU9gFevs
cLELdwlh5TaUPKLx9UC/zs7iLQjjUakuSBpfLTbN4cwd8bQ6ktwOIShM5fQVLUNdpMF4br/fOniO
gYYPGnqdnnhaSXgo8q2MkHv/mGbXwTfZHvMo9rDu/+mAXeRTRakV1nUQDue9Wr1RYDrdAlCuvJ2I
Z8nrrFVYxvlRj2VtDF3Y5jGIS+6ud1TCEZj40pXR18gsnVDDEuSS6488LbBBPUuCi6CByD1nsbds
JgLXV7lfcYSiDFMbvMKwJi794EAwecQqNpVsZYUYqbLkhOY8IteY3cvyxcMQlKxw7ZYYqSO2djHb
vLFPxRo9wowi7Yc0WOtKA3DBjpFXc0FGcx/gVTKEb8NkLGncNY/7YgqmXPplMM5sUXcyKeljfZqh
+oqby6ohUGP3bhQIswItjRmDDl8ofaXFTVcI3ImCwaNL+To7qopy1hkuz3XgFzKGSrOL9BrsIo2w
KfYAL01jIrHWqczm0zBge+5ph5BO1cHd6pI8XmuuqWVEmVgkUL8pBHbpdBEkc7TrNiizHZIONbqS
ZmfUGNlEKHYLhbkNMe70I2kNuZcrgbzlBXeoz6TMFw3sJwEoX3fkqEhr8qYiUPvMoxY4yD9U8l2e
QgrCR9VZChyqedxfQYX2b47jIaiX/6eCqU7x1qDjmbAR5sDkP7AUNNuESoEYUplbTHloaupO995b
wLdiYAqOdgjijt/vsW4xJrMLptX5LaV4X7UWEBOb7nC5Q5+ojbnaPK+AImQ2I9FW6Uc9iaUScqpZ
WO5BzbTMUFwindoMppt9cCBqLyXqTCT1YKIIp7E2zuF8sXMrpa4UILJKMM1574Za821vVZM8gQer
FfhbzJL2n4syl/CMHtFCjSEWkTklU+Ti8IfS4mD2Ssv8ARso8K06I56PasDBzUOx29/oa1Aomp2G
6q/598FwQ9tO8rtkWlzdXxbeogLQJdr+8X6yuhKSKFJrMP3O6LAk4rIIrO5KY8jfKtHCA5x/4csP
EXny7J8ntMFFyvOTwPoAa/HEftVT/UcIdYQUVMnrntMJAeyVgsPzRIt8cNV8g9eC41VahkN8T5Dk
s6riLFKdvM6QuA9axzarjkIFTdOycypBBfuIQ0WwShY8mfPP1ErSQzN+Ceeh/pCqwJp8GuhfPgPf
NJiDsi4gkPbciPJTrISwPzcUF/PuN0Lx5gmreQgcBACVFIB4Y6PE8ofVYP9DCjmvIbthgMbhmBk4
fTPoUxeOEAv9bYHdverU0cObtKHrZ0/lk6pn9wbC+6+KEG54ums759sEC9scy7W2Q3jX1OM8KiW1
ZAtNlr170n4xIPlqbloknKqCbhzymAkP8L1tu5YhaK/NLvuRp6B4lkbZSJPXztKVvB8CBEYhwh9k
ATJXA71TTjBgVueVIrHNPdNw47rVp0Ojvi2NJYXi9/+ysEbrJUPOlD+zed+SHsR4mK4NU+4WGCcd
Sf6YErPCaXZXclGo04+cGIJsDRiEXjyB9CtjKEsJnreozEwDP+UF1tnd4dwS4deNzLJoHyCtXAX6
OBKFKBgkvMyNY9p3T3ZrVZA+C+AQWW9t4z3BwZpmJQT2Oj84JHnk2tUkYqZDYM6qLVZ+3OAH2w2R
ptoGoagZAIbMnCwQdxmU6lvgPGRKAXEttUwm6CUu0Lmk/P3AHRT+sfqgw4A9Ch88315lgvffGeC8
GFbxS2w3xkOGGlRNdHy5jlsKFj+5PlkB5DeN80KZmBKyGbCpY0zl00eF6l1Yx9zxbJGBMkGaeiOb
rw6sOA3vM51d4pxE4OiKCG2QeiQ4npqHJE2xyXidpZzhnobop4zPbbMcasdPJikvBD8v3+d7sVbu
vSlNC0qw4zt2rYw03ASnlfu2n3BywrDvrnZ5OcWsS7ODknNBoi7ZFDl/BgZNhU0M6kw4lB3yTR6h
MrpPQg3aYektT7icvCU4ov2p3BrVtqZ1XIo1YVl/0piPawRxBq7ii0Tku5MPZ9z+iFNAKAeuYtDj
YsjRY/2pELa6l/xJOfW8owIvxvsSQBODlNRm7Ol69oSL/MhioLYpGVFv5+UPe/ICU5g+jZizZ5Ke
Vn7XEWr2PG39SWKHoO2kpBLAnxfUa1/yk+Gb3tSMGFg0sB73V6hcm1f9vNE6JLxsrIOWWhsjmom+
fPrPE2xLOTMNIwMkLLhzvIFlhOC1RrKcyiXIUUjY0az5trJgIVKnRAvRxHXT3LuHMZEuj1kgqC9G
BfHVP0Li4nzkbMc2Xi700Uk6nPl+rLVArl9zNjvVyNWJWsDYKC1rMDS0OZXhIWgs0P2+Q4GCDPSJ
Lus84oYRf7rXFC/gdQx8J9p1i93lIMaE4kK+KmY//B1CDb0Q4yyN+aLXIsM/lrnl0k9xve/e7/Zh
NmNgjYOcHtJL/ELa2Y7kHRMdWyYmrBG62hzUkgXJWc4m+vSsl+ba5X02sSCySyOLqQW/pcEa1zov
7t2tQxxtYAuDY7NcSmwwwczpkZCqoWLmEHUtVmuYYJCK66ltrfeJS1y95XO3cQBCst4SqAL1Yzh+
Z6goxT3QbEDrTYKu+OMGSgR6g53bmPqTvru9yh7N51rncr7G6pW/Ry4eCAU4L9stiiMyenRM7Q8I
g18sBG8D9VXd/pk7Isav+PPPCR87Lmmb6RVxoNl8vUp1gEiIWyKjOnVqCpw99MipP6SaXJ31gRh0
MGhg6xGrkh+VuRx7LYAZpXTKrMhW1IQDskUelDtXD4Wr6PBol4mAXX+G547PLlbD4xh+MMi2yiTe
+ey6/Mbw2Ir9H5uJBxaZ4o0wqItZEvlO5t/v1ypnk8h4NYZzcJempGrNQpEutoMEDYjRuel99PdX
8BE0wAQ+p14UtOEQ8tDkT+uOrftzbjrq0OsNd5s9semMeEMiF45PgX9/CcfUVbOe/wxP48m6Pk/k
AasJKnJuld2+56zLExyk+WLq9sMFwTnn82YTVR++0QnW+OEM2Fdt03O8FNaNjnoGEGNaO9cRTOFw
CcSaPF9qsiHtuS6WvW3Vh1VQAJvPGIz+nm+j0zy9OpjTI1Kp7sbvK9B4oZkHy5dyUzf+DdHfYunX
4e11QL4ROHl7P7KSePDFjAe9G2uhCDKXsWqy0DLOc8lNLJLLJ891uAqks9Z93DfVMg295DQszNjP
rVpR8ymu7RDCxVRTkK+DL9e7DgE35I+ZbpV2aHBfacMQecUwVupSiaXTx0qS1nDXlG4Rnlm6qmrB
OnXus2yjTTvB7RU/aXgpRwzSMw9TT5Y4af4UNY7sih9ExOxZbncpd1Dg80o+veS50gv3TJLXYKvk
p9wMfIpRc60ARpvyipRuIRpORUJh36l4IH1JSPg0+PZRZUC4+lbOCcTijyOHqJzmGJzZKiHj3Ufl
zzP98AsSspI9zsMXcfpo/bOzTQz6r4rIjwVYGuZL8lAuv4ppcv1SVThDSNF+up1kJ/u2xm/QJ7aa
BTXsGyJ5N8pH1+g1Fd4C1iviJlzpW+Xw1Kdl6U+Lw1YQoxd1IKMAykyPhGBviggClNDyn4qKzFAg
28fO5tR+VS8YBsW1u+o4kwNMZee2zAVNaP39ab0o3+63FiegbfOB7oRRtfSa4QO7tt9SmJZ2rK81
ij02VucfR9qpeZu3z2pUAWjdXIFj+SP06lbxajijiUjqS+EUhm9/d+Q2EsWESbi6OYLbVNwz7L6U
lB76ALmU2Ooy18Favwt5br2DYkDC83k5o/LA6QtEutyTQ7MFA1T0+r86FBM0mRzQp2BTvjIw+sbH
wAN/GEMMUT7L5QsSkIvnd78ZAR3P6zB4T/j0Qbf43cvme6BpAEMflPXU1qoPpHxFV1WhVeVDofk2
bSF8uDsdBLn0npYd2Lw3XYTIs5KDHI+jWfOtnEAW9LDEtNkI/W/3Tu+ii4NLPE2B6Zk+s3oIhQK3
zaJ29SfH9aUJ9fFP45YD0nHYNbW8z94SqHdHQlp7Wrm6KIvYqteMZIjAvHhEymMjvxcWKoTKdEDN
D9RbkOArhgNS8Ik067mspVRgrKFgA58WXXqkm0Qcz1EqhNgnRk2EBoAOF889XlYXfN0G46WhFxrq
cUqYA+GyibHiOe+3t5Imu2ckW5U7MN+E5+ksgo9l0wPZzqDoWnfkzHoq4uMMe5DDZ7kru8tGjqLi
vRdlx4g+IGR1jar91BIRFBZosWI9UAnp7/ZbPQ3bbzFDwMuzg6I4uqnVa8/R1KCQeFKkMutcDcGH
gvVllBQyR2hjyl6dFI9edYTXqB44BN1X6RO8uLn67nJYVC9Z19Hx02mvK34ot4DNq2oTh3IkVcpZ
h08UFa0/F8AaPNjHe6DxgOIEzikdJMbMOqbRsHPV4AzBzaUDeVszhwKN8QHCC0t62zZCcl8M8GyL
UOrdzuzRBebEC5lkjdrH2YRSzkk0r/uNHAYKfpGb/k3RMbF/9HzAb3fX21tXbmEA2f0tBEQzljJZ
gkuHT/XQOERf5QOPnwF7z3yhxxok5tTOkHvqC/Zd61Vn5ctLMgg4dglQyJSlR70ox0GUaisjRzq+
q4CQLsoPAr9fwfBHhmZx/119jphzurdixyiZugoAF/g9GfKY6YnkYyeXFSGe8sF9f2Yjj7NJvx09
n/Qt9yB3X8XX2eS/igOcpon29RnGrbmoQhpB2SvgDu7yYQF9SNHaAyL2d73wOp0c9v0e9sht1jr3
I+Hb1dDlTurPbflbCo/e8AYna/P/su+VxTDIzLwGYY0poHVc6T/yTT5QVAC4NzUVaQM6tPxrME8m
fagF7SYjwXmyqPW/uJNwCfcrYfltBOba7EJGebfVjOIKqXQTEYw1VtfG5JHxTZOiCh1vWqHxHm94
WJ0M8Olu2cNo2605w5qYM4o7Rd2cg1r+D74/eVD1+wllX9MiwUSCiDCSlq1m/57Q1v5CjZS7KSWT
gjwVcs/6RqM+Tgq33SxlaevJ1xQbqn4xwVsQqFjJ/QDZUBWUlloxC+AU7TUIMBTbIirtwv5sgkKh
IPWkiPq1qqIqjfras0w782Qr9nTAkRKuFwzutm+sTAU5nuevVbzA0O5SPOv+at6QaamAGJs/bo3g
1eMaw8AI/GjfXiJhZokD539RzI9o98VjOf6xtGOV8qq4QQt+R2p/24RQP/oHB+LEueiGcrG/kAXK
VEkSvgFmxM0sJ48NC3zGyO7ck6rYxI4S5rXxf/l0r0IbHnn6UCrKBi5UeLktiut993GB2mQSien2
n5BllPZrx14wZV2rd/bvB+eEOScP2juGyl9AoEVBgAoGtQDdkyn+KfR93gVZZ5vHMXb/qp4jzlRc
fR0uta6Vco+vLiY/N9mS4kxPLDeLxe+3Rk+hK0HSylv1gR6tzR9GeyLeWvmWWkf8cBqsiwT5Q+uL
rJtUIApWUNn7xl83RKc26MMXUmXiqyMiwelgyQyE7NY6WwlvWFfmbnw0XVy/8oc89w2QM4zcYo7w
YELytOZejrVys4q0i+cD7CuTraoWN+hYRc2bM7nkNvyYPNnbVLkGVp9iPkfegpqDGL/WVuQTeYZq
mjhMoAScpGGu97j/v00ZZuBhuF0aWvk++8C6RpQwOponCCVnGvTJuMHCpvn0S4pDvNvbTFE0m5qA
uJ2vdHOBc3REAflUMQBGXopDtUoVAvUxbu6k4UGInmNONmeulzvo0ucjITmyGwkhSk6La2I1a9M1
erCnFPx3dAhuJlAFG08g7KszAUd6MuSHlOhDF+OEmOrTVxj2gh3TQCRBUPXqXyciDiYSOtYuNmKy
BAmbUTKBlcTOmnMOlcoZG5lKiC7WCirYmL5LVveMIP4/wJM4oMDXxuc8uNY044UuveyYBa2DIABO
yzKwyhi8kmTf7Cjm4CSF4XZSAnWErVNSb1XCtUhK86ekG9/V3kefyZh4KTKjrHlgJTq9vQxvJ90O
aNjw7goiv6pxPdQYAyC2SPcEmBURiGM0uLAJztv3NrwQoFm0Vqu7ZXiNSrRTu9H2Mont+j2ev6tH
/6hrWhkCvQ2EKWwReOt7POZd0q5dt61g+Rej3O10fPHTni028pIsKSC9zijHfspHoDqpZRTXGQze
TmRQCpsdtqvfU8AXZLoxLpV7CFDAFOn5xF5/jliPQ7RS4p16+dBwBZ+XQ+gSAByd3kj6sa+Avjc9
tNHQyIYCD/pixlFDKzb9D/r6bj8+N7NsX1V9a7OZkFQRQcUc3lvZ2ISCxrwY+km+lUSlsVMVvdou
f9VD3NRu3N5UsMw52fLvPNoMcSB5279eC2b6sl21Iud85mZeZk6J7clwwGTj1LBzuAeFt8y6RJhL
RLgoBkrpG1N83THKAy5Y8YQWy5F5Vw0xLmDZlNz1bLk/1fNyl0sxfD9BZo6vW84MqQUE+mVielK0
dsCcct5mqFrps5+84j65tU1p9zxCOFoI+KfgvAdLFvKUrs8MX5C51hvEv4aVoJmNFnKDoPl6cuIF
u6QTK7tMD1VSUO5m114vH8m+hA6b3PoyklJfs0sog91iIzr3OpozobaqEFVe5yfOioSBklHLRTO2
OdBGBm8XRjLUwJNLz2GM1BkpyVAGLVIj+zVRKIm62suVSiP+eBj59r8fPd9FoSKkMBdFMe5Th1Ck
yDsq3jQINP/OgIPf8UNmhLEou4GEVJSioacmz0fFS4lwC2Iv07AxLNoTz+Z0wgmnlfrQ0WS6Cd6y
XrpKI0cvVYXFGaaSpvEyGYzXrTcnesIZm8OJ+xaTKS9Tjy+0+njry94ORlgerj7SAsIedAMacuhh
Z5sltslcj3WRQILO/rOgFPOVYFAlWvr4i21OwjbtRApalyddxVK0LjKqHJFP3XCU0WFUN0ojP8AN
8r4O+UCnfsRl2ALfiFz7iv4GfTqzu04UHgmNcVwH89AmheDR8pINrn89ha3DzQSKwJ3XpTK8TUnJ
htVQ7etEqaWH74u7iE++TNQOD2fm9quNwR86axWBXleiU0XfqZOthkUh1Zvqk+Cf9xLMNcMiqo8x
gq7bvtWAdC9J69vRA11lqaHOoFsxsR1K9jsiVnMPPkX8OUVWdXmtIVTVE4hwkW7zjjQF2PYN7QDr
Nft/pz9DDzqs4Gf1KxPeNso4p/CvLZe2UpuHQOvNJpVIVyqLGOLNUx6Brzw/+czSF+cA9LLSn3Ah
n3dHBrNLHCibhUtYLrpJN/K/9t3Bfbthpz879N/Mlti69oSAXl7Vq/k2mnwojVRgpLklOgXdR9g6
UBFvvofTuNjt5dLthxKfc7uP2gKZeySthwptZ/KiownhdenhfwODmYxlQFSUOXw6qpIy7KA3cU+H
iDH0xdsAGFkth8/YhJRyde0wIFQ7jjYhonC7AP5Z2gTDv3GeI6N6aFjIc+szq70f+a90pViDhsDT
PI6ygnyFWolqy7apVcmcKULEvfatJ6nJ6KIH5Mq+cb4jrZrC0gHzek+Pv4FtpPuAqDEqAYOs6PIs
Vvsp0LaNDjys1ScSllXbmNn13l9IhqcznebDlWJL7V+9pj6Tf0RNjGizBrDiOh7QLb0ObVg9CoFl
CCJMVRBKUBP0nTgWkBJX/rMlluuthan/LUfVlvOjkNBHM75N9syYjWl5Cjxt3KL3vkWybgAFAueH
ZwZrW1dCQZqJnQtxC9sn4UcenStQrpOFXMQBTXuZ5tGIGdsOLov0AQmTiunffJ4Ky/mGJti51RXK
8JNHNLDCbXywiYgcZuCdW8LsJr/ptntNs6kOG+P/wJcTRrzJmJTTwcQ2qZYtdhdRE+zdH3x3Y/4k
JkCKN59XCNPpXaEDvxt652MfD6aCjDJ29DNPiqckIPbK5741VwvZoGGf26gV7jw445EhuYI4Wuci
3uK/nA53Dkg0bpUgZDwf0aDyxJEtXvQ9zHDdEIGb53Q61nsr9mlfBo43VbjZh3Fz1Y1HlvMk+K4f
m4hqqpELrmbVM/NeK6iXsMnGT3EnXUuEQ0t/Zdaeo4lNXGabVHkXWJjERyroO/ybGQU+Pwvn209K
cMNZuXcCANRsRQ6JhrDBrYxPflVt0sgMXQWsguhAKn091cmr+nglwP2uXOO4FzKz+dgb3rxluQaN
IV0+rtNiDkeffuxJOLjuKGjdlf77kriIePniZwfqHIUe5h7qM3Q2rVC9gwHFOw8Rp/RAVYCNKSUK
E0r28tlt6RHg8s5qGoLskhrzKCKJOk61qK3cuvWLuncGchwAE0lEXpVOjNUObquPmn+CyVJYLn9E
Fd4rAEx69qb7/5so/RWdqjhRIBGEXIDdkr+jXF7jeYK0gNIyBl0cu59qBaqhEQcriKqCPkGnO+rN
5pw+pgPfkxXWUcY8IXKgpY0s+GmqgM6/tk+swBZ+khbwbI3AbbnPQvU44/zWPWIMKsYJPCWqGpAq
CirqBB1qR27Vv94+/Wdy6upSfenAN1K6k2p3nXjOjpQkdHTc+CXjWEf9YMg8pgpgW3nu0uG20yFL
lZiAEUpN5GivyFxGA2jYoKU0DUsAocIBmc5BdjToTEHkMTjrSYovaRSsYRWDszvQ9PzdPaJcOUKi
wsvE5BF73+3HedmzOja5SQrVhahfueuaW74BVvnuh+hS15bqNIadu+Q+6pLe+NOJIHV0Y35sLycv
MkyIUcr808cqVbIYS0xrDKB2S57HRQ5R2D2I/Mi+oOR3BEEHixrgtNR9RckLR8wsHCQ7AFpsZm8J
aCLPPO+nurc29EB7XSRRpbbHOHADwxEJx/9lVG+rtxUoV2nwjQgoVss89+UtFb7jj7Nl30wVEp2q
KprvY2BLVMiXnv0ovMDIkegWG8fTgRGTHouvroL+xfJuz539cVn/fG/QPoAEPQ2hqjy360oVr+MN
/rxb8vaqZrIm7AI/bzEZmtQ2wW49VNimX7tmDTT2cqh8TqRzQmAbX0n0z3h0XFYhOUBEztYz3fNt
Et/4iS7C0sWnOeSQTDrJhBSLg6z6crDkq3/VWXT7LTKLDel57cqABUixndAW2+3kNBr6vzhYOt7A
ibKBFDW9kqV/MSPz8X/I/3XFIXQ4moWhANyXBqcgMPmfq83d4yN4aMl+W9SWSFAygeZHQCwOQRDv
ari9CXMg1Ys3ZL9ZWN2yNcLlhR7Vwmt/MiOc3AVoDKBKyFWgGO9n31Ug2BU3ztvyq2pn8ulg26mc
o80YChml7IzO8e3oVfUwDibXeG0C8APpvfEVGqza0T62OgpHOubPLt5XAbNztGkyGoUnTu92nEp6
B5UHBk2Iq9COTgwGdzGAeM+pFNxFmsorSchq3rqfJidxgDia6W8+PHE7lvFENqpDv3IdIWuIZ8oW
nIMFYLvfFm1bv+g/1uYGlpQ3U1Q2bbedeMx+/PTtQXRagvPTwyCAVqxpg1uvG8xkHiBKpRbP05uM
v0icAZE1rcfGdhJRz6iooPDyBkQc7Q4eA5i9Vf4Ti+VWxzS5v9G8GOYvjfJP4DGFxwBwcoVDM+P5
Cqf//EDVFvJJuvLqTN25MDvoFAmIT4P0f4I09KnExFyE8Ol+F1TAAb74gq9N84EhJ6bPnrfYxW8g
AFbZUt7C5cNk9b9/OiyQtRcp08Jr1PBtIO+jvM+VGiiP6QbfWUt/GXNE1WUt37f4SBduxu+pDKZn
mw4RTEgEbD/GnoMcX3s7AfytYYCtg3QieiV4alOvAc89b7IaaLhNEsPozRRB2sJDladmTZtQ20aP
Tvczx2pZdMObDYtXs3NTeB5UnqLt0lQpr5zD74wAvUpZUC9+tKlaw0Do6lVfNoRFsLCSJJ6PaSeI
K7XKIox28cbZqFeubgqpx2W+sOQub5elh0HcMqwQsR2Q8o06UJaXuxAtCZ7Twgz1/S6l+QgXs4uy
bjJ/+/79dmTyzUPx8ZgN6aU7R9xr68yRZ8KEzVH2duZi90/RiTQDDhiNi4ajXNW43yr5t4xi1xhk
0dGbett/sUAp3YuDNgdU4Ai8UsZ20KNLFr+HtpZHXRfLKHd3OeWSTFZjiY/BRjiTcydVCkG9vGdb
oz/inXDAR5N3drAnCifg8BSGhrwwDJofoGkSHD3nQKWWInkVTuA9eAPbCJ04eFlpeN7bfWCLeiJd
mID584sWl2URuZpucBC71G3fcHpXKScMb/Ls7cA9xNDfJdlB7qFrgIlc5NCbOENmajB36BKNWByG
Azso/7h2wWw4b3Md/ztBIcX3cMBRPl4ug+AFhdN/jayDkp8BbSbZPKBxP+uOdzJYwqjPchpxAket
a+BYdHheuqoKuGM1dIoFo9sj7L6ms+H7PY3pUBQGzwMDH1BrN8JMWvELpF4MUHrP6sYkqNRMKLHc
98cxyDiRHOpuFZQQ9TNX924NYM0n2n0129wrGeZwfqrO2RQ1Wh3LMXtZeu8oxNtfWCsxqwDxsSzK
1rdEJNpSrVdWxjP9kxMGMlZIp0kK+VHrBf4Lu0WHNpGbFGxigrj0b6LdXglELqMGLS0xiL7rTKTF
Vxjh+2kdA82qr0/yOUWn1mJ1Z+JPauo8pM9L6f02TCgoc/UMjNhqfXC8fZ7clqNw4TGna/bQEFep
ESJfj15DDwbFXUq+LzuC5t7MzUy2BxGXyPesJ9dR3InxqH6ERVZIL7AHFs8GSrkNje9IB4ujRQvH
aBsuMXVSE4JjbqCa64vFkhIepr4ATEHf+1TMQ0Lrl+aW7PXV/wey6E9HbckKQUax3ASi3htkkZmL
buGMhj7167+c9VfaDQ2bCg4pwi7E3PO8egInIgxpqZVJBxyj44yPiD2CHc0v7UPyO16k9PubUhdM
ShFv7RGfoJfVd5A9sLOKyR8ZBtJFm7oz0GKoUh/lso2U4qXdNhakItmgQvOD5b1TmFM7JDHBLM+0
sRAfTvdRTYW/+AIMuOsZ+3OQlqwXm4U2OzDAwy+wPIktzQpHnoTwWTlbcQclQVvmMgEN7OWJlvAp
5AVFXxoJKTArsbGP8w1bMymaNfqFlDuCnOK1uaa/UoO0vY2mbv3iYasszqkSaydYQqwZc6meh04m
qrKdLlOt9ENA6O1dgf1tyd5EZ4kBKaAKojUfJfAEuaH8s0tSDRl7xBR2gely5WAQR+Lj/W5GNQ02
cmFmDaFMpEbswtGzLVZ/L0fEsrVTp6OMiprQZP155DuOsU0oGEhlAkgfe0iRyJyfri2bWnofDubu
4F55kPpoq2XGbhfik7GiIw/89AJxnS+H5PjoUjKktik5IpAPsWgk+KM1kwb363vmCam+Y/vbYpG2
AjNjL4Xih34JanWAvVCevjj/wEmLXKggObys/77TwONCtDobIkNTQBRF6jyB6GIszTOgl2WpY/Qt
9RcQdZ5MvY827Ga8IT+pM62FHZf68drXlOMfsCudEYfm/WaZaFqDLoGAY17LVA95bL1y0hltErkP
K8MR60uJTZBhjniPnAKn9heaAsj2fzaXukpgCVm4l/U4qWe8aofRlycKCl2gdkDAbxOUTbpYi3K4
7S6sAYmwETe9U+72raPnzcBt19TXMf6+kxgzBkAmP1lu7q6zcdzK+fQ6gGnxex7MPPA6ZNvo0eS5
UkQBQALbbQdNlpKQ9T4FExwXn0Yb2M0dODgFV/aSOVm4ZQlaFomy4SqCywLCDQp2IFYDOAMaAcXo
FCQq4fbJlOePvDbhT4SclW7ryDrF8+t16Al2Zb9K9x9LASDh/lRHVv3zzaOFkbcpuyQEJEUSW9Tl
Lg2wMwLQqzLqKTkS5fJ1yXRLVaymtN/XiBGtlx1tkpfQZ58WOPQsxM/ueOevbsej9xDKYiCDwttf
kQm3qtr2fMYMcOJMZqqSsdvPoPh4PVHGcO4a5Mq/UwfXt9BsvtC4ZnxI7VrR1XHhx5QfTeSdN75H
69pGkHkqbURQZLrDj7uC0apVmj2LbUSLHC9xtPUj1SXrwBbrd9HXSC1SDLWMAK0wIAEnjh9YsEPU
crCxnOFnXOc18Qk0Z5E8VezzmJF7aWd8PYMzHcjMjhVDdqYZI1yOcnP+TT2oSbKG2ap2YfU11taI
pG2mCm8Pg8bEn2J5voBHVCJHa0NP79yRpzlAurJ/nvcqhWaui3i7NzsG5SQDDhRvDJGINKCX3JAB
TJO39OjtSB14HsUA3jVtduDKmXb/KgioU3wtavKQ29JRMzlUP/h+DEUs1gERublTb4wHyJSAVRev
411AY/3933mg2azOCOuPjR92MlgYGQpkk1Q5OWEkktj3v6Hcz8faAbevgrWl9LbU8MTUrdTfhAKT
Pm6w18yjAoaWNm6q/g+At0OepvDjNu0OoNgatol3B3RSoVo/zrvMds2ZtICtzc9j75/sSlTv19MS
6VvKDbl9zVzkpiXFZFDCzknzncNKzO0ijHdLY3M1JYwYga1QsneBjEaVuZ1S6eJn7EWZOtS4qHDA
WZC6NTvtaO6a+iq+H2ubnFO6K7amyI1ZzPvRz5yio5hLLPdwRYS3iyP6nIzV818glYJcNM2lzk+f
4W9m3H6nFqH0/Qczh8JnCzBoy+7vUuLKc63nTw05pMcPkqIbvSd5REFKB3KZMkBO3XyhXBoX7qgA
YIGF8SrTrdBHob8qeix4GhzsvgToY+mE4c5B1PkuJxIRAFv5wMgI452iJ9vnaALWnIhATqIAO94F
V3/Rglw2LCsYRYQphmhN+HaY9Py/wxeEScueiZIpBQtMxl/f8u9mE09pWoeOkmHZZI9Kpp1GaY7+
SP1OzQ+A3JADVZcC9rQ0P2XrhNR74f7E3ibOJSBymT1IZDcH5ekLTaV1MESnxRfkcQbfmB1FGL0S
AoWTSgSbBduo25bCx8kZRwUKZF/A9ByhJTW+J61MaSfafMF1Qyl1b0eIf1kSGKSenqm6hO4APrxW
1bhh+dg406x7LEtu8GJ+6ADqISuYgwEedOBpPlDUBoqBG6zZWLhPTmFaB5rwCuQocoFOKTn7/xi2
v3ximQ3a2pIIUw6ioSGvGiXDedIzp+dQD9ms3VUrspJvAgLKi9WgE7Q/4tfBiMfevo8bLZpltUmW
DnXAixFzrIxax93v+CFtHuqCKrekrtgVgxA1HgyANmDvAQl/qYbpMyCs2L1kmRDKEXOGOV1UUGrV
63TUZUQ1kvMhaPiFOUwkJ9XKLYssHcPNdThVJiHzwHbRE7wxlwZ/UXnxEqRxtTZyPJdeLwXikPZu
kMmhH6AgIsGPf6fXrNEXSGYdV/YIvzeWYY8tndNHUERu31sHMTnQc1KdSTbQ8kHdNGTT/LmTjjpq
LHL5POFR2gVzND1XPfTfw0VsCoGYhepoqfZV///7SLgQImK2bdf/qPrXwp1cp5m/dGLt58t7PBJS
omHLyNoJrO5G6sPNjMrN8s3app54KxRh/wK/BJRyoLdCcRAJZ73nXD2ZVijk75ddGC3GuAOkroos
JSne51Nd+RiyAZsqNqrmW9qmswLdXOu1vpWuEAMFnAZPXm/xK+cyNVfnCWukHyIwsZul3isZAOC6
UX3C8xVVHHifp+1XhVNwQemQMbQ3vnsETRrj881x01PWj0YuAIKEy5PWmlDO1mjegoJFIz/nuqlp
QnE4lHE2do37xq4yIdOjQjYHOoh3l0x4jahDyiU8XySbcamdukFk8MrtJ8H32oJySrN6Ut418vcz
wb6lVBoz/sZh/CW35NvoxQWisQrl6zmwY74EAyQ+vAVHrt8uDM0JCKmTPpDkeNeotPHrBrr5MvV2
EBmUtGP4V7R8qL7ssS8+WHdJnQLgbw5w1Toigk8G6p5wbLGy7pAPr/hcKLdEVkKGs7lx7dKbt5OQ
czFAfcqPjUB9nNbjdqlJeNSIGIGsnfDjAcT82vufsfIjw2ky2AaXtB0sN1R/jrO+IX/kODDDHLHM
HfmQYdx24osDHAdPIbkUTxQO8mJ7e+4LSPNsUGZQBIb2OXq4/ncGyrq/Dl856tPGwd2j8d/Ikt1M
w46mG3IEVZa6Ro3VP4OYY1w/AI163LK5aq589MoLMC++ofoMZ32u5GFLvtdny/W+S4CSkYDHKPT7
mccfjxuosNhsItzu8Tu102bURd4+2tfvuG93dOk8vija3xe7kW8aGm1/Ay22iF3tm8FppQKaEcV3
U4gBaM5FURZYZGJGOXTi+QQo+SzZZBm6jORGMxzKBM0pdD9djyoDHRqab65qjbw5vWSR+QrzIFNO
03lhNpUIbep5YplZue04ahYGY4hlWr4q8Ibm1vTkmZWTSXc52ht/ToDsxOX9sWRkFhBfACeFQalE
kcudHGRITLbUV12p5kS06KOLGREdDVxLG6bi0xhE0mCG+PofiLlG97gnxDX34XZzD5cEs/0KymOm
yF06TwZsEkK28wuy15MAj+BBbZYszzNhL1t9liZLmu+TAv8JT7pWPtizULQiYXPPhqS52iCtVWV6
gl4HUrPBFEe1r1u69i4fIXi2BLyrUmM4AQp2Uv+4gQVCFkeSc1jFOZh5fRUQjHHa+5lBjSrErPst
ZvMYci8oQrOi6tjuI+8C2mmQvXQxpejvEIIUpxorxI8nhQKgSWm5pKBhB5RXRMrPg13SwizS75A/
oHKgk6nU4jURGxL4t7XE4oy5FAQsCtxqadP8/ICaGUAcN+lOFRh0UM086qZv1gB9Xd9GOuJh5QtL
RFDT0zG1XwOOgayEPIgy/W2RDM58TR7mOyH4MZvd4HTpjWW9ls+9tX3xcT8GZw6XgzrJruulwtEW
qXXg+e0kaior0ChodN1VLoq7m4iinpCB26A2aepjaFdGCuVeDrpUBNa4sPpcod5ZFT4x2zi0fzVb
W7un+sBlRKqTwtPMZDW+fCbGbwmM34pxVLsyrZ6GUW/cdVCM3c0pUfBHOCvwZSN/iUcjJ44LDcnF
OYfYB1ylxTFjMUpSGV26Anz/AR/IjpamnBbT0pI6ZXPg5GabYhLGlybHeIoWzPrR0tvm43LptJSL
IBNcwFDxKJQyI28mSVC1b4khHdqY/A9Cl90QSm2gmGJveHVA2MSf8RXd72LE74mp4xrI1zPHw4Cs
kXP+eFUqhsWyatR4sTozs8VJ3lUI4UcUjhvGl0CLaHdp7lWJLE2Kw6nv3dfU+Fw4Ig7qvnvszLEH
XzhWSaCDY9HeY0cafAjjsfH+KQ/C/tPulYylGeMSGvqXL/eeNXwgHLOa4uAmX/ZyhZSu1EvtDMJf
Dtn/6hhcstE93xAzL7640XMXRfuIK6hiNNP6+Pyj9brw6VYStICLLVQ5WtiQU0DLZqZVRAHPO6N8
Tq9IAbnyl0mKgcBjxYnFTg4e/xb7wX+7VM09Otw2jlitCFeUEb2Q4Qkqj18GC6eqpIExlqQcgd8E
doPuxrrJ5VCvs++fneIlwQs9i2Lrk1YFmQdbiaKreY+FE6k087MGHSWTogADiZ1nRaJKzsBiVcy+
1tTylqtUTnyouAlq7Jzrm5zmzWkpU4/41Nizc4NGHhj1Fg+AyMdLHXDtUYStu/DrRsgyvhZ2es+3
b8Qh6w9ufNHF/nQ7+j+y5YDFZqhCVH9rHkpAXsnolG4DSrGaXa9PTeAIJg9bMBfXdsWSSUiAE7nX
Q3sLzX3NVeAt7D32XEYXnq9fZ67UXC1AYMUTYaB2q6WeSHPchrS8Z+SPU0uOYe5r/oF4PD8KCntK
ckcKUGTzNUhGzGbKaS+TB5jNktTlQ48pgtBQzH5u7bTXvNVJ5UNuDKZs0ElkgdgcTB9wI+0MkaeY
gOqpr9xib67ysSoeIBkDrWAcgWr20wGOdr6nUoFOgrZ4Vz01gNqGKLDCCXbOAE8iTfFsgvAVdwtY
fuqrBqqWuFxAp9EyUspMQhXLlTT83XDhEpYMkHGu8c/K6XcR4GzviiINP7kPpmj3mDDkZwFk10dk
uGYIihlGkEN2ihmuum+/yT0F8HwqNkmb5nJEtspW2mth/LMR/gHqEgX4HdHa7XBsYL4j6yKZovIL
9OnE8QbQILzlgk90+wYqDSWUUcxheu5yxqYseMhFrWEnZMtQPAKxjObvjBJp1ZrIxN5N6l3HbuEq
Zv7pwVUOjGJ9Kb/ocWqA12FTGwLTL4gBTj2iYn/sRoHwOLFAA3vwP2Zozo5U4kw+bChcHnP14lfA
40qAMpSbhMTOdLHw3EEYNzbWsOGy5AwkcLGAiQr6qbuYOeYEfxLV5sQaizK4CjULO8wPQiwkIRUh
BeYeyyHXvzkz6e6PaUN0IKmvqnAWDFDE4V68mibDWTL3RH8ZgTp1pnrQ8w3lCegr9bvHqeMDSLKc
DC3s3BAmGMwb1MdkQ2kBO5g80iuwYgSkOLyem7C4LhCSjhYIVN8Uy/VY6oyOS2rn+yd4rTIp2BcB
NGkcwGcsD0K3grRzXpc/cb2JG4v56Xp/Tjw0OTl/vJTW8ai1JT8BjN/h7McrTwO1qrAyg9gR1mPK
lsj/Pd8cBH5j1pCOik6+Y9djrLMjGV4apjQgd+Ai6GHwpNGPljVMwZ0stO3JdSNA954q7II+R7La
sBWmFQ4hl95KvXCChPD+QpvPn5C3wOG9SkvAz++DvGrgkDI7ueug3xAoGDaY8cu7/NbHjOsi/gix
xtbMsBiIjVG8mGbqBaCbh769bBD8r7tcALMhm6vfHyUqBeGItG8QYDwvsyUZ+fBKwJQb9LWRsTqo
d8TSMz3nyRTAJljgIcm8ewq9iTA62jts1NBBffsfFjPuizgn2ZXjzf6o4Kjbsk1aRpREUXJLSSHS
dzZHc7j97t70tZIvUqolxn+fnwfNtO+//G1sIoWGErwZPOX6oyTJ4rp+5JF3cKQFM3J2vIs/Qejn
hg0mZmjhFfEnG2gp5c7WSw04HwPvf5LsPXZMZ9GTRglt5ngPbXrWZxosXByZT83t+1nfS7KhOe3K
4V4KhlWTVJ2GMssuAZLkscsVcBVmYw/a6dcF92tq8r6euC9cQs4O1UAzme0wc96GS1+hVHgeGm6D
sZU8v1uqLqPQWxwgxF5AsUnMQLSQ8cNX9Ki5Ls3/bvny6yXQWiG86eC+G1HIGE/0WkUBAuqmEkEQ
ouek9km5Vs3099Y1bMsUFIFdXkgvZ8SGJlRi5kLRN6Fp4f8544WB6uCC8NKmBMKfyVTwWUceuUd1
zvRJ23bQi3V4PCz9B+ehFvLiWqu4TlNJBIOmyITyjhTWNdx+faTc9VppeC3DGD+Zqwej5s7zQ3Ho
c3j/l29Vr+5BeOZ2nB/4O3chFTmO5gfTfAzWJcyBusKVI0VZ1dqzpuUWuyPPoDRY/zKQpMC9yBRl
ijjWDtKIEzLnOMnZWxfuC3h5NaKNFIwOMAJvTxOAw/joqdLr5F9iOWJBPDsOpb21lBAgU7U+gpKR
+qcN4vOsPSuZwTBvaZ1agJHGpInwpm1rLx8yGh+g2LUrSwwYW7lLIukF5rJbyZZzi5sgy2qtwqRW
+2ajpzffT0/IzrJth4Zz6oo86rRIJ7SEmSFsPep6JCjkJXOWqEKxG/DbEvdH77pQOC8aQLUmXn+J
/ocSxGsjBGmDZTRax8EDuYKjawedyHFMZi4Lg6M3siR0or1oA7ehSTPNcwlkDJrCNdmGxaVrNL8Y
5BrQ+sHTV11VlWb9qQXAnLJc+GcAC87fCt3Gbif7s31XuazXqOkcInf/4nO4SQ7MQ15WwXgAu/ms
NgbHTpDX/J9TEj4VF2cRCbp2LqRyvNS4VwCZNB/L65gxZlGSRuqivFEwsCq0GrUn5UJGIHzKjt+e
i3eKtE+e/ZDRZsxu2HAh3WtDk7dnHoBsid3ZSBtN2ioHmbgTC82e1QySv+zOLnCnAE+pY62nMwET
yCK8HuBt746VVmrfeT0v0UwUpqJuqw/Bledo2AdmBxrcGfazrduNUFVIYPaxD6+PcPhlyd5md+Cm
MxFVWGikLJPGdTGwwEwa8LyFODfz6kNuOICdLJcTk5HfMffYOkNQiDkNj4WxWw3PPkng1gTSy5DZ
z387V9QyZ1/IYai7xt51XWTyDKVU6Z04PkYcd5ZBj9NXZQZHcsSLz9GqUiMddtpfWFr8hw7M8oV9
gb02OOmzQP/sJSlI2FE1lkbGt/d/IkiAzUjRyQTBr2+L6KwDGXc5XNznxL7pZGK0L0+dQf5X1wUx
UdQkjEH3QU+z92OzK/USQW8Ksxv1CmT7fGwc4dDH2tkU+xV28os2cc6/8hGnumVbmgyrUlA9dN15
JJS3D8/1Kb0sEqZ1Q3fCz2PWcMxR8Nr1opNjt3b3+GmJ8aRZYIgxroLWse2/LrefX0jhYtJvacNW
mUtaSjndNoSqdVQVYDVXOS/5sdE3KTRBk/OsZSnJS+ep3r1vidg87KVMsUFOoiocAOsl7C/hlhTQ
9quYVxY10KqsNrc/L2d/4xs2qEkzUsPWeKtLReYadH36eXVWAD0TfnonHj1IlTc8BFulNUEE2SO6
cnxbapr1qR1hRaTYpUUBzD/cCtSZCpfdY4A7VFSe3iSgdFTTBEhPvM9l0DT/t8BDrXjxBpq4Yl64
irO3xkWccMV8xKGeaLA8eeQLdaieAtxh0HsoUeW9juVFOYJvrj78J42mmXWfXrl0lgJwmWzSj9Ki
lpSdVbfeFQU0cjAs6AWgQCjjUUgssMqbDHUgFKHuzMTcY+OQSN/KXtbqZDpvs1CMZrdlF/uy2JFD
YNZ4rKni2Q7a60IQvAms5mtUXPwI6AI7epS/OecmPWD1lym9P/swXhazywzxKGvKYieolLEOG5uh
/ulY1BK622SI3c4ZwkuRXljRu9gNciL5AEgNHIOXYtP6P1woHS9zyEkctljb8PfDT4VLYDxLsmCg
eN6HOVY4qAb6JgmrusLr+sPIizyPh58RYTOuy4rE2kQ21bVoJjV7o2Ce3Z0b5aF03dhmiWeQXuXi
JX5vMY6e1nz+7AwxuKHmgP7LUwS1tCBfCj+k1upMO+TCoNEcGc5zC2vjSA0ajUCBE+MVCkSPKLrr
FdASg70MdzZbUVKx8cHovn7MbyGAZXtfbfsgKGfD784uVu2MUa+DqtMqhXN0UzIuZkhmHCUmFIAm
MoSfBwDZbMgvepxtcN3bYkGeXcCzsB5NTvT3j0tFPSEyBxIpr6T8EEH/fiPD28p7jUuyy9Zm7bmF
lmCfCmdA+ZS2N/N/FVtcchFZnlVvslm9f5X4+hjPfHIXv8GsPXPo8Kam57HpyeWjbC2Ux/iYWYL9
gFb6X/asksp8QqxuJyf2Zx6OVMsjhuOBunPmL/BQCM+huArXqmkWeSeHNTlSOsTmmFURRZ//a3ss
aMGd7uRpbf3hsGFjfIcD3jEzA4R8Rl7FexNzAUy09Kohb0vO/D+d+iAe9JoQfXRVjH4f+c40aG+a
pPAOApSEncR8Z95Lgb3gtgbkMa449BnZQvxe6fb50IVGqSuuyH/mdc0ZIyUwcpWmIGApz+rYvKsO
95vGRZCCrt6EU/alcHTFikgGJVb/WxoamesbtYiHc9JxTZhl846pBa1rm0Js7A3omhRyhFj0YkFw
tUMlNc34UigYsuIDBHI5c1KhPz5002He2kw4Lky8ww1FPScON0UPFkRwQrsSiqsf4QZbEjiak6XZ
sx4+ox04png2ZWVkbKMOlswk+1Bv5KoeNt/OGr1HxgPP3A27EHSQ3eSoZOoS8CUUPmhy5SC7Tury
B58kLBSB0TPc2lmGvjKDdvJgB81om/BdT1uNk9QjA7lU6xAGwwK7OZaDUzOgfjflT27que824ZUM
21e9CENxzFgm3hr9hSHxHJvYlTDZXBEODAwij85A/BOTkoeU74TTtaknWiFIcdoL56SbcY1ViTUN
r180NaW2nQsVkdMRqI8bSV16QcPEpcLZI17BylI6RMHF86ZNYkW4LhGXLQpRaDBkBQ3D2I28pp+v
hgUtResP3Mbl8azMxlsB4YbWAle0IitAkYfvxd7VDWvNCosiU5lygA4GYn6muG/EOUA22cXO3/6D
uNZoAR/W8eaBV4g0WCmEwj/bHC0F9dOPZqF+OQMCuD/mjcrapmELRkOB8Z9nxJYfr8dGnpUcCPNA
KJoTnzEqwC/EMBrztgsQ7R9hByBXqhWePpJr9SyGsEA4ZY6jdHMveDiajfYmGy5UPhKPPwZ1EkCa
q6aNkzW2fLdiKmuTqOX6SBHuRtovJSvkYSbvk48cCqOeKLNWDlWTz/5gg7qrBUHnHiXVoBo9xvEN
TyuhnvRv+Q==
`protect end_protected

